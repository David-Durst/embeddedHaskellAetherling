// Latency = 4
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset(reset), // @[:@1297.4]
    .io_in_x289_TREADY(dontcare), // @[:@1298.4]
    .io_in_x289_TDATA({I_0,I_1,I_2,I_3}), // @[:@1298.4]
    .io_in_x289_TID(8'h0),
    .io_in_x289_TDEST(8'h0),
    .io_in_x290_TVALID(valid_down), // @[:@1298.4]
    .io_in_x290_TDATA({O_0,O_1,O_2,O_3}), // @[:@1298.4]
    .io_in_x290_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x297_ctrchain cchain ( // @[:@2879.2]
    .clock(CLK), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule


module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 325:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh45); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh45); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [31:0] io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@512.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@512.4]
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@512.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign io_rdata = SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@539.4]
  assign SRAMVerilogAWS_wdata = 32'h0; // @[SRAM.scala 175:20:@526.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@527.4]
  assign SRAMVerilogAWS_wen = 1'h0; // @[SRAM.scala 173:18:@524.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@529.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@528.4]
  assign SRAMVerilogAWS_waddr = 21'h0; // @[SRAM.scala 174:20:@525.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@523.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@553.2]
  input         clock, // @[:@554.4]
  input         reset, // @[:@555.4]
  input         io_flow, // @[:@556.4]
  input  [20:0] io_in, // @[:@556.4]
  output [20:0] io_out // @[:@556.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@558.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@558.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@571.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@570.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@569.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@568.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@567.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@565.4]
endmodule
module Mem1D( // @[:@573.2]
  input         clock, // @[:@574.4]
  input         reset, // @[:@575.4]
  input  [20:0] io_r_ofs_0, // @[:@576.4]
  input         io_r_backpressure, // @[:@576.4]
  output [31:0] io_output // @[:@576.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@580.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@580.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@580.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@580.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@583.4]
  SRAM SRAM ( // @[MemPrimitives.scala 715:21:@580.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@583.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@596.4]
  assign SRAM_clock = clock; // @[:@581.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@590.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@595.4]
  assign RetimeWrapper_clock = clock; // @[:@584.4]
  assign RetimeWrapper_reset = reset; // @[:@585.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@587.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@586.4]
endmodule
module StickySelects( // @[:@598.2]
  input   io_ins_0, // @[:@601.4]
  output  io_outs_0 // @[:@601.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@603.4]
endmodule
module RetimeWrapper_6( // @[:@617.2]
  input   clock, // @[:@618.4]
  input   reset, // @[:@619.4]
  input   io_flow, // @[:@620.4]
  input   io_in, // @[:@620.4]
  output  io_out // @[:@620.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@622.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@622.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@635.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@634.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@633.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@632.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@631.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@629.4]
endmodule
module x291_outbuf_0( // @[:@637.2]
  input         clock, // @[:@638.4]
  input         reset, // @[:@639.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@640.4]
  input         io_rPort_0_en_0, // @[:@640.4]
  input         io_rPort_0_backpressure, // @[:@640.4]
  output [31:0] io_rPort_0_output_0 // @[:@640.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@655.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@655.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@655.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@695.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@685.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@687.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@655.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@681.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@695.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@685.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@687.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@702.4]
  assign Mem1D_clock = clock; // @[:@656.4]
  assign Mem1D_reset = reset; // @[:@657.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 131:28:@691.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 132:32:@692.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@684.4]
  assign RetimeWrapper_clock = clock; // @[:@696.4]
  assign RetimeWrapper_reset = reset; // @[:@697.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@699.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@698.4]
endmodule
module x632_sm( // @[:@846.2]
  input   clock, // @[:@847.4]
  input   reset, // @[:@848.4]
  input   io_enable, // @[:@849.4]
  output  io_done, // @[:@849.4]
  input   io_ctrDone, // @[:@849.4]
  output  io_ctrInc, // @[:@849.4]
  input   io_parentAck, // @[:@849.4]
  input   io_doneIn_0, // @[:@849.4]
  input   io_doneIn_1, // @[:@849.4]
  output  io_enableOut_0, // @[:@849.4]
  output  io_enableOut_1, // @[:@849.4]
  output  io_childAck_0, // @[:@849.4]
  output  io_childAck_1 // @[:@849.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@852.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@855.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@858.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@861.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@893.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1011.4]
  wire  allDone; // @[Controllers.scala 80:47:@864.4]
  wire  synchronize; // @[Controllers.scala 146:56:@918.4]
  wire  _T_127; // @[Controllers.scala 150:35:@920.4]
  wire  _T_129; // @[Controllers.scala 150:60:@921.4]
  wire  _T_130; // @[Controllers.scala 150:58:@922.4]
  wire  _T_132; // @[Controllers.scala 150:76:@923.4]
  wire  _T_133; // @[Controllers.scala 150:74:@924.4]
  wire  _T_135; // @[Controllers.scala 150:97:@925.4]
  wire  _T_136; // @[Controllers.scala 150:95:@926.4]
  wire  _T_152; // @[Controllers.scala 150:35:@944.4]
  wire  _T_154; // @[Controllers.scala 150:60:@945.4]
  wire  _T_155; // @[Controllers.scala 150:58:@946.4]
  wire  _T_157; // @[Controllers.scala 150:76:@947.4]
  wire  _T_158; // @[Controllers.scala 150:74:@948.4]
  wire  _T_161; // @[Controllers.scala 150:95:@950.4]
  wire  _T_179; // @[Controllers.scala 213:68:@972.4]
  wire  _T_181; // @[Controllers.scala 213:90:@974.4]
  wire  _T_183; // @[Controllers.scala 213:132:@976.4]
  wire  _T_184; // @[Controllers.scala 213:130:@977.4]
  wire  _T_185; // @[Controllers.scala 213:156:@978.4]
  wire  _T_187; // @[Controllers.scala 213:68:@981.4]
  wire  _T_189; // @[Controllers.scala 213:90:@983.4]
  wire  _T_196; // @[package.scala 100:49:@989.4]
  reg  _T_199; // @[package.scala 48:56:@990.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@992.4]
  reg  _T_213; // @[package.scala 48:56:@1008.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@852.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@855.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@858.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@861.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@890.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@893.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@994.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1011.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@864.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@918.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@920.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@921.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@922.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@923.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@924.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@925.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@926.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@944.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@945.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@946.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@947.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@948.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@950.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@972.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@974.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@976.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@977.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@978.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@981.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@983.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@989.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@992.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1018.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@917.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@980.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@988.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@969.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@971.4]
  assign active_0_clock = clock; // @[:@853.4]
  assign active_0_reset = reset; // @[:@854.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@929.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@933.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@867.4]
  assign active_1_clock = clock; // @[:@856.4]
  assign active_1_reset = reset; // @[:@857.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@953.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@957.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@868.4]
  assign done_0_clock = clock; // @[:@859.4]
  assign done_0_reset = reset; // @[:@860.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@943.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@879.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@869.4]
  assign done_1_clock = clock; // @[:@862.4]
  assign done_1_reset = reset; // @[:@863.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@967.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@888.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@870.4]
  assign iterDone_0_clock = clock; // @[:@891.4]
  assign iterDone_0_reset = reset; // @[:@892.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@939.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@906.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@896.4]
  assign iterDone_1_clock = clock; // @[:@894.4]
  assign iterDone_1_reset = reset; // @[:@895.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@963.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@915.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@897.4]
  assign RetimeWrapper_clock = clock; // @[:@995.4]
  assign RetimeWrapper_reset = reset; // @[:@996.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@998.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@997.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1012.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1013.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1015.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1014.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x555_outr_UnitPipe_sm( // @[:@1435.2]
  input   clock, // @[:@1436.4]
  input   reset, // @[:@1437.4]
  input   io_enable, // @[:@1438.4]
  output  io_done, // @[:@1438.4]
  input   io_parentAck, // @[:@1438.4]
  input   io_doneIn_0, // @[:@1438.4]
  input   io_doneIn_1, // @[:@1438.4]
  output  io_enableOut_0, // @[:@1438.4]
  output  io_enableOut_1, // @[:@1438.4]
  output  io_childAck_0, // @[:@1438.4]
  output  io_childAck_1, // @[:@1438.4]
  input   io_ctrCopyDone_0, // @[:@1438.4]
  input   io_ctrCopyDone_1 // @[:@1438.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1441.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1444.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1447.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1450.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1482.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1688.4]
  wire  allDone; // @[Controllers.scala 80:47:@1453.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1507.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1508.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1509.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1510.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1511.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1514.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1516.4]
  wire  _T_148; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1531.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1532.4]
  wire  _T_160; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  wire  _T_178; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1563.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1564.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1576.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1577.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1578.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1579.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1580.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1583.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1585.4]
  wire  _T_216; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1600.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1601.4]
  wire  _T_228; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  wire  _T_246; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1632.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1633.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1649.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1651.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1653.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1658.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1660.4]
  wire  _T_282; // @[package.scala 100:49:@1666.4]
  reg  _T_285; // @[package.scala 48:56:@1667.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1669.4]
  reg  _T_299; // @[package.scala 48:56:@1685.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1441.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1444.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1447.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1450.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1479.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1482.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1523.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1537.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1555.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1592.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1606.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1624.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1671.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1688.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1453.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1507.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1508.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1509.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1510.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1511.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1514.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1516.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1531.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1532.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1563.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1564.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1576.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1577.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1578.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1579.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1580.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1583.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1585.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1600.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1601.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1632.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1633.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1649.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1651.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1653.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1658.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1660.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1666.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1669.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1695.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1657.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1665.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1646.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1648.4]
  assign active_0_clock = clock; // @[:@1442.4]
  assign active_0_reset = reset; // @[:@1443.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1518.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1522.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1456.4]
  assign active_1_clock = clock; // @[:@1445.4]
  assign active_1_reset = reset; // @[:@1446.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1587.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1591.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1457.4]
  assign done_0_clock = clock; // @[:@1448.4]
  assign done_0_reset = reset; // @[:@1449.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1568.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1468.4 Controllers.scala 170:32:@1575.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1458.4]
  assign done_1_clock = clock; // @[:@1451.4]
  assign done_1_reset = reset; // @[:@1452.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1637.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1477.4 Controllers.scala 170:32:@1644.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1459.4]
  assign iterDone_0_clock = clock; // @[:@1480.4]
  assign iterDone_0_reset = reset; // @[:@1481.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1536.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1495.4 Controllers.scala 168:36:@1552.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1485.4]
  assign iterDone_1_clock = clock; // @[:@1483.4]
  assign iterDone_1_reset = reset; // @[:@1484.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1605.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1504.4 Controllers.scala 168:36:@1621.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1486.4]
  assign RetimeWrapper_clock = clock; // @[:@1524.4]
  assign RetimeWrapper_reset = reset; // @[:@1525.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1527.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1526.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1538.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1539.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1541.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1540.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1556.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1557.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1559.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1558.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1593.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1594.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1596.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1595.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1607.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1608.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1610.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1609.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1625.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1626.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1628.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1627.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1672.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1673.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1675.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1674.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1689.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1690.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1692.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1691.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1924.2]
  input   clock, // @[:@1925.4]
  input   reset, // @[:@1926.4]
  input   io_input_inc_en_0, // @[:@1927.4]
  input   io_input_dinc_en_0, // @[:@1927.4]
  output  io_output_full // @[:@1927.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1929.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1930.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1931.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1932.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1932.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1933.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1934.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1935.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1935.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1936.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1937.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1930.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1931.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1932.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1932.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1933.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1934.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1935.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1935.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1936.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1937.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1951.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x292_fifoinraw_0( // @[:@2074.2]
  input   clock, // @[:@2075.4]
  input   reset // @[:@2076.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2121.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2121.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2122.4]
  assign elements_reset = reset; // @[:@2123.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 394:79:@2133.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2134.4]
endmodule
module x293_fifoinpacked_0( // @[:@2497.2]
  input   clock, // @[:@2498.4]
  input   reset, // @[:@2499.4]
  input   io_wPort_0_en_0, // @[:@2500.4]
  output  io_full, // @[:@2500.4]
  input   io_active_0_in, // @[:@2500.4]
  output  io_active_0_out // @[:@2500.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2544.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2544.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 439:39:@2618.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 437:129:@2616.4]
  assign elements_clock = clock; // @[:@2545.4]
  assign elements_reset = reset; // @[:@2546.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 394:79:@2556.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2557.4]
endmodule
module FF_7( // @[:@3047.2]
  input         clock, // @[:@3048.4]
  input         reset, // @[:@3049.4]
  output [12:0] io_rPort_0_output_0, // @[:@3050.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3050.4]
  input         io_wPort_0_reset, // @[:@3050.4]
  input         io_wPort_0_en_0 // @[:@3050.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 321:19:@3065.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 325:32:@3067.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 325:12:@3068.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@3067.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 325:12:@3068.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@3070.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3085.2]
  input         clock, // @[:@3086.4]
  input         reset, // @[:@3087.4]
  input         io_setup_saturate, // @[:@3088.4]
  input         io_input_reset, // @[:@3088.4]
  input         io_input_enable, // @[:@3088.4]
  output [12:0] io_output_count_0, // @[:@3088.4]
  output        io_output_oobs_0, // @[:@3088.4]
  output        io_output_done, // @[:@3088.4]
  output        io_output_saturated // @[:@3088.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3101.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3117.4]
  wire  _T_36; // @[Counter.scala 264:45:@3120.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3145.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3146.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3147.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3148.4]
  wire  _T_57; // @[Counter.scala 293:18:@3150.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3158.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3160.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3161.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3162.4]
  wire  _T_75; // @[Counter.scala 322:102:@3166.4]
  wire  _T_77; // @[Counter.scala 322:130:@3167.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3101.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3117.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3120.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3145.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3146.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3147.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3148.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3150.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3158.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3160.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3161.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3162.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3166.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3167.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3165.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3169.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3171.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3174.4]
  assign bases_0_clock = clock; // @[:@3102.4]
  assign bases_0_reset = reset; // @[:@3103.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3164.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3143.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3144.4]
  assign SRFF_clock = clock; // @[:@3118.4]
  assign SRFF_reset = reset; // @[:@3119.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3122.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3124.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3125.4]
endmodule
module SingleCounter_2( // @[:@3214.2]
  input         clock, // @[:@3215.4]
  input         reset, // @[:@3216.4]
  input         io_setup_saturate, // @[:@3217.4]
  input         io_input_reset, // @[:@3217.4]
  input         io_input_enable, // @[:@3217.4]
  output [12:0] io_output_count_0, // @[:@3217.4]
  output        io_output_oobs_0, // @[:@3217.4]
  output        io_output_done // @[:@3217.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3230.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3246.4]
  wire  _T_36; // @[Counter.scala 264:45:@3249.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3274.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3275.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3276.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3277.4]
  wire  _T_57; // @[Counter.scala 293:18:@3279.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3287.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3289.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3290.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3291.4]
  wire  _T_75; // @[Counter.scala 322:102:@3295.4]
  wire  _T_77; // @[Counter.scala 322:130:@3296.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3230.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3246.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3249.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3274.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh4); // @[Counter.scala 291:33:@3275.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh4); // @[Counter.scala 291:33:@3276.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3277.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3279.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3287.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3289.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3290.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3291.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3295.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3296.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3294.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3298.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3300.4]
  assign bases_0_clock = clock; // @[:@3231.4]
  assign bases_0_reset = reset; // @[:@3232.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3293.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3272.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3273.4]
  assign SRFF_clock = clock; // @[:@3247.4]
  assign SRFF_reset = reset; // @[:@3248.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3251.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3253.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3254.4]
endmodule
module x297_ctrchain( // @[:@3305.2]
  input         clock, // @[:@3306.4]
  input         reset, // @[:@3307.4]
  input         io_input_reset, // @[:@3308.4]
  input         io_input_enable, // @[:@3308.4]
  output [12:0] io_output_counts_1, // @[:@3308.4]
  output [12:0] io_output_counts_0, // @[:@3308.4]
  output        io_output_oobs_0, // @[:@3308.4]
  output        io_output_oobs_1, // @[:@3308.4]
  output        io_output_done // @[:@3308.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3310.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3313.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3313.4]
  wire  isDone; // @[Counter.scala 541:51:@3330.4]
  reg  wasDone; // @[Counter.scala 542:24:@3331.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3339.4]
  wire  _T_66; // @[Counter.scala 546:80:@3340.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3345.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3346.4]
  wire  _T_74; // @[Counter.scala 551:19:@3347.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3310.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3313.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3330.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3339.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3340.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3346.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3347.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3352.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3349.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3351.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3354.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3342.4]
  assign ctrs_0_clock = clock; // @[:@3311.4]
  assign ctrs_0_reset = reset; // @[:@3312.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3327.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3319.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3326.4]
  assign ctrs_1_clock = clock; // @[:@3314.4]
  assign ctrs_1_reset = reset; // @[:@3315.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3329.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3323.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3324.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3394.2]
  input   clock, // @[:@3395.4]
  input   reset, // @[:@3396.4]
  input   io_flow, // @[:@3397.4]
  input   io_in, // @[:@3397.4]
  output  io_out // @[:@3397.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@3399.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3412.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3411.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3410.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3409.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3408.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3406.4]
endmodule
module RetimeWrapper_25( // @[:@3522.2]
  input   clock, // @[:@3523.4]
  input   reset, // @[:@3524.4]
  input   io_flow, // @[:@3525.4]
  input   io_in, // @[:@3525.4]
  output  io_out // @[:@3525.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3527.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3540.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3539.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3538.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3537.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3536.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3534.4]
endmodule
module x323_inr_Foreach_sm( // @[:@3542.2]
  input   clock, // @[:@3543.4]
  input   reset, // @[:@3544.4]
  input   io_enable, // @[:@3545.4]
  output  io_done, // @[:@3545.4]
  output  io_doneLatch, // @[:@3545.4]
  input   io_ctrDone, // @[:@3545.4]
  output  io_datapathEn, // @[:@3545.4]
  output  io_ctrInc, // @[:@3545.4]
  output  io_ctrRst, // @[:@3545.4]
  input   io_parentAck, // @[:@3545.4]
  input   io_backpressure, // @[:@3545.4]
  input   io_break // @[:@3545.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3547.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3547.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3550.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3550.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3642.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3555.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3556.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3557.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3558.4]
  wire  _T_100; // @[package.scala 100:49:@3575.4]
  reg  _T_103; // @[package.scala 48:56:@3576.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  wire  _T_110; // @[package.scala 100:49:@3591.4]
  reg  _T_113; // @[package.scala 48:56:@3592.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3594.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3599.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3600.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3603.4]
  wire  _T_124; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  wire  _T_126; // @[package.scala 100:49:@3613.4]
  reg  _T_129; // @[package.scala 48:56:@3614.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3636.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3638.4]
  reg  _T_153; // @[package.scala 48:56:@3639.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3649.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3650.4]
  SRFF active ( // @[Controllers.scala 261:22:@3547.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3550.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3584.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3606.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3618.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3626.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3642.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3555.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3556.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3557.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3558.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3575.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3591.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3594.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3599.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3600.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3603.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3613.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3638.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3649.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3650.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3617.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3652.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3602.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3605.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3597.4]
  assign active_clock = clock; // @[:@3548.4]
  assign active_reset = reset; // @[:@3549.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3560.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3564.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3565.4]
  assign done_clock = clock; // @[:@3551.4]
  assign done_reset = reset; // @[:@3552.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3580.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3573.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3574.4]
  assign RetimeWrapper_clock = clock; // @[:@3585.4]
  assign RetimeWrapper_reset = reset; // @[:@3586.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3588.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3587.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3607.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3608.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3610.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3609.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3619.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3620.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3622.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3621.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3627.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3628.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3630.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3629.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3643.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3644.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3646.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3645.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@3759.2]
  input  [31:0] io_a, // @[:@3762.4]
  output [31:0] io_b // @[:@3762.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@3775.4]
endmodule
module _( // @[:@3777.2]
  input  [31:0] io_b, // @[:@3780.4]
  output [31:0] io_result // @[:@3780.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3785.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3785.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@3785.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3793.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3788.4]
endmodule
module fix2fixBox_2( // @[:@3831.2]
  input  [31:0] io_a, // @[:@3834.4]
  output [32:0] io_b // @[:@3834.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3844.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3844.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@3849.4]
endmodule
module __2( // @[:@3851.2]
  input  [31:0] io_b, // @[:@3854.4]
  output [32:0] io_result // @[:@3854.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3859.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3859.4]
  fix2fixBox_2 fix2fixBox ( // @[BigIPZynq.scala 219:30:@3859.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3867.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3862.4]
endmodule
module RetimeWrapper_29( // @[:@3919.2]
  input         clock, // @[:@3920.4]
  input         reset, // @[:@3921.4]
  input         io_flow, // @[:@3922.4]
  input  [31:0] io_in, // @[:@3922.4]
  output [31:0] io_out // @[:@3922.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3924.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3937.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3936.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3935.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3934.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3933.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3931.4]
endmodule
module fix2fixBox_4( // @[:@3939.2]
  input         clock, // @[:@3940.4]
  input         reset, // @[:@3941.4]
  input  [32:0] io_a, // @[:@3942.4]
  input         io_flow, // @[:@3942.4]
  output [31:0] io_b // @[:@3942.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3955.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3955.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3962.4]
  assign RetimeWrapper_clock = clock; // @[:@3956.4]
  assign RetimeWrapper_reset = reset; // @[:@3957.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3959.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3958.4]
endmodule
module x604_sub( // @[:@3964.2]
  input         clock, // @[:@3965.4]
  input         reset, // @[:@3966.4]
  input  [31:0] io_a, // @[:@3967.4]
  input  [31:0] io_b, // @[:@3967.4]
  input         io_flow, // @[:@3967.4]
  output [31:0] io_result // @[:@3967.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3975.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3975.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3982.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3982.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4001.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4001.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4001.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@3989.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@3990.4]
  __2 _ ( // @[Math.scala 720:24:@3975.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@3982.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@4001.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@3989.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@3990.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4009.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3978.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3985.4]
  assign fix2fixBox_clock = clock; // @[:@4002.4]
  assign fix2fixBox_reset = reset; // @[:@4003.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4004.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4007.4]
endmodule
module x303_sum( // @[:@4176.2]
  input         clock, // @[:@4177.4]
  input         reset, // @[:@4178.4]
  input  [31:0] io_a, // @[:@4179.4]
  input  [31:0] io_b, // @[:@4179.4]
  input         io_flow, // @[:@4179.4]
  output [31:0] io_result // @[:@4179.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4187.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@4187.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4194.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@4194.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4212.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4212.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4212.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4201.4]
  __2 _ ( // @[Math.scala 720:24:@4187.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@4194.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@4212.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4201.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4220.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@4190.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@4197.4]
  assign fix2fixBox_clock = clock; // @[:@4213.4]
  assign fix2fixBox_reset = reset; // @[:@4214.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4215.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4218.4]
endmodule
module x323_inr_Foreach_kernelx323_inr_Foreach_concrete1( // @[:@5894.2]
  input         clock, // @[:@5895.4]
  input         reset, // @[:@5896.4]
  output        io_in_x293_fifoinpacked_0_wPort_0_en_0, // @[:@5897.4]
  input         io_in_x293_fifoinpacked_0_full, // @[:@5897.4]
  output        io_in_x293_fifoinpacked_0_active_0_in, // @[:@5897.4]
  input         io_in_x293_fifoinpacked_0_active_0_out, // @[:@5897.4]
  input         io_sigsIn_backpressure, // @[:@5897.4]
  input         io_sigsIn_datapathEn, // @[:@5897.4]
  input         io_sigsIn_break, // @[:@5897.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@5897.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@5897.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@5897.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@5897.4]
  input         io_rr // @[:@5897.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@5931.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@5931.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@5943.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@5943.4]
  wire  x604_sub_1_clock; // @[Math.scala 191:24:@5970.4]
  wire  x604_sub_1_reset; // @[Math.scala 191:24:@5970.4]
  wire [31:0] x604_sub_1_io_a; // @[Math.scala 191:24:@5970.4]
  wire [31:0] x604_sub_1_io_b; // @[Math.scala 191:24:@5970.4]
  wire  x604_sub_1_io_flow; // @[Math.scala 191:24:@5970.4]
  wire [31:0] x604_sub_1_io_result; // @[Math.scala 191:24:@5970.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5980.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5980.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@5980.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@5980.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@5980.4]
  wire  x303_sum_1_clock; // @[Math.scala 150:24:@5989.4]
  wire  x303_sum_1_reset; // @[Math.scala 150:24:@5989.4]
  wire [31:0] x303_sum_1_io_a; // @[Math.scala 150:24:@5989.4]
  wire [31:0] x303_sum_1_io_b; // @[Math.scala 150:24:@5989.4]
  wire  x303_sum_1_io_flow; // @[Math.scala 150:24:@5989.4]
  wire [31:0] x303_sum_1_io_result; // @[Math.scala 150:24:@5989.4]
  wire  x304_sum_1_clock; // @[Math.scala 150:24:@6001.4]
  wire  x304_sum_1_reset; // @[Math.scala 150:24:@6001.4]
  wire [31:0] x304_sum_1_io_a; // @[Math.scala 150:24:@6001.4]
  wire [31:0] x304_sum_1_io_b; // @[Math.scala 150:24:@6001.4]
  wire  x304_sum_1_io_flow; // @[Math.scala 150:24:@6001.4]
  wire [31:0] x304_sum_1_io_result; // @[Math.scala 150:24:@6001.4]
  wire  x606_sum_1_clock; // @[Math.scala 150:24:@6016.4]
  wire  x606_sum_1_reset; // @[Math.scala 150:24:@6016.4]
  wire [31:0] x606_sum_1_io_a; // @[Math.scala 150:24:@6016.4]
  wire [31:0] x606_sum_1_io_b; // @[Math.scala 150:24:@6016.4]
  wire  x606_sum_1_io_flow; // @[Math.scala 150:24:@6016.4]
  wire [31:0] x606_sum_1_io_result; // @[Math.scala 150:24:@6016.4]
  wire [31:0] x307_1_io_b; // @[Math.scala 720:24:@6037.4]
  wire [31:0] x307_1_io_result; // @[Math.scala 720:24:@6037.4]
  wire  x308_sum_1_clock; // @[Math.scala 150:24:@6048.4]
  wire  x308_sum_1_reset; // @[Math.scala 150:24:@6048.4]
  wire [31:0] x308_sum_1_io_a; // @[Math.scala 150:24:@6048.4]
  wire [31:0] x308_sum_1_io_b; // @[Math.scala 150:24:@6048.4]
  wire  x308_sum_1_io_flow; // @[Math.scala 150:24:@6048.4]
  wire [31:0] x308_sum_1_io_result; // @[Math.scala 150:24:@6048.4]
  wire  x609_sum_1_clock; // @[Math.scala 150:24:@6063.4]
  wire  x609_sum_1_reset; // @[Math.scala 150:24:@6063.4]
  wire [31:0] x609_sum_1_io_a; // @[Math.scala 150:24:@6063.4]
  wire [31:0] x609_sum_1_io_b; // @[Math.scala 150:24:@6063.4]
  wire  x609_sum_1_io_flow; // @[Math.scala 150:24:@6063.4]
  wire [31:0] x609_sum_1_io_result; // @[Math.scala 150:24:@6063.4]
  wire [31:0] x311_1_io_b; // @[Math.scala 720:24:@6084.4]
  wire [31:0] x311_1_io_result; // @[Math.scala 720:24:@6084.4]
  wire  x312_sum_1_clock; // @[Math.scala 150:24:@6095.4]
  wire  x312_sum_1_reset; // @[Math.scala 150:24:@6095.4]
  wire [31:0] x312_sum_1_io_a; // @[Math.scala 150:24:@6095.4]
  wire [31:0] x312_sum_1_io_b; // @[Math.scala 150:24:@6095.4]
  wire  x312_sum_1_io_flow; // @[Math.scala 150:24:@6095.4]
  wire [31:0] x312_sum_1_io_result; // @[Math.scala 150:24:@6095.4]
  wire  x612_sum_1_clock; // @[Math.scala 150:24:@6110.4]
  wire  x612_sum_1_reset; // @[Math.scala 150:24:@6110.4]
  wire [31:0] x612_sum_1_io_a; // @[Math.scala 150:24:@6110.4]
  wire [31:0] x612_sum_1_io_b; // @[Math.scala 150:24:@6110.4]
  wire  x612_sum_1_io_flow; // @[Math.scala 150:24:@6110.4]
  wire [31:0] x612_sum_1_io_result; // @[Math.scala 150:24:@6110.4]
  wire [31:0] x315_1_io_b; // @[Math.scala 720:24:@6131.4]
  wire [31:0] x315_1_io_result; // @[Math.scala 720:24:@6131.4]
  wire  x316_sum_1_clock; // @[Math.scala 150:24:@6142.4]
  wire  x316_sum_1_reset; // @[Math.scala 150:24:@6142.4]
  wire [31:0] x316_sum_1_io_a; // @[Math.scala 150:24:@6142.4]
  wire [31:0] x316_sum_1_io_b; // @[Math.scala 150:24:@6142.4]
  wire  x316_sum_1_io_flow; // @[Math.scala 150:24:@6142.4]
  wire [31:0] x316_sum_1_io_result; // @[Math.scala 150:24:@6142.4]
  wire  x615_sum_1_clock; // @[Math.scala 150:24:@6157.4]
  wire  x615_sum_1_reset; // @[Math.scala 150:24:@6157.4]
  wire [31:0] x615_sum_1_io_a; // @[Math.scala 150:24:@6157.4]
  wire [31:0] x615_sum_1_io_b; // @[Math.scala 150:24:@6157.4]
  wire  x615_sum_1_io_flow; // @[Math.scala 150:24:@6157.4]
  wire [31:0] x615_sum_1_io_result; // @[Math.scala 150:24:@6157.4]
  wire [31:0] x319_1_io_b; // @[Math.scala 720:24:@6178.4]
  wire [31:0] x319_1_io_result; // @[Math.scala 720:24:@6178.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6197.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6197.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6197.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6197.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6197.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6206.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6206.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6206.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6206.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6206.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6217.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6217.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6217.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6217.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6217.4]
  wire  _T_327; // @[sm_x323_inr_Foreach.scala 62:18:@5956.4]
  wire  _T_328; // @[sm_x323_inr_Foreach.scala 62:55:@5957.4]
  wire [31:0] b298_number; // @[Math.scala 723:22:@5936.4 Math.scala 724:14:@5937.4]
  wire [42:0] _GEN_0; // @[Math.scala 461:32:@5961.4]
  wire [42:0] _T_331; // @[Math.scala 461:32:@5961.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@5966.4]
  wire [38:0] _T_334; // @[Math.scala 461:32:@5966.4]
  wire [31:0] x304_sum_number; // @[Math.scala 154:22:@6007.4 Math.scala 155:14:@6008.4]
  wire [33:0] _GEN_2; // @[Math.scala 461:32:@6012.4]
  wire [33:0] _T_353; // @[Math.scala 461:32:@6012.4]
  wire [31:0] x606_sum_number; // @[Math.scala 154:22:@6022.4 Math.scala 155:14:@6023.4]
  wire [31:0] _T_364; // @[Math.scala 406:49:@6029.4]
  wire [31:0] _T_366; // @[Math.scala 406:56:@6031.4]
  wire [31:0] _T_367; // @[Math.scala 406:56:@6032.4]
  wire [31:0] x308_sum_number; // @[Math.scala 154:22:@6054.4 Math.scala 155:14:@6055.4]
  wire [33:0] _GEN_3; // @[Math.scala 461:32:@6059.4]
  wire [33:0] _T_381; // @[Math.scala 461:32:@6059.4]
  wire [31:0] x609_sum_number; // @[Math.scala 154:22:@6069.4 Math.scala 155:14:@6070.4]
  wire [31:0] _T_392; // @[Math.scala 406:49:@6076.4]
  wire [31:0] _T_394; // @[Math.scala 406:56:@6078.4]
  wire [31:0] _T_395; // @[Math.scala 406:56:@6079.4]
  wire [31:0] x312_sum_number; // @[Math.scala 154:22:@6101.4 Math.scala 155:14:@6102.4]
  wire [33:0] _GEN_4; // @[Math.scala 461:32:@6106.4]
  wire [33:0] _T_409; // @[Math.scala 461:32:@6106.4]
  wire [31:0] x612_sum_number; // @[Math.scala 154:22:@6116.4 Math.scala 155:14:@6117.4]
  wire [31:0] _T_420; // @[Math.scala 406:49:@6123.4]
  wire [31:0] _T_422; // @[Math.scala 406:56:@6125.4]
  wire [31:0] _T_423; // @[Math.scala 406:56:@6126.4]
  wire [31:0] x316_sum_number; // @[Math.scala 154:22:@6148.4 Math.scala 155:14:@6149.4]
  wire [33:0] _GEN_5; // @[Math.scala 461:32:@6153.4]
  wire [33:0] _T_437; // @[Math.scala 461:32:@6153.4]
  wire [31:0] x615_sum_number; // @[Math.scala 154:22:@6163.4 Math.scala 155:14:@6164.4]
  wire [31:0] _T_448; // @[Math.scala 406:49:@6170.4]
  wire [31:0] _T_450; // @[Math.scala 406:56:@6172.4]
  wire [31:0] _T_451; // @[Math.scala 406:56:@6173.4]
  wire  _T_475; // @[sm_x323_inr_Foreach.scala 123:131:@6214.4]
  wire  _T_479; // @[package.scala 96:25:@6222.4 package.scala 96:25:@6223.4]
  wire  _T_481; // @[implicits.scala 55:10:@6224.4]
  wire  _T_482; // @[sm_x323_inr_Foreach.scala 123:148:@6225.4]
  wire  _T_484; // @[sm_x323_inr_Foreach.scala 123:236:@6227.4]
  wire  _T_485; // @[sm_x323_inr_Foreach.scala 123:255:@6228.4]
  wire  x635_b300_D4; // @[package.scala 96:25:@6202.4 package.scala 96:25:@6203.4]
  wire  _T_488; // @[sm_x323_inr_Foreach.scala 123:291:@6230.4]
  wire  x636_b301_D4; // @[package.scala 96:25:@6211.4 package.scala 96:25:@6212.4]
  _ _ ( // @[Math.scala 720:24:@5931.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@5943.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x604_sub x604_sub_1 ( // @[Math.scala 191:24:@5970.4]
    .clock(x604_sub_1_clock),
    .reset(x604_sub_1_reset),
    .io_a(x604_sub_1_io_a),
    .io_b(x604_sub_1_io_b),
    .io_flow(x604_sub_1_io_flow),
    .io_result(x604_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@5980.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x303_sum x303_sum_1 ( // @[Math.scala 150:24:@5989.4]
    .clock(x303_sum_1_clock),
    .reset(x303_sum_1_reset),
    .io_a(x303_sum_1_io_a),
    .io_b(x303_sum_1_io_b),
    .io_flow(x303_sum_1_io_flow),
    .io_result(x303_sum_1_io_result)
  );
  x303_sum x304_sum_1 ( // @[Math.scala 150:24:@6001.4]
    .clock(x304_sum_1_clock),
    .reset(x304_sum_1_reset),
    .io_a(x304_sum_1_io_a),
    .io_b(x304_sum_1_io_b),
    .io_flow(x304_sum_1_io_flow),
    .io_result(x304_sum_1_io_result)
  );
  x303_sum x606_sum_1 ( // @[Math.scala 150:24:@6016.4]
    .clock(x606_sum_1_clock),
    .reset(x606_sum_1_reset),
    .io_a(x606_sum_1_io_a),
    .io_b(x606_sum_1_io_b),
    .io_flow(x606_sum_1_io_flow),
    .io_result(x606_sum_1_io_result)
  );
  _ x307_1 ( // @[Math.scala 720:24:@6037.4]
    .io_b(x307_1_io_b),
    .io_result(x307_1_io_result)
  );
  x303_sum x308_sum_1 ( // @[Math.scala 150:24:@6048.4]
    .clock(x308_sum_1_clock),
    .reset(x308_sum_1_reset),
    .io_a(x308_sum_1_io_a),
    .io_b(x308_sum_1_io_b),
    .io_flow(x308_sum_1_io_flow),
    .io_result(x308_sum_1_io_result)
  );
  x303_sum x609_sum_1 ( // @[Math.scala 150:24:@6063.4]
    .clock(x609_sum_1_clock),
    .reset(x609_sum_1_reset),
    .io_a(x609_sum_1_io_a),
    .io_b(x609_sum_1_io_b),
    .io_flow(x609_sum_1_io_flow),
    .io_result(x609_sum_1_io_result)
  );
  _ x311_1 ( // @[Math.scala 720:24:@6084.4]
    .io_b(x311_1_io_b),
    .io_result(x311_1_io_result)
  );
  x303_sum x312_sum_1 ( // @[Math.scala 150:24:@6095.4]
    .clock(x312_sum_1_clock),
    .reset(x312_sum_1_reset),
    .io_a(x312_sum_1_io_a),
    .io_b(x312_sum_1_io_b),
    .io_flow(x312_sum_1_io_flow),
    .io_result(x312_sum_1_io_result)
  );
  x303_sum x612_sum_1 ( // @[Math.scala 150:24:@6110.4]
    .clock(x612_sum_1_clock),
    .reset(x612_sum_1_reset),
    .io_a(x612_sum_1_io_a),
    .io_b(x612_sum_1_io_b),
    .io_flow(x612_sum_1_io_flow),
    .io_result(x612_sum_1_io_result)
  );
  _ x315_1 ( // @[Math.scala 720:24:@6131.4]
    .io_b(x315_1_io_b),
    .io_result(x315_1_io_result)
  );
  x303_sum x316_sum_1 ( // @[Math.scala 150:24:@6142.4]
    .clock(x316_sum_1_clock),
    .reset(x316_sum_1_reset),
    .io_a(x316_sum_1_io_a),
    .io_b(x316_sum_1_io_b),
    .io_flow(x316_sum_1_io_flow),
    .io_result(x316_sum_1_io_result)
  );
  x303_sum x615_sum_1 ( // @[Math.scala 150:24:@6157.4]
    .clock(x615_sum_1_clock),
    .reset(x615_sum_1_reset),
    .io_a(x615_sum_1_io_a),
    .io_b(x615_sum_1_io_b),
    .io_flow(x615_sum_1_io_flow),
    .io_result(x615_sum_1_io_result)
  );
  _ x319_1 ( // @[Math.scala 720:24:@6178.4]
    .io_b(x319_1_io_b),
    .io_result(x319_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@6197.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@6206.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@6217.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_327 = ~ io_in_x293_fifoinpacked_0_full; // @[sm_x323_inr_Foreach.scala 62:18:@5956.4]
  assign _T_328 = ~ io_in_x293_fifoinpacked_0_active_0_out; // @[sm_x323_inr_Foreach.scala 62:55:@5957.4]
  assign b298_number = __io_result; // @[Math.scala 723:22:@5936.4 Math.scala 724:14:@5937.4]
  assign _GEN_0 = {{11'd0}, b298_number}; // @[Math.scala 461:32:@5961.4]
  assign _T_331 = _GEN_0 << 11; // @[Math.scala 461:32:@5961.4]
  assign _GEN_1 = {{7'd0}, b298_number}; // @[Math.scala 461:32:@5966.4]
  assign _T_334 = _GEN_1 << 7; // @[Math.scala 461:32:@5966.4]
  assign x304_sum_number = x304_sum_1_io_result; // @[Math.scala 154:22:@6007.4 Math.scala 155:14:@6008.4]
  assign _GEN_2 = {{2'd0}, x304_sum_number}; // @[Math.scala 461:32:@6012.4]
  assign _T_353 = _GEN_2 << 2; // @[Math.scala 461:32:@6012.4]
  assign x606_sum_number = x606_sum_1_io_result; // @[Math.scala 154:22:@6022.4 Math.scala 155:14:@6023.4]
  assign _T_364 = $signed(x606_sum_number); // @[Math.scala 406:49:@6029.4]
  assign _T_366 = $signed(_T_364) & $signed(32'shff); // @[Math.scala 406:56:@6031.4]
  assign _T_367 = $signed(_T_366); // @[Math.scala 406:56:@6032.4]
  assign x308_sum_number = x308_sum_1_io_result; // @[Math.scala 154:22:@6054.4 Math.scala 155:14:@6055.4]
  assign _GEN_3 = {{2'd0}, x308_sum_number}; // @[Math.scala 461:32:@6059.4]
  assign _T_381 = _GEN_3 << 2; // @[Math.scala 461:32:@6059.4]
  assign x609_sum_number = x609_sum_1_io_result; // @[Math.scala 154:22:@6069.4 Math.scala 155:14:@6070.4]
  assign _T_392 = $signed(x609_sum_number); // @[Math.scala 406:49:@6076.4]
  assign _T_394 = $signed(_T_392) & $signed(32'shff); // @[Math.scala 406:56:@6078.4]
  assign _T_395 = $signed(_T_394); // @[Math.scala 406:56:@6079.4]
  assign x312_sum_number = x312_sum_1_io_result; // @[Math.scala 154:22:@6101.4 Math.scala 155:14:@6102.4]
  assign _GEN_4 = {{2'd0}, x312_sum_number}; // @[Math.scala 461:32:@6106.4]
  assign _T_409 = _GEN_4 << 2; // @[Math.scala 461:32:@6106.4]
  assign x612_sum_number = x612_sum_1_io_result; // @[Math.scala 154:22:@6116.4 Math.scala 155:14:@6117.4]
  assign _T_420 = $signed(x612_sum_number); // @[Math.scala 406:49:@6123.4]
  assign _T_422 = $signed(_T_420) & $signed(32'shff); // @[Math.scala 406:56:@6125.4]
  assign _T_423 = $signed(_T_422); // @[Math.scala 406:56:@6126.4]
  assign x316_sum_number = x316_sum_1_io_result; // @[Math.scala 154:22:@6148.4 Math.scala 155:14:@6149.4]
  assign _GEN_5 = {{2'd0}, x316_sum_number}; // @[Math.scala 461:32:@6153.4]
  assign _T_437 = _GEN_5 << 2; // @[Math.scala 461:32:@6153.4]
  assign x615_sum_number = x615_sum_1_io_result; // @[Math.scala 154:22:@6163.4 Math.scala 155:14:@6164.4]
  assign _T_448 = $signed(x615_sum_number); // @[Math.scala 406:49:@6170.4]
  assign _T_450 = $signed(_T_448) & $signed(32'shff); // @[Math.scala 406:56:@6172.4]
  assign _T_451 = $signed(_T_450); // @[Math.scala 406:56:@6173.4]
  assign _T_475 = ~ io_sigsIn_break; // @[sm_x323_inr_Foreach.scala 123:131:@6214.4]
  assign _T_479 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@6222.4 package.scala 96:25:@6223.4]
  assign _T_481 = io_rr ? _T_479 : 1'h0; // @[implicits.scala 55:10:@6224.4]
  assign _T_482 = _T_475 & _T_481; // @[sm_x323_inr_Foreach.scala 123:148:@6225.4]
  assign _T_484 = _T_482 & _T_475; // @[sm_x323_inr_Foreach.scala 123:236:@6227.4]
  assign _T_485 = _T_484 & io_sigsIn_backpressure; // @[sm_x323_inr_Foreach.scala 123:255:@6228.4]
  assign x635_b300_D4 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6202.4 package.scala 96:25:@6203.4]
  assign _T_488 = _T_485 & x635_b300_D4; // @[sm_x323_inr_Foreach.scala 123:291:@6230.4]
  assign x636_b301_D4 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@6211.4 package.scala 96:25:@6212.4]
  assign io_in_x293_fifoinpacked_0_wPort_0_en_0 = _T_488 & x636_b301_D4; // @[MemInterfaceType.scala 93:57:@6234.4]
  assign io_in_x293_fifoinpacked_0_active_0_in = x635_b300_D4 & x636_b301_D4; // @[MemInterfaceType.scala 147:18:@6237.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@5934.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@5946.4]
  assign x604_sub_1_clock = clock; // @[:@5971.4]
  assign x604_sub_1_reset = reset; // @[:@5972.4]
  assign x604_sub_1_io_a = _T_331[31:0]; // @[Math.scala 192:17:@5973.4]
  assign x604_sub_1_io_b = _T_334[31:0]; // @[Math.scala 193:17:@5974.4]
  assign x604_sub_1_io_flow = _T_327 | _T_328; // @[Math.scala 194:20:@5975.4]
  assign RetimeWrapper_clock = clock; // @[:@5981.4]
  assign RetimeWrapper_reset = reset; // @[:@5982.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5984.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@5983.4]
  assign x303_sum_1_clock = clock; // @[:@5990.4]
  assign x303_sum_1_reset = reset; // @[:@5991.4]
  assign x303_sum_1_io_a = x604_sub_1_io_result; // @[Math.scala 151:17:@5992.4]
  assign x303_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@5993.4]
  assign x303_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5994.4]
  assign x304_sum_1_clock = clock; // @[:@6002.4]
  assign x304_sum_1_reset = reset; // @[:@6003.4]
  assign x304_sum_1_io_a = x303_sum_1_io_result; // @[Math.scala 151:17:@6004.4]
  assign x304_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@6005.4]
  assign x304_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6006.4]
  assign x606_sum_1_clock = clock; // @[:@6017.4]
  assign x606_sum_1_reset = reset; // @[:@6018.4]
  assign x606_sum_1_io_a = _T_353[31:0]; // @[Math.scala 151:17:@6019.4]
  assign x606_sum_1_io_b = x304_sum_1_io_result; // @[Math.scala 152:17:@6020.4]
  assign x606_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6021.4]
  assign x307_1_io_b = $unsigned(_T_367); // @[Math.scala 721:17:@6040.4]
  assign x308_sum_1_clock = clock; // @[:@6049.4]
  assign x308_sum_1_reset = reset; // @[:@6050.4]
  assign x308_sum_1_io_a = x303_sum_1_io_result; // @[Math.scala 151:17:@6051.4]
  assign x308_sum_1_io_b = 32'h2; // @[Math.scala 152:17:@6052.4]
  assign x308_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6053.4]
  assign x609_sum_1_clock = clock; // @[:@6064.4]
  assign x609_sum_1_reset = reset; // @[:@6065.4]
  assign x609_sum_1_io_a = _T_381[31:0]; // @[Math.scala 151:17:@6066.4]
  assign x609_sum_1_io_b = x308_sum_1_io_result; // @[Math.scala 152:17:@6067.4]
  assign x609_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6068.4]
  assign x311_1_io_b = $unsigned(_T_395); // @[Math.scala 721:17:@6087.4]
  assign x312_sum_1_clock = clock; // @[:@6096.4]
  assign x312_sum_1_reset = reset; // @[:@6097.4]
  assign x312_sum_1_io_a = x303_sum_1_io_result; // @[Math.scala 151:17:@6098.4]
  assign x312_sum_1_io_b = 32'h3; // @[Math.scala 152:17:@6099.4]
  assign x312_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6100.4]
  assign x612_sum_1_clock = clock; // @[:@6111.4]
  assign x612_sum_1_reset = reset; // @[:@6112.4]
  assign x612_sum_1_io_a = _T_409[31:0]; // @[Math.scala 151:17:@6113.4]
  assign x612_sum_1_io_b = x312_sum_1_io_result; // @[Math.scala 152:17:@6114.4]
  assign x612_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6115.4]
  assign x315_1_io_b = $unsigned(_T_423); // @[Math.scala 721:17:@6134.4]
  assign x316_sum_1_clock = clock; // @[:@6143.4]
  assign x316_sum_1_reset = reset; // @[:@6144.4]
  assign x316_sum_1_io_a = x303_sum_1_io_result; // @[Math.scala 151:17:@6145.4]
  assign x316_sum_1_io_b = 32'h4; // @[Math.scala 152:17:@6146.4]
  assign x316_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6147.4]
  assign x615_sum_1_clock = clock; // @[:@6158.4]
  assign x615_sum_1_reset = reset; // @[:@6159.4]
  assign x615_sum_1_io_a = _T_437[31:0]; // @[Math.scala 151:17:@6160.4]
  assign x615_sum_1_io_b = x316_sum_1_io_result; // @[Math.scala 152:17:@6161.4]
  assign x615_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@6162.4]
  assign x319_1_io_b = $unsigned(_T_451); // @[Math.scala 721:17:@6181.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6198.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6199.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@6201.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@6200.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6207.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6208.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@6210.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@6209.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6218.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6219.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@6221.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@6220.4]
endmodule
module RetimeWrapper_48( // @[:@7355.2]
  input   clock, // @[:@7356.4]
  input   reset, // @[:@7357.4]
  input   io_flow, // @[:@7358.4]
  input   io_in, // @[:@7358.4]
  output  io_out // @[:@7358.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@7360.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@7360.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@7360.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7360.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7360.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7360.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(70)) sr ( // @[RetimeShiftRegister.scala 15:20:@7360.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7373.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7372.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@7371.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7370.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7369.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7367.4]
endmodule
module RetimeWrapper_52( // @[:@7483.2]
  input   clock, // @[:@7484.4]
  input   reset, // @[:@7485.4]
  input   io_flow, // @[:@7486.4]
  input   io_in, // @[:@7486.4]
  output  io_out // @[:@7486.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@7488.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@7488.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@7488.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7488.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7488.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7488.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(69)) sr ( // @[RetimeShiftRegister.scala 15:20:@7488.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7501.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7500.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@7499.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7498.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7497.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7495.4]
endmodule
module x553_inr_Foreach_SAMPLER_BOX_sm( // @[:@7503.2]
  input   clock, // @[:@7504.4]
  input   reset, // @[:@7505.4]
  input   io_enable, // @[:@7506.4]
  output  io_done, // @[:@7506.4]
  output  io_doneLatch, // @[:@7506.4]
  input   io_ctrDone, // @[:@7506.4]
  output  io_datapathEn, // @[:@7506.4]
  output  io_ctrInc, // @[:@7506.4]
  output  io_ctrRst, // @[:@7506.4]
  input   io_parentAck, // @[:@7506.4]
  input   io_backpressure, // @[:@7506.4]
  input   io_break // @[:@7506.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@7508.4]
  wire  active_reset; // @[Controllers.scala 261:22:@7508.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@7508.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@7508.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@7508.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@7508.4]
  wire  done_clock; // @[Controllers.scala 262:20:@7511.4]
  wire  done_reset; // @[Controllers.scala 262:20:@7511.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@7511.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@7511.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@7511.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@7511.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7545.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7545.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@7545.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@7545.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@7545.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@7567.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@7567.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@7567.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@7567.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@7567.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@7579.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@7579.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@7579.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@7579.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@7579.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@7587.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@7587.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@7587.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@7587.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@7587.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@7603.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@7603.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@7603.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@7603.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@7603.4]
  wire  _T_80; // @[Controllers.scala 264:48:@7516.4]
  wire  _T_81; // @[Controllers.scala 264:46:@7517.4]
  wire  _T_82; // @[Controllers.scala 264:62:@7518.4]
  wire  _T_83; // @[Controllers.scala 264:60:@7519.4]
  wire  _T_100; // @[package.scala 100:49:@7536.4]
  reg  _T_103; // @[package.scala 48:56:@7537.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@7550.4 package.scala 96:25:@7551.4]
  wire  _T_110; // @[package.scala 100:49:@7552.4]
  reg  _T_113; // @[package.scala 48:56:@7553.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@7555.4]
  wire  _T_118; // @[Controllers.scala 283:41:@7560.4]
  wire  _T_119; // @[Controllers.scala 283:59:@7561.4]
  wire  _T_121; // @[Controllers.scala 284:37:@7564.4]
  wire  _T_124; // @[package.scala 96:25:@7572.4 package.scala 96:25:@7573.4]
  wire  _T_126; // @[package.scala 100:49:@7574.4]
  reg  _T_129; // @[package.scala 48:56:@7575.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@7597.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@7599.4]
  reg  _T_153; // @[package.scala 48:56:@7600.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@7608.4 package.scala 96:25:@7609.4]
  wire  _T_158; // @[Controllers.scala 292:61:@7610.4]
  wire  _T_159; // @[Controllers.scala 292:24:@7611.4]
  SRFF active ( // @[Controllers.scala 261:22:@7508.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@7511.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_48 RetimeWrapper ( // @[package.scala 93:22:@7545.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_1 ( // @[package.scala 93:22:@7567.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@7579.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@7587.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_4 ( // @[package.scala 93:22:@7603.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@7516.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@7517.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@7518.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@7519.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@7536.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@7550.4 package.scala 96:25:@7551.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@7552.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@7555.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@7560.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@7561.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@7564.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@7572.4 package.scala 96:25:@7573.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@7574.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@7599.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@7608.4 package.scala 96:25:@7609.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@7610.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@7611.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@7578.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@7613.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@7563.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@7566.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@7558.4]
  assign active_clock = clock; // @[:@7509.4]
  assign active_reset = reset; // @[:@7510.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@7521.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@7525.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@7526.4]
  assign done_clock = clock; // @[:@7512.4]
  assign done_reset = reset; // @[:@7513.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@7541.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@7534.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@7535.4]
  assign RetimeWrapper_clock = clock; // @[:@7546.4]
  assign RetimeWrapper_reset = reset; // @[:@7547.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@7549.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@7548.4]
  assign RetimeWrapper_1_clock = clock; // @[:@7568.4]
  assign RetimeWrapper_1_reset = reset; // @[:@7569.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@7571.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@7570.4]
  assign RetimeWrapper_2_clock = clock; // @[:@7580.4]
  assign RetimeWrapper_2_reset = reset; // @[:@7581.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@7583.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@7582.4]
  assign RetimeWrapper_3_clock = clock; // @[:@7588.4]
  assign RetimeWrapper_3_reset = reset; // @[:@7589.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@7591.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@7590.4]
  assign RetimeWrapper_4_clock = clock; // @[:@7604.4]
  assign RetimeWrapper_4_reset = reset; // @[:@7605.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@7607.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@7606.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module RetimeWrapper_56( // @[:@7804.2]
  input          clock, // @[:@7805.4]
  input          reset, // @[:@7806.4]
  input          io_flow, // @[:@7807.4]
  input  [127:0] io_in, // @[:@7807.4]
  output [127:0] io_out // @[:@7807.4]
);
  wire [127:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@7809.4]
  wire [127:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@7809.4]
  wire [127:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@7809.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7809.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7809.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7809.4]
  RetimeShiftRegister #(.WIDTH(128), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@7809.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7822.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7821.4]
  assign sr_init = 128'h0; // @[RetimeShiftRegister.scala 19:16:@7820.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7819.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7818.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7816.4]
endmodule
module SRAM_1( // @[:@7840.2]
  input         clock, // @[:@7841.4]
  input         reset, // @[:@7842.4]
  input  [8:0]  io_raddr, // @[:@7843.4]
  input         io_wen, // @[:@7843.4]
  input  [8:0]  io_waddr, // @[:@7843.4]
  input  [31:0] io_wdata, // @[:@7843.4]
  output [31:0] io_rdata, // @[:@7843.4]
  input         io_backpressure // @[:@7843.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@7845.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@7845.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@7845.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@7845.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@7845.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@7845.4]
  wire [8:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@7845.4]
  wire [8:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@7845.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@7845.4]
  wire  _T_19; // @[SRAM.scala 182:49:@7863.4]
  wire  _T_20; // @[SRAM.scala 182:37:@7864.4]
  reg  _T_23; // @[SRAM.scala 182:29:@7865.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@7867.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(320), .AWIDTH(9)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@7845.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@7863.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@7864.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@7872.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@7859.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@7860.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@7857.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@7862.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@7861.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@7858.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@7856.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@7855.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_57( // @[:@7886.2]
  input        clock, // @[:@7887.4]
  input        reset, // @[:@7888.4]
  input        io_flow, // @[:@7889.4]
  input  [8:0] io_in, // @[:@7889.4]
  output [8:0] io_out // @[:@7889.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@7891.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@7891.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@7891.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7891.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7891.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7891.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@7891.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7904.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7903.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@7902.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7901.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7900.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7898.4]
endmodule
module Mem1D_5( // @[:@7906.2]
  input         clock, // @[:@7907.4]
  input         reset, // @[:@7908.4]
  input  [8:0]  io_r_ofs_0, // @[:@7909.4]
  input         io_r_backpressure, // @[:@7909.4]
  input  [8:0]  io_w_ofs_0, // @[:@7909.4]
  input  [31:0] io_w_data_0, // @[:@7909.4]
  input         io_w_en_0, // @[:@7909.4]
  output [31:0] io_output // @[:@7909.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@7913.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 715:21:@7913.4]
  wire [8:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@7913.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 715:21:@7913.4]
  wire [8:0] SRAM_io_waddr; // @[MemPrimitives.scala 715:21:@7913.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 715:21:@7913.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@7913.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@7913.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7916.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7916.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@7916.4]
  wire [8:0] RetimeWrapper_io_in; // @[package.scala 93:22:@7916.4]
  wire [8:0] RetimeWrapper_io_out; // @[package.scala 93:22:@7916.4]
  wire  wInBound; // @[MemPrimitives.scala 702:32:@7911.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 715:21:@7913.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_57 RetimeWrapper ( // @[package.scala 93:22:@7916.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 9'h140; // @[MemPrimitives.scala 702:32:@7911.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@7929.4]
  assign SRAM_clock = clock; // @[:@7914.4]
  assign SRAM_reset = reset; // @[:@7915.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@7923.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 719:22:@7926.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 718:22:@7924.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 720:22:@7927.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@7928.4]
  assign RetimeWrapper_clock = clock; // @[:@7917.4]
  assign RetimeWrapper_reset = reset; // @[:@7918.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@7920.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@7919.4]
endmodule
module StickySelects_1( // @[:@10392.2]
  input   clock, // @[:@10393.4]
  input   reset, // @[:@10394.4]
  input   io_ins_0, // @[:@10395.4]
  input   io_ins_1, // @[:@10395.4]
  input   io_ins_2, // @[:@10395.4]
  input   io_ins_3, // @[:@10395.4]
  input   io_ins_4, // @[:@10395.4]
  input   io_ins_5, // @[:@10395.4]
  input   io_ins_6, // @[:@10395.4]
  input   io_ins_7, // @[:@10395.4]
  input   io_ins_8, // @[:@10395.4]
  output  io_outs_0, // @[:@10395.4]
  output  io_outs_1, // @[:@10395.4]
  output  io_outs_2, // @[:@10395.4]
  output  io_outs_3, // @[:@10395.4]
  output  io_outs_4, // @[:@10395.4]
  output  io_outs_5, // @[:@10395.4]
  output  io_outs_6, // @[:@10395.4]
  output  io_outs_7, // @[:@10395.4]
  output  io_outs_8 // @[:@10395.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@10397.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@10398.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@10399.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@10400.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@10401.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@10402.4]
  reg [31:0] _RAND_5;
  reg  _T_37; // @[StickySelects.scala 37:46:@10403.4]
  reg [31:0] _RAND_6;
  reg  _T_40; // @[StickySelects.scala 37:46:@10404.4]
  reg [31:0] _RAND_7;
  reg  _T_43; // @[StickySelects.scala 37:46:@10405.4]
  reg [31:0] _RAND_8;
  wire  _T_44; // @[StickySelects.scala 47:46:@10406.4]
  wire  _T_45; // @[StickySelects.scala 47:46:@10407.4]
  wire  _T_46; // @[StickySelects.scala 47:46:@10408.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@10409.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@10410.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@10411.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@10412.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@10413.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@10414.4]
  wire  _T_53; // @[StickySelects.scala 47:46:@10416.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@10417.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@10418.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@10419.4]
  wire  _T_57; // @[StickySelects.scala 47:46:@10420.4]
  wire  _T_58; // @[StickySelects.scala 47:46:@10421.4]
  wire  _T_59; // @[StickySelects.scala 47:46:@10422.4]
  wire  _T_60; // @[StickySelects.scala 49:53:@10423.4]
  wire  _T_61; // @[StickySelects.scala 49:21:@10424.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@10426.4]
  wire  _T_63; // @[StickySelects.scala 47:46:@10427.4]
  wire  _T_64; // @[StickySelects.scala 47:46:@10428.4]
  wire  _T_65; // @[StickySelects.scala 47:46:@10429.4]
  wire  _T_66; // @[StickySelects.scala 47:46:@10430.4]
  wire  _T_67; // @[StickySelects.scala 47:46:@10431.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@10432.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@10433.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@10434.4]
  wire  _T_72; // @[StickySelects.scala 47:46:@10437.4]
  wire  _T_73; // @[StickySelects.scala 47:46:@10438.4]
  wire  _T_74; // @[StickySelects.scala 47:46:@10439.4]
  wire  _T_75; // @[StickySelects.scala 47:46:@10440.4]
  wire  _T_76; // @[StickySelects.scala 47:46:@10441.4]
  wire  _T_77; // @[StickySelects.scala 47:46:@10442.4]
  wire  _T_78; // @[StickySelects.scala 49:53:@10443.4]
  wire  _T_79; // @[StickySelects.scala 49:21:@10444.4]
  wire  _T_82; // @[StickySelects.scala 47:46:@10448.4]
  wire  _T_83; // @[StickySelects.scala 47:46:@10449.4]
  wire  _T_84; // @[StickySelects.scala 47:46:@10450.4]
  wire  _T_85; // @[StickySelects.scala 47:46:@10451.4]
  wire  _T_86; // @[StickySelects.scala 47:46:@10452.4]
  wire  _T_87; // @[StickySelects.scala 49:53:@10453.4]
  wire  _T_88; // @[StickySelects.scala 49:21:@10454.4]
  wire  _T_92; // @[StickySelects.scala 47:46:@10459.4]
  wire  _T_93; // @[StickySelects.scala 47:46:@10460.4]
  wire  _T_94; // @[StickySelects.scala 47:46:@10461.4]
  wire  _T_95; // @[StickySelects.scala 47:46:@10462.4]
  wire  _T_96; // @[StickySelects.scala 49:53:@10463.4]
  wire  _T_97; // @[StickySelects.scala 49:21:@10464.4]
  wire  _T_102; // @[StickySelects.scala 47:46:@10470.4]
  wire  _T_103; // @[StickySelects.scala 47:46:@10471.4]
  wire  _T_104; // @[StickySelects.scala 47:46:@10472.4]
  wire  _T_105; // @[StickySelects.scala 49:53:@10473.4]
  wire  _T_106; // @[StickySelects.scala 49:21:@10474.4]
  wire  _T_112; // @[StickySelects.scala 47:46:@10481.4]
  wire  _T_113; // @[StickySelects.scala 47:46:@10482.4]
  wire  _T_114; // @[StickySelects.scala 49:53:@10483.4]
  wire  _T_115; // @[StickySelects.scala 49:21:@10484.4]
  wire  _T_122; // @[StickySelects.scala 47:46:@10492.4]
  wire  _T_123; // @[StickySelects.scala 49:53:@10493.4]
  wire  _T_124; // @[StickySelects.scala 49:21:@10494.4]
  assign _T_44 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@10406.4]
  assign _T_45 = _T_44 | io_ins_3; // @[StickySelects.scala 47:46:@10407.4]
  assign _T_46 = _T_45 | io_ins_4; // @[StickySelects.scala 47:46:@10408.4]
  assign _T_47 = _T_46 | io_ins_5; // @[StickySelects.scala 47:46:@10409.4]
  assign _T_48 = _T_47 | io_ins_6; // @[StickySelects.scala 47:46:@10410.4]
  assign _T_49 = _T_48 | io_ins_7; // @[StickySelects.scala 47:46:@10411.4]
  assign _T_50 = _T_49 | io_ins_8; // @[StickySelects.scala 47:46:@10412.4]
  assign _T_51 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@10413.4]
  assign _T_52 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 49:21:@10414.4]
  assign _T_53 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@10416.4]
  assign _T_54 = _T_53 | io_ins_3; // @[StickySelects.scala 47:46:@10417.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@10418.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@10419.4]
  assign _T_57 = _T_56 | io_ins_6; // @[StickySelects.scala 47:46:@10420.4]
  assign _T_58 = _T_57 | io_ins_7; // @[StickySelects.scala 47:46:@10421.4]
  assign _T_59 = _T_58 | io_ins_8; // @[StickySelects.scala 47:46:@10422.4]
  assign _T_60 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@10423.4]
  assign _T_61 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 49:21:@10424.4]
  assign _T_62 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@10426.4]
  assign _T_63 = _T_62 | io_ins_3; // @[StickySelects.scala 47:46:@10427.4]
  assign _T_64 = _T_63 | io_ins_4; // @[StickySelects.scala 47:46:@10428.4]
  assign _T_65 = _T_64 | io_ins_5; // @[StickySelects.scala 47:46:@10429.4]
  assign _T_66 = _T_65 | io_ins_6; // @[StickySelects.scala 47:46:@10430.4]
  assign _T_67 = _T_66 | io_ins_7; // @[StickySelects.scala 47:46:@10431.4]
  assign _T_68 = _T_67 | io_ins_8; // @[StickySelects.scala 47:46:@10432.4]
  assign _T_69 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@10433.4]
  assign _T_70 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 49:21:@10434.4]
  assign _T_72 = _T_62 | io_ins_2; // @[StickySelects.scala 47:46:@10437.4]
  assign _T_73 = _T_72 | io_ins_4; // @[StickySelects.scala 47:46:@10438.4]
  assign _T_74 = _T_73 | io_ins_5; // @[StickySelects.scala 47:46:@10439.4]
  assign _T_75 = _T_74 | io_ins_6; // @[StickySelects.scala 47:46:@10440.4]
  assign _T_76 = _T_75 | io_ins_7; // @[StickySelects.scala 47:46:@10441.4]
  assign _T_77 = _T_76 | io_ins_8; // @[StickySelects.scala 47:46:@10442.4]
  assign _T_78 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@10443.4]
  assign _T_79 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 49:21:@10444.4]
  assign _T_82 = _T_72 | io_ins_3; // @[StickySelects.scala 47:46:@10448.4]
  assign _T_83 = _T_82 | io_ins_5; // @[StickySelects.scala 47:46:@10449.4]
  assign _T_84 = _T_83 | io_ins_6; // @[StickySelects.scala 47:46:@10450.4]
  assign _T_85 = _T_84 | io_ins_7; // @[StickySelects.scala 47:46:@10451.4]
  assign _T_86 = _T_85 | io_ins_8; // @[StickySelects.scala 47:46:@10452.4]
  assign _T_87 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@10453.4]
  assign _T_88 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 49:21:@10454.4]
  assign _T_92 = _T_82 | io_ins_4; // @[StickySelects.scala 47:46:@10459.4]
  assign _T_93 = _T_92 | io_ins_6; // @[StickySelects.scala 47:46:@10460.4]
  assign _T_94 = _T_93 | io_ins_7; // @[StickySelects.scala 47:46:@10461.4]
  assign _T_95 = _T_94 | io_ins_8; // @[StickySelects.scala 47:46:@10462.4]
  assign _T_96 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@10463.4]
  assign _T_97 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 49:21:@10464.4]
  assign _T_102 = _T_92 | io_ins_5; // @[StickySelects.scala 47:46:@10470.4]
  assign _T_103 = _T_102 | io_ins_7; // @[StickySelects.scala 47:46:@10471.4]
  assign _T_104 = _T_103 | io_ins_8; // @[StickySelects.scala 47:46:@10472.4]
  assign _T_105 = io_ins_6 | _T_37; // @[StickySelects.scala 49:53:@10473.4]
  assign _T_106 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 49:21:@10474.4]
  assign _T_112 = _T_102 | io_ins_6; // @[StickySelects.scala 47:46:@10481.4]
  assign _T_113 = _T_112 | io_ins_8; // @[StickySelects.scala 47:46:@10482.4]
  assign _T_114 = io_ins_7 | _T_40; // @[StickySelects.scala 49:53:@10483.4]
  assign _T_115 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 49:21:@10484.4]
  assign _T_122 = _T_112 | io_ins_7; // @[StickySelects.scala 47:46:@10492.4]
  assign _T_123 = io_ins_8 | _T_43; // @[StickySelects.scala 49:53:@10493.4]
  assign _T_124 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 49:21:@10494.4]
  assign io_outs_0 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 53:57:@10496.4]
  assign io_outs_1 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 53:57:@10497.4]
  assign io_outs_2 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 53:57:@10498.4]
  assign io_outs_3 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 53:57:@10499.4]
  assign io_outs_4 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 53:57:@10500.4]
  assign io_outs_5 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 53:57:@10501.4]
  assign io_outs_6 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 53:57:@10502.4]
  assign io_outs_7 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 53:57:@10503.4]
  assign io_outs_8 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 53:57:@10504.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_37 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_40 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_43 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_51;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_59) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_60;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_69;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_77) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_78;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_86) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_87;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_95) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_96;
      end
    end
    if (reset) begin
      _T_37 <= 1'h0;
    end else begin
      if (_T_104) begin
        _T_37 <= io_ins_6;
      end else begin
        _T_37 <= _T_105;
      end
    end
    if (reset) begin
      _T_40 <= 1'h0;
    end else begin
      if (_T_113) begin
        _T_40 <= io_ins_7;
      end else begin
        _T_40 <= _T_114;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_122) begin
        _T_43 <= io_ins_8;
      end else begin
        _T_43 <= _T_123;
      end
    end
  end
endmodule
module x334_lb_0( // @[:@20040.2]
  input         clock, // @[:@20041.4]
  input         reset, // @[:@20042.4]
  input  [2:0]  io_rPort_17_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_17_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_17_ofs_0, // @[:@20043.4]
  input         io_rPort_17_en_0, // @[:@20043.4]
  input         io_rPort_17_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_17_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_16_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_16_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_16_ofs_0, // @[:@20043.4]
  input         io_rPort_16_en_0, // @[:@20043.4]
  input         io_rPort_16_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_16_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_15_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_15_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_15_ofs_0, // @[:@20043.4]
  input         io_rPort_15_en_0, // @[:@20043.4]
  input         io_rPort_15_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_15_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_14_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_14_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_14_ofs_0, // @[:@20043.4]
  input         io_rPort_14_en_0, // @[:@20043.4]
  input         io_rPort_14_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_14_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_13_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_13_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_13_ofs_0, // @[:@20043.4]
  input         io_rPort_13_en_0, // @[:@20043.4]
  input         io_rPort_13_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_13_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_12_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_12_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_12_ofs_0, // @[:@20043.4]
  input         io_rPort_12_en_0, // @[:@20043.4]
  input         io_rPort_12_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_12_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_11_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_11_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_11_ofs_0, // @[:@20043.4]
  input         io_rPort_11_en_0, // @[:@20043.4]
  input         io_rPort_11_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_11_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_10_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_10_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_10_ofs_0, // @[:@20043.4]
  input         io_rPort_10_en_0, // @[:@20043.4]
  input         io_rPort_10_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_10_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_9_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_9_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_9_ofs_0, // @[:@20043.4]
  input         io_rPort_9_en_0, // @[:@20043.4]
  input         io_rPort_9_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_9_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_8_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_8_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_8_ofs_0, // @[:@20043.4]
  input         io_rPort_8_en_0, // @[:@20043.4]
  input         io_rPort_8_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_8_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_7_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_7_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_7_ofs_0, // @[:@20043.4]
  input         io_rPort_7_en_0, // @[:@20043.4]
  input         io_rPort_7_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_7_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_6_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_6_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_6_ofs_0, // @[:@20043.4]
  input         io_rPort_6_en_0, // @[:@20043.4]
  input         io_rPort_6_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_6_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_5_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_5_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_5_ofs_0, // @[:@20043.4]
  input         io_rPort_5_en_0, // @[:@20043.4]
  input         io_rPort_5_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_5_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_4_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_4_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_4_ofs_0, // @[:@20043.4]
  input         io_rPort_4_en_0, // @[:@20043.4]
  input         io_rPort_4_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_4_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_3_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_3_ofs_0, // @[:@20043.4]
  input         io_rPort_3_en_0, // @[:@20043.4]
  input         io_rPort_3_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_3_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_2_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_2_ofs_0, // @[:@20043.4]
  input         io_rPort_2_en_0, // @[:@20043.4]
  input         io_rPort_2_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_2_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_1_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_1_ofs_0, // @[:@20043.4]
  input         io_rPort_1_en_0, // @[:@20043.4]
  input         io_rPort_1_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_1_output_0, // @[:@20043.4]
  input  [2:0]  io_rPort_0_banks_1, // @[:@20043.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@20043.4]
  input  [8:0]  io_rPort_0_ofs_0, // @[:@20043.4]
  input         io_rPort_0_en_0, // @[:@20043.4]
  input         io_rPort_0_backpressure, // @[:@20043.4]
  output [31:0] io_rPort_0_output_0, // @[:@20043.4]
  input  [2:0]  io_wPort_3_banks_1, // @[:@20043.4]
  input  [2:0]  io_wPort_3_banks_0, // @[:@20043.4]
  input  [8:0]  io_wPort_3_ofs_0, // @[:@20043.4]
  input  [31:0] io_wPort_3_data_0, // @[:@20043.4]
  input         io_wPort_3_en_0, // @[:@20043.4]
  input  [2:0]  io_wPort_2_banks_1, // @[:@20043.4]
  input  [2:0]  io_wPort_2_banks_0, // @[:@20043.4]
  input  [8:0]  io_wPort_2_ofs_0, // @[:@20043.4]
  input  [31:0] io_wPort_2_data_0, // @[:@20043.4]
  input         io_wPort_2_en_0, // @[:@20043.4]
  input  [2:0]  io_wPort_1_banks_1, // @[:@20043.4]
  input  [2:0]  io_wPort_1_banks_0, // @[:@20043.4]
  input  [8:0]  io_wPort_1_ofs_0, // @[:@20043.4]
  input  [31:0] io_wPort_1_data_0, // @[:@20043.4]
  input         io_wPort_1_en_0, // @[:@20043.4]
  input  [2:0]  io_wPort_0_banks_1, // @[:@20043.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@20043.4]
  input  [8:0]  io_wPort_0_ofs_0, // @[:@20043.4]
  input  [31:0] io_wPort_0_data_0, // @[:@20043.4]
  input         io_wPort_0_en_0 // @[:@20043.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@20186.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@20186.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20186.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20186.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20186.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@20186.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@20186.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@20186.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@20202.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@20202.4]
  wire [8:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20202.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20202.4]
  wire [8:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20202.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@20202.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@20202.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@20202.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@20218.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@20218.4]
  wire [8:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20218.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20218.4]
  wire [8:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20218.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@20218.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@20218.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@20218.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@20234.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@20234.4]
  wire [8:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20234.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20234.4]
  wire [8:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20234.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@20234.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@20234.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@20234.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@20250.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@20250.4]
  wire [8:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20250.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20250.4]
  wire [8:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20250.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@20250.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@20250.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@20250.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@20266.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@20266.4]
  wire [8:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20266.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20266.4]
  wire [8:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20266.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@20266.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@20266.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@20266.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@20282.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@20282.4]
  wire [8:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20282.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20282.4]
  wire [8:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20282.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@20282.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@20282.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@20282.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@20298.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@20298.4]
  wire [8:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20298.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20298.4]
  wire [8:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20298.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@20298.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@20298.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@20298.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@20314.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@20314.4]
  wire [8:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20314.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20314.4]
  wire [8:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20314.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@20314.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@20314.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@20314.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@20330.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@20330.4]
  wire [8:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20330.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20330.4]
  wire [8:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20330.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@20330.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@20330.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@20330.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@20346.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@20346.4]
  wire [8:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20346.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20346.4]
  wire [8:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20346.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@20346.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@20346.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@20346.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@20362.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@20362.4]
  wire [8:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20362.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20362.4]
  wire [8:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20362.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@20362.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@20362.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@20362.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@20378.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@20378.4]
  wire [8:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20378.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20378.4]
  wire [8:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20378.4]
  wire [31:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@20378.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@20378.4]
  wire [31:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@20378.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@20394.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@20394.4]
  wire [8:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20394.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20394.4]
  wire [8:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20394.4]
  wire [31:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@20394.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@20394.4]
  wire [31:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@20394.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@20410.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@20410.4]
  wire [8:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20410.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20410.4]
  wire [8:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20410.4]
  wire [31:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@20410.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@20410.4]
  wire [31:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@20410.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@20426.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@20426.4]
  wire [8:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20426.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20426.4]
  wire [8:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20426.4]
  wire [31:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@20426.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@20426.4]
  wire [31:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@20426.4]
  wire  Mem1D_16_clock; // @[MemPrimitives.scala 64:21:@20442.4]
  wire  Mem1D_16_reset; // @[MemPrimitives.scala 64:21:@20442.4]
  wire [8:0] Mem1D_16_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20442.4]
  wire  Mem1D_16_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20442.4]
  wire [8:0] Mem1D_16_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20442.4]
  wire [31:0] Mem1D_16_io_w_data_0; // @[MemPrimitives.scala 64:21:@20442.4]
  wire  Mem1D_16_io_w_en_0; // @[MemPrimitives.scala 64:21:@20442.4]
  wire [31:0] Mem1D_16_io_output; // @[MemPrimitives.scala 64:21:@20442.4]
  wire  Mem1D_17_clock; // @[MemPrimitives.scala 64:21:@20458.4]
  wire  Mem1D_17_reset; // @[MemPrimitives.scala 64:21:@20458.4]
  wire [8:0] Mem1D_17_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20458.4]
  wire  Mem1D_17_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20458.4]
  wire [8:0] Mem1D_17_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20458.4]
  wire [31:0] Mem1D_17_io_w_data_0; // @[MemPrimitives.scala 64:21:@20458.4]
  wire  Mem1D_17_io_w_en_0; // @[MemPrimitives.scala 64:21:@20458.4]
  wire [31:0] Mem1D_17_io_output; // @[MemPrimitives.scala 64:21:@20458.4]
  wire  Mem1D_18_clock; // @[MemPrimitives.scala 64:21:@20474.4]
  wire  Mem1D_18_reset; // @[MemPrimitives.scala 64:21:@20474.4]
  wire [8:0] Mem1D_18_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20474.4]
  wire  Mem1D_18_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20474.4]
  wire [8:0] Mem1D_18_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20474.4]
  wire [31:0] Mem1D_18_io_w_data_0; // @[MemPrimitives.scala 64:21:@20474.4]
  wire  Mem1D_18_io_w_en_0; // @[MemPrimitives.scala 64:21:@20474.4]
  wire [31:0] Mem1D_18_io_output; // @[MemPrimitives.scala 64:21:@20474.4]
  wire  Mem1D_19_clock; // @[MemPrimitives.scala 64:21:@20490.4]
  wire  Mem1D_19_reset; // @[MemPrimitives.scala 64:21:@20490.4]
  wire [8:0] Mem1D_19_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20490.4]
  wire  Mem1D_19_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20490.4]
  wire [8:0] Mem1D_19_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20490.4]
  wire [31:0] Mem1D_19_io_w_data_0; // @[MemPrimitives.scala 64:21:@20490.4]
  wire  Mem1D_19_io_w_en_0; // @[MemPrimitives.scala 64:21:@20490.4]
  wire [31:0] Mem1D_19_io_output; // @[MemPrimitives.scala 64:21:@20490.4]
  wire  Mem1D_20_clock; // @[MemPrimitives.scala 64:21:@20506.4]
  wire  Mem1D_20_reset; // @[MemPrimitives.scala 64:21:@20506.4]
  wire [8:0] Mem1D_20_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20506.4]
  wire  Mem1D_20_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20506.4]
  wire [8:0] Mem1D_20_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20506.4]
  wire [31:0] Mem1D_20_io_w_data_0; // @[MemPrimitives.scala 64:21:@20506.4]
  wire  Mem1D_20_io_w_en_0; // @[MemPrimitives.scala 64:21:@20506.4]
  wire [31:0] Mem1D_20_io_output; // @[MemPrimitives.scala 64:21:@20506.4]
  wire  Mem1D_21_clock; // @[MemPrimitives.scala 64:21:@20522.4]
  wire  Mem1D_21_reset; // @[MemPrimitives.scala 64:21:@20522.4]
  wire [8:0] Mem1D_21_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20522.4]
  wire  Mem1D_21_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20522.4]
  wire [8:0] Mem1D_21_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20522.4]
  wire [31:0] Mem1D_21_io_w_data_0; // @[MemPrimitives.scala 64:21:@20522.4]
  wire  Mem1D_21_io_w_en_0; // @[MemPrimitives.scala 64:21:@20522.4]
  wire [31:0] Mem1D_21_io_output; // @[MemPrimitives.scala 64:21:@20522.4]
  wire  Mem1D_22_clock; // @[MemPrimitives.scala 64:21:@20538.4]
  wire  Mem1D_22_reset; // @[MemPrimitives.scala 64:21:@20538.4]
  wire [8:0] Mem1D_22_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20538.4]
  wire  Mem1D_22_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20538.4]
  wire [8:0] Mem1D_22_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20538.4]
  wire [31:0] Mem1D_22_io_w_data_0; // @[MemPrimitives.scala 64:21:@20538.4]
  wire  Mem1D_22_io_w_en_0; // @[MemPrimitives.scala 64:21:@20538.4]
  wire [31:0] Mem1D_22_io_output; // @[MemPrimitives.scala 64:21:@20538.4]
  wire  Mem1D_23_clock; // @[MemPrimitives.scala 64:21:@20554.4]
  wire  Mem1D_23_reset; // @[MemPrimitives.scala 64:21:@20554.4]
  wire [8:0] Mem1D_23_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@20554.4]
  wire  Mem1D_23_io_r_backpressure; // @[MemPrimitives.scala 64:21:@20554.4]
  wire [8:0] Mem1D_23_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@20554.4]
  wire [31:0] Mem1D_23_io_w_data_0; // @[MemPrimitives.scala 64:21:@20554.4]
  wire  Mem1D_23_io_w_en_0; // @[MemPrimitives.scala 64:21:@20554.4]
  wire [31:0] Mem1D_23_io_output; // @[MemPrimitives.scala 64:21:@20554.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_6; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_7; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_ins_8; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_6; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_7; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_io_outs_8; // @[MemPrimitives.scala 124:33:@21062.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_6; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_7; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_ins_8; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_6; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_7; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_1_io_outs_8; // @[MemPrimitives.scala 124:33:@21151.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_ins_8; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_2_io_outs_8; // @[MemPrimitives.scala 124:33:@21240.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_ins_8; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_3_io_outs_8; // @[MemPrimitives.scala 124:33:@21329.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_6; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_7; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_ins_8; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_6; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_7; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_4_io_outs_8; // @[MemPrimitives.scala 124:33:@21418.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_6; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_7; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_ins_8; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_6; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_7; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_5_io_outs_8; // @[MemPrimitives.scala 124:33:@21507.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_ins_8; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_6_io_outs_8; // @[MemPrimitives.scala 124:33:@21596.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_ins_8; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_7_io_outs_8; // @[MemPrimitives.scala 124:33:@21685.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_6; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_7; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_ins_8; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_6; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_7; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_8_io_outs_8; // @[MemPrimitives.scala 124:33:@21774.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_6; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_7; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_ins_8; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_6; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_7; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_9_io_outs_8; // @[MemPrimitives.scala 124:33:@21863.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_ins_8; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_10_io_outs_8; // @[MemPrimitives.scala 124:33:@21952.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_ins_8; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_11_io_outs_8; // @[MemPrimitives.scala 124:33:@22041.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_6; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_7; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_ins_8; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_6; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_7; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_12_io_outs_8; // @[MemPrimitives.scala 124:33:@22130.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_6; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_7; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_ins_8; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_6; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_7; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_13_io_outs_8; // @[MemPrimitives.scala 124:33:@22219.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_6; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_7; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_ins_8; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_6; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_7; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_14_io_outs_8; // @[MemPrimitives.scala 124:33:@22308.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_6; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_7; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_ins_8; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_6; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_7; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_15_io_outs_8; // @[MemPrimitives.scala 124:33:@22397.4]
  wire  StickySelects_16_clock; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_reset; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_0; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_1; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_2; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_3; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_4; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_5; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_6; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_7; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_ins_8; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_0; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_1; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_2; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_3; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_4; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_5; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_6; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_7; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_16_io_outs_8; // @[MemPrimitives.scala 124:33:@22486.4]
  wire  StickySelects_17_clock; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_reset; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_0; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_1; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_2; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_3; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_4; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_5; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_6; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_7; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_ins_8; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_0; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_1; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_2; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_3; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_4; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_5; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_6; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_7; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_17_io_outs_8; // @[MemPrimitives.scala 124:33:@22575.4]
  wire  StickySelects_18_clock; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_reset; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_0; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_1; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_2; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_3; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_4; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_5; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_6; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_7; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_ins_8; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_0; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_1; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_2; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_3; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_4; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_5; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_6; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_7; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_18_io_outs_8; // @[MemPrimitives.scala 124:33:@22664.4]
  wire  StickySelects_19_clock; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_reset; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_0; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_1; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_2; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_3; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_4; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_5; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_6; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_7; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_ins_8; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_0; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_1; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_2; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_3; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_4; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_5; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_6; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_7; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_19_io_outs_8; // @[MemPrimitives.scala 124:33:@22753.4]
  wire  StickySelects_20_clock; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_reset; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_0; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_1; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_2; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_3; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_4; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_5; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_6; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_7; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_ins_8; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_0; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_1; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_2; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_3; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_4; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_5; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_6; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_7; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_20_io_outs_8; // @[MemPrimitives.scala 124:33:@22842.4]
  wire  StickySelects_21_clock; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_reset; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_0; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_1; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_2; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_3; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_4; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_5; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_6; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_7; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_ins_8; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_0; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_1; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_2; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_3; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_4; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_5; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_6; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_7; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_21_io_outs_8; // @[MemPrimitives.scala 124:33:@22931.4]
  wire  StickySelects_22_clock; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_reset; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_0; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_1; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_2; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_3; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_4; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_5; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_6; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_7; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_ins_8; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_0; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_1; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_2; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_3; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_4; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_5; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_6; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_7; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_22_io_outs_8; // @[MemPrimitives.scala 124:33:@23020.4]
  wire  StickySelects_23_clock; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_reset; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_0; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_1; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_2; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_3; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_4; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_5; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_6; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_7; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_ins_8; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_0; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_1; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_2; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_3; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_4; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_5; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_6; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_7; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  StickySelects_23_io_outs_8; // @[MemPrimitives.scala 124:33:@23109.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@23199.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@23199.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@23199.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@23199.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@23199.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@23207.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@23207.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@23207.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@23207.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@23207.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@23215.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@23215.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@23215.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@23215.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@23215.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@23223.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@23223.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@23223.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@23223.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@23223.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@23231.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@23231.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@23231.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@23231.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@23231.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@23239.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@23239.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@23239.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@23239.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@23239.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@23247.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@23247.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@23247.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@23247.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@23247.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@23255.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@23255.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@23255.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@23255.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@23255.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@23263.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@23263.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@23263.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@23263.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@23263.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@23271.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@23271.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@23271.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@23271.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@23271.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@23279.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@23279.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@23279.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@23279.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@23279.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@23287.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@23287.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@23287.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@23287.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@23287.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@23343.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@23343.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@23343.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@23343.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@23343.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@23351.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@23351.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@23351.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@23351.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@23351.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@23359.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@23359.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@23359.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@23359.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@23359.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@23367.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@23367.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@23367.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@23367.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@23367.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@23375.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@23375.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@23375.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@23375.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@23375.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@23383.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@23383.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@23383.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@23383.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@23383.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@23391.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@23391.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@23391.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@23391.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@23391.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@23399.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@23399.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@23399.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@23399.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@23399.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@23407.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@23407.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@23407.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@23407.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@23407.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@23415.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@23415.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@23415.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@23415.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@23415.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@23423.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@23423.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@23423.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@23423.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@23423.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@23431.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@23431.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@23431.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@23431.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@23431.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@23487.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@23487.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@23487.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@23487.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@23487.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@23495.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@23495.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@23495.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@23495.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@23495.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@23503.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@23503.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@23503.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@23503.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@23503.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@23511.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@23511.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@23511.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@23511.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@23511.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@23519.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@23519.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@23519.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@23519.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@23519.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@23527.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@23527.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@23527.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@23527.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@23527.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@23535.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@23535.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@23535.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@23535.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@23535.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@23543.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@23543.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@23543.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@23543.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@23543.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@23551.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@23551.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@23551.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@23551.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@23551.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@23559.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@23559.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@23559.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@23559.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@23559.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@23567.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@23567.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@23567.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@23567.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@23567.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@23575.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@23575.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@23575.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@23575.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@23575.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@23631.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@23631.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@23631.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@23631.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@23631.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@23639.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@23639.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@23639.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@23639.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@23639.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@23647.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@23647.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@23647.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@23647.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@23647.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@23655.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@23655.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@23655.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@23655.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@23655.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@23663.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@23663.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@23663.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@23663.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@23663.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@23671.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@23671.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@23671.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@23671.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@23671.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@23679.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@23679.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@23679.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@23679.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@23679.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@23687.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@23687.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@23687.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@23687.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@23687.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@23695.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@23695.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@23695.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@23695.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@23695.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@23703.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@23703.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@23703.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@23703.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@23703.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@23711.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@23711.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@23711.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@23711.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@23711.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@23719.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@23719.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@23719.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@23719.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@23719.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@23775.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@23775.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@23775.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@23775.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@23775.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@23783.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@23783.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@23783.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@23783.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@23783.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@23791.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@23791.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@23791.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@23791.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@23791.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@23799.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@23799.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@23799.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@23799.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@23799.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@23807.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@23807.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@23807.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@23807.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@23807.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@23815.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@23815.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@23815.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@23815.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@23815.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@23823.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@23823.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@23823.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@23823.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@23823.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@23831.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@23831.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@23831.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@23831.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@23831.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@23839.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@23839.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@23839.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@23839.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@23839.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@23847.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@23847.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@23847.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@23847.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@23847.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@23855.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@23855.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@23855.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@23855.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@23855.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@23863.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@23863.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@23863.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@23863.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@23863.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@23919.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@23919.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@23919.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@23919.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@23919.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@23927.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@23927.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@23927.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@23927.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@23927.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@23935.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@23935.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@23935.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@23935.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@23935.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@23943.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@23943.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@23943.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@23943.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@23943.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@23951.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@23951.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@23951.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@23951.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@23951.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@23959.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@23959.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@23959.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@23959.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@23959.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@23967.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@23967.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@23967.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@23967.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@23967.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@23975.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@23975.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@23975.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@23975.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@23975.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@23983.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@23983.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@23983.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@23983.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@23983.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@23991.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@23991.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@23991.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@23991.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@23991.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@23999.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@23999.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@23999.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@23999.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@23999.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@24007.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@24007.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@24007.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@24007.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@24007.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@24063.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@24063.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@24063.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@24063.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@24063.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@24071.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@24071.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@24071.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@24071.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@24071.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@24079.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@24079.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@24079.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@24079.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@24079.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@24087.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@24087.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@24087.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@24087.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@24087.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@24095.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@24095.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@24095.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@24095.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@24095.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@24103.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@24103.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@24103.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@24103.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@24103.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@24111.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@24111.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@24111.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@24111.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@24111.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@24119.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@24119.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@24119.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@24119.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@24119.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@24127.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@24127.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@24127.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@24127.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@24127.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@24135.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@24135.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@24135.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@24135.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@24135.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@24143.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@24143.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@24143.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@24143.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@24143.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@24151.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@24151.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@24151.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@24151.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@24151.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@24207.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@24207.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@24207.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@24207.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@24207.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@24215.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@24215.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@24215.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@24215.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@24215.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@24223.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@24223.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@24223.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@24223.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@24223.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@24231.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@24231.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@24231.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@24231.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@24231.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@24239.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@24239.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@24239.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@24239.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@24239.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@24247.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@24247.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@24247.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@24247.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@24247.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@24255.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@24255.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@24255.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@24255.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@24255.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@24263.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@24263.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@24263.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@24263.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@24263.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@24271.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@24271.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@24271.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@24271.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@24271.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@24279.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@24279.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@24279.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@24279.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@24279.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@24287.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@24287.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@24287.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@24287.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@24287.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@24295.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@24295.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@24295.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@24295.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@24295.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@24351.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@24351.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@24351.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@24351.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@24351.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@24359.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@24359.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@24359.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@24359.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@24359.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@24367.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@24367.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@24367.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@24367.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@24367.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@24375.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@24375.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@24375.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@24375.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@24375.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@24383.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@24383.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@24383.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@24383.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@24383.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@24391.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@24391.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@24391.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@24391.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@24391.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@24399.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@24399.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@24399.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@24399.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@24399.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@24407.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@24407.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@24407.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@24407.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@24407.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@24415.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@24415.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@24415.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@24415.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@24415.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@24423.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@24423.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@24423.4]
  wire  RetimeWrapper_105_io_in; // @[package.scala 93:22:@24423.4]
  wire  RetimeWrapper_105_io_out; // @[package.scala 93:22:@24423.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@24431.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@24431.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@24431.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@24431.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@24431.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@24439.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@24439.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@24439.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@24439.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@24439.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@24495.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@24495.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@24495.4]
  wire  RetimeWrapper_108_io_in; // @[package.scala 93:22:@24495.4]
  wire  RetimeWrapper_108_io_out; // @[package.scala 93:22:@24495.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@24503.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@24503.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@24503.4]
  wire  RetimeWrapper_109_io_in; // @[package.scala 93:22:@24503.4]
  wire  RetimeWrapper_109_io_out; // @[package.scala 93:22:@24503.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@24511.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@24511.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@24511.4]
  wire  RetimeWrapper_110_io_in; // @[package.scala 93:22:@24511.4]
  wire  RetimeWrapper_110_io_out; // @[package.scala 93:22:@24511.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@24519.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@24519.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@24519.4]
  wire  RetimeWrapper_111_io_in; // @[package.scala 93:22:@24519.4]
  wire  RetimeWrapper_111_io_out; // @[package.scala 93:22:@24519.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@24527.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@24527.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@24527.4]
  wire  RetimeWrapper_112_io_in; // @[package.scala 93:22:@24527.4]
  wire  RetimeWrapper_112_io_out; // @[package.scala 93:22:@24527.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@24535.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@24535.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@24535.4]
  wire  RetimeWrapper_113_io_in; // @[package.scala 93:22:@24535.4]
  wire  RetimeWrapper_113_io_out; // @[package.scala 93:22:@24535.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@24543.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@24543.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@24543.4]
  wire  RetimeWrapper_114_io_in; // @[package.scala 93:22:@24543.4]
  wire  RetimeWrapper_114_io_out; // @[package.scala 93:22:@24543.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@24551.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@24551.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@24551.4]
  wire  RetimeWrapper_115_io_in; // @[package.scala 93:22:@24551.4]
  wire  RetimeWrapper_115_io_out; // @[package.scala 93:22:@24551.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@24559.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@24559.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@24559.4]
  wire  RetimeWrapper_116_io_in; // @[package.scala 93:22:@24559.4]
  wire  RetimeWrapper_116_io_out; // @[package.scala 93:22:@24559.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@24567.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@24567.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@24567.4]
  wire  RetimeWrapper_117_io_in; // @[package.scala 93:22:@24567.4]
  wire  RetimeWrapper_117_io_out; // @[package.scala 93:22:@24567.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@24575.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@24575.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@24575.4]
  wire  RetimeWrapper_118_io_in; // @[package.scala 93:22:@24575.4]
  wire  RetimeWrapper_118_io_out; // @[package.scala 93:22:@24575.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@24583.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@24583.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@24583.4]
  wire  RetimeWrapper_119_io_in; // @[package.scala 93:22:@24583.4]
  wire  RetimeWrapper_119_io_out; // @[package.scala 93:22:@24583.4]
  wire  RetimeWrapper_120_clock; // @[package.scala 93:22:@24639.4]
  wire  RetimeWrapper_120_reset; // @[package.scala 93:22:@24639.4]
  wire  RetimeWrapper_120_io_flow; // @[package.scala 93:22:@24639.4]
  wire  RetimeWrapper_120_io_in; // @[package.scala 93:22:@24639.4]
  wire  RetimeWrapper_120_io_out; // @[package.scala 93:22:@24639.4]
  wire  RetimeWrapper_121_clock; // @[package.scala 93:22:@24647.4]
  wire  RetimeWrapper_121_reset; // @[package.scala 93:22:@24647.4]
  wire  RetimeWrapper_121_io_flow; // @[package.scala 93:22:@24647.4]
  wire  RetimeWrapper_121_io_in; // @[package.scala 93:22:@24647.4]
  wire  RetimeWrapper_121_io_out; // @[package.scala 93:22:@24647.4]
  wire  RetimeWrapper_122_clock; // @[package.scala 93:22:@24655.4]
  wire  RetimeWrapper_122_reset; // @[package.scala 93:22:@24655.4]
  wire  RetimeWrapper_122_io_flow; // @[package.scala 93:22:@24655.4]
  wire  RetimeWrapper_122_io_in; // @[package.scala 93:22:@24655.4]
  wire  RetimeWrapper_122_io_out; // @[package.scala 93:22:@24655.4]
  wire  RetimeWrapper_123_clock; // @[package.scala 93:22:@24663.4]
  wire  RetimeWrapper_123_reset; // @[package.scala 93:22:@24663.4]
  wire  RetimeWrapper_123_io_flow; // @[package.scala 93:22:@24663.4]
  wire  RetimeWrapper_123_io_in; // @[package.scala 93:22:@24663.4]
  wire  RetimeWrapper_123_io_out; // @[package.scala 93:22:@24663.4]
  wire  RetimeWrapper_124_clock; // @[package.scala 93:22:@24671.4]
  wire  RetimeWrapper_124_reset; // @[package.scala 93:22:@24671.4]
  wire  RetimeWrapper_124_io_flow; // @[package.scala 93:22:@24671.4]
  wire  RetimeWrapper_124_io_in; // @[package.scala 93:22:@24671.4]
  wire  RetimeWrapper_124_io_out; // @[package.scala 93:22:@24671.4]
  wire  RetimeWrapper_125_clock; // @[package.scala 93:22:@24679.4]
  wire  RetimeWrapper_125_reset; // @[package.scala 93:22:@24679.4]
  wire  RetimeWrapper_125_io_flow; // @[package.scala 93:22:@24679.4]
  wire  RetimeWrapper_125_io_in; // @[package.scala 93:22:@24679.4]
  wire  RetimeWrapper_125_io_out; // @[package.scala 93:22:@24679.4]
  wire  RetimeWrapper_126_clock; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_126_reset; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_126_io_flow; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_126_io_in; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_126_io_out; // @[package.scala 93:22:@24687.4]
  wire  RetimeWrapper_127_clock; // @[package.scala 93:22:@24695.4]
  wire  RetimeWrapper_127_reset; // @[package.scala 93:22:@24695.4]
  wire  RetimeWrapper_127_io_flow; // @[package.scala 93:22:@24695.4]
  wire  RetimeWrapper_127_io_in; // @[package.scala 93:22:@24695.4]
  wire  RetimeWrapper_127_io_out; // @[package.scala 93:22:@24695.4]
  wire  RetimeWrapper_128_clock; // @[package.scala 93:22:@24703.4]
  wire  RetimeWrapper_128_reset; // @[package.scala 93:22:@24703.4]
  wire  RetimeWrapper_128_io_flow; // @[package.scala 93:22:@24703.4]
  wire  RetimeWrapper_128_io_in; // @[package.scala 93:22:@24703.4]
  wire  RetimeWrapper_128_io_out; // @[package.scala 93:22:@24703.4]
  wire  RetimeWrapper_129_clock; // @[package.scala 93:22:@24711.4]
  wire  RetimeWrapper_129_reset; // @[package.scala 93:22:@24711.4]
  wire  RetimeWrapper_129_io_flow; // @[package.scala 93:22:@24711.4]
  wire  RetimeWrapper_129_io_in; // @[package.scala 93:22:@24711.4]
  wire  RetimeWrapper_129_io_out; // @[package.scala 93:22:@24711.4]
  wire  RetimeWrapper_130_clock; // @[package.scala 93:22:@24719.4]
  wire  RetimeWrapper_130_reset; // @[package.scala 93:22:@24719.4]
  wire  RetimeWrapper_130_io_flow; // @[package.scala 93:22:@24719.4]
  wire  RetimeWrapper_130_io_in; // @[package.scala 93:22:@24719.4]
  wire  RetimeWrapper_130_io_out; // @[package.scala 93:22:@24719.4]
  wire  RetimeWrapper_131_clock; // @[package.scala 93:22:@24727.4]
  wire  RetimeWrapper_131_reset; // @[package.scala 93:22:@24727.4]
  wire  RetimeWrapper_131_io_flow; // @[package.scala 93:22:@24727.4]
  wire  RetimeWrapper_131_io_in; // @[package.scala 93:22:@24727.4]
  wire  RetimeWrapper_131_io_out; // @[package.scala 93:22:@24727.4]
  wire  RetimeWrapper_132_clock; // @[package.scala 93:22:@24783.4]
  wire  RetimeWrapper_132_reset; // @[package.scala 93:22:@24783.4]
  wire  RetimeWrapper_132_io_flow; // @[package.scala 93:22:@24783.4]
  wire  RetimeWrapper_132_io_in; // @[package.scala 93:22:@24783.4]
  wire  RetimeWrapper_132_io_out; // @[package.scala 93:22:@24783.4]
  wire  RetimeWrapper_133_clock; // @[package.scala 93:22:@24791.4]
  wire  RetimeWrapper_133_reset; // @[package.scala 93:22:@24791.4]
  wire  RetimeWrapper_133_io_flow; // @[package.scala 93:22:@24791.4]
  wire  RetimeWrapper_133_io_in; // @[package.scala 93:22:@24791.4]
  wire  RetimeWrapper_133_io_out; // @[package.scala 93:22:@24791.4]
  wire  RetimeWrapper_134_clock; // @[package.scala 93:22:@24799.4]
  wire  RetimeWrapper_134_reset; // @[package.scala 93:22:@24799.4]
  wire  RetimeWrapper_134_io_flow; // @[package.scala 93:22:@24799.4]
  wire  RetimeWrapper_134_io_in; // @[package.scala 93:22:@24799.4]
  wire  RetimeWrapper_134_io_out; // @[package.scala 93:22:@24799.4]
  wire  RetimeWrapper_135_clock; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_135_reset; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_135_io_flow; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_135_io_in; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_135_io_out; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_136_clock; // @[package.scala 93:22:@24815.4]
  wire  RetimeWrapper_136_reset; // @[package.scala 93:22:@24815.4]
  wire  RetimeWrapper_136_io_flow; // @[package.scala 93:22:@24815.4]
  wire  RetimeWrapper_136_io_in; // @[package.scala 93:22:@24815.4]
  wire  RetimeWrapper_136_io_out; // @[package.scala 93:22:@24815.4]
  wire  RetimeWrapper_137_clock; // @[package.scala 93:22:@24823.4]
  wire  RetimeWrapper_137_reset; // @[package.scala 93:22:@24823.4]
  wire  RetimeWrapper_137_io_flow; // @[package.scala 93:22:@24823.4]
  wire  RetimeWrapper_137_io_in; // @[package.scala 93:22:@24823.4]
  wire  RetimeWrapper_137_io_out; // @[package.scala 93:22:@24823.4]
  wire  RetimeWrapper_138_clock; // @[package.scala 93:22:@24831.4]
  wire  RetimeWrapper_138_reset; // @[package.scala 93:22:@24831.4]
  wire  RetimeWrapper_138_io_flow; // @[package.scala 93:22:@24831.4]
  wire  RetimeWrapper_138_io_in; // @[package.scala 93:22:@24831.4]
  wire  RetimeWrapper_138_io_out; // @[package.scala 93:22:@24831.4]
  wire  RetimeWrapper_139_clock; // @[package.scala 93:22:@24839.4]
  wire  RetimeWrapper_139_reset; // @[package.scala 93:22:@24839.4]
  wire  RetimeWrapper_139_io_flow; // @[package.scala 93:22:@24839.4]
  wire  RetimeWrapper_139_io_in; // @[package.scala 93:22:@24839.4]
  wire  RetimeWrapper_139_io_out; // @[package.scala 93:22:@24839.4]
  wire  RetimeWrapper_140_clock; // @[package.scala 93:22:@24847.4]
  wire  RetimeWrapper_140_reset; // @[package.scala 93:22:@24847.4]
  wire  RetimeWrapper_140_io_flow; // @[package.scala 93:22:@24847.4]
  wire  RetimeWrapper_140_io_in; // @[package.scala 93:22:@24847.4]
  wire  RetimeWrapper_140_io_out; // @[package.scala 93:22:@24847.4]
  wire  RetimeWrapper_141_clock; // @[package.scala 93:22:@24855.4]
  wire  RetimeWrapper_141_reset; // @[package.scala 93:22:@24855.4]
  wire  RetimeWrapper_141_io_flow; // @[package.scala 93:22:@24855.4]
  wire  RetimeWrapper_141_io_in; // @[package.scala 93:22:@24855.4]
  wire  RetimeWrapper_141_io_out; // @[package.scala 93:22:@24855.4]
  wire  RetimeWrapper_142_clock; // @[package.scala 93:22:@24863.4]
  wire  RetimeWrapper_142_reset; // @[package.scala 93:22:@24863.4]
  wire  RetimeWrapper_142_io_flow; // @[package.scala 93:22:@24863.4]
  wire  RetimeWrapper_142_io_in; // @[package.scala 93:22:@24863.4]
  wire  RetimeWrapper_142_io_out; // @[package.scala 93:22:@24863.4]
  wire  RetimeWrapper_143_clock; // @[package.scala 93:22:@24871.4]
  wire  RetimeWrapper_143_reset; // @[package.scala 93:22:@24871.4]
  wire  RetimeWrapper_143_io_flow; // @[package.scala 93:22:@24871.4]
  wire  RetimeWrapper_143_io_in; // @[package.scala 93:22:@24871.4]
  wire  RetimeWrapper_143_io_out; // @[package.scala 93:22:@24871.4]
  wire  RetimeWrapper_144_clock; // @[package.scala 93:22:@24927.4]
  wire  RetimeWrapper_144_reset; // @[package.scala 93:22:@24927.4]
  wire  RetimeWrapper_144_io_flow; // @[package.scala 93:22:@24927.4]
  wire  RetimeWrapper_144_io_in; // @[package.scala 93:22:@24927.4]
  wire  RetimeWrapper_144_io_out; // @[package.scala 93:22:@24927.4]
  wire  RetimeWrapper_145_clock; // @[package.scala 93:22:@24935.4]
  wire  RetimeWrapper_145_reset; // @[package.scala 93:22:@24935.4]
  wire  RetimeWrapper_145_io_flow; // @[package.scala 93:22:@24935.4]
  wire  RetimeWrapper_145_io_in; // @[package.scala 93:22:@24935.4]
  wire  RetimeWrapper_145_io_out; // @[package.scala 93:22:@24935.4]
  wire  RetimeWrapper_146_clock; // @[package.scala 93:22:@24943.4]
  wire  RetimeWrapper_146_reset; // @[package.scala 93:22:@24943.4]
  wire  RetimeWrapper_146_io_flow; // @[package.scala 93:22:@24943.4]
  wire  RetimeWrapper_146_io_in; // @[package.scala 93:22:@24943.4]
  wire  RetimeWrapper_146_io_out; // @[package.scala 93:22:@24943.4]
  wire  RetimeWrapper_147_clock; // @[package.scala 93:22:@24951.4]
  wire  RetimeWrapper_147_reset; // @[package.scala 93:22:@24951.4]
  wire  RetimeWrapper_147_io_flow; // @[package.scala 93:22:@24951.4]
  wire  RetimeWrapper_147_io_in; // @[package.scala 93:22:@24951.4]
  wire  RetimeWrapper_147_io_out; // @[package.scala 93:22:@24951.4]
  wire  RetimeWrapper_148_clock; // @[package.scala 93:22:@24959.4]
  wire  RetimeWrapper_148_reset; // @[package.scala 93:22:@24959.4]
  wire  RetimeWrapper_148_io_flow; // @[package.scala 93:22:@24959.4]
  wire  RetimeWrapper_148_io_in; // @[package.scala 93:22:@24959.4]
  wire  RetimeWrapper_148_io_out; // @[package.scala 93:22:@24959.4]
  wire  RetimeWrapper_149_clock; // @[package.scala 93:22:@24967.4]
  wire  RetimeWrapper_149_reset; // @[package.scala 93:22:@24967.4]
  wire  RetimeWrapper_149_io_flow; // @[package.scala 93:22:@24967.4]
  wire  RetimeWrapper_149_io_in; // @[package.scala 93:22:@24967.4]
  wire  RetimeWrapper_149_io_out; // @[package.scala 93:22:@24967.4]
  wire  RetimeWrapper_150_clock; // @[package.scala 93:22:@24975.4]
  wire  RetimeWrapper_150_reset; // @[package.scala 93:22:@24975.4]
  wire  RetimeWrapper_150_io_flow; // @[package.scala 93:22:@24975.4]
  wire  RetimeWrapper_150_io_in; // @[package.scala 93:22:@24975.4]
  wire  RetimeWrapper_150_io_out; // @[package.scala 93:22:@24975.4]
  wire  RetimeWrapper_151_clock; // @[package.scala 93:22:@24983.4]
  wire  RetimeWrapper_151_reset; // @[package.scala 93:22:@24983.4]
  wire  RetimeWrapper_151_io_flow; // @[package.scala 93:22:@24983.4]
  wire  RetimeWrapper_151_io_in; // @[package.scala 93:22:@24983.4]
  wire  RetimeWrapper_151_io_out; // @[package.scala 93:22:@24983.4]
  wire  RetimeWrapper_152_clock; // @[package.scala 93:22:@24991.4]
  wire  RetimeWrapper_152_reset; // @[package.scala 93:22:@24991.4]
  wire  RetimeWrapper_152_io_flow; // @[package.scala 93:22:@24991.4]
  wire  RetimeWrapper_152_io_in; // @[package.scala 93:22:@24991.4]
  wire  RetimeWrapper_152_io_out; // @[package.scala 93:22:@24991.4]
  wire  RetimeWrapper_153_clock; // @[package.scala 93:22:@24999.4]
  wire  RetimeWrapper_153_reset; // @[package.scala 93:22:@24999.4]
  wire  RetimeWrapper_153_io_flow; // @[package.scala 93:22:@24999.4]
  wire  RetimeWrapper_153_io_in; // @[package.scala 93:22:@24999.4]
  wire  RetimeWrapper_153_io_out; // @[package.scala 93:22:@24999.4]
  wire  RetimeWrapper_154_clock; // @[package.scala 93:22:@25007.4]
  wire  RetimeWrapper_154_reset; // @[package.scala 93:22:@25007.4]
  wire  RetimeWrapper_154_io_flow; // @[package.scala 93:22:@25007.4]
  wire  RetimeWrapper_154_io_in; // @[package.scala 93:22:@25007.4]
  wire  RetimeWrapper_154_io_out; // @[package.scala 93:22:@25007.4]
  wire  RetimeWrapper_155_clock; // @[package.scala 93:22:@25015.4]
  wire  RetimeWrapper_155_reset; // @[package.scala 93:22:@25015.4]
  wire  RetimeWrapper_155_io_flow; // @[package.scala 93:22:@25015.4]
  wire  RetimeWrapper_155_io_in; // @[package.scala 93:22:@25015.4]
  wire  RetimeWrapper_155_io_out; // @[package.scala 93:22:@25015.4]
  wire  RetimeWrapper_156_clock; // @[package.scala 93:22:@25071.4]
  wire  RetimeWrapper_156_reset; // @[package.scala 93:22:@25071.4]
  wire  RetimeWrapper_156_io_flow; // @[package.scala 93:22:@25071.4]
  wire  RetimeWrapper_156_io_in; // @[package.scala 93:22:@25071.4]
  wire  RetimeWrapper_156_io_out; // @[package.scala 93:22:@25071.4]
  wire  RetimeWrapper_157_clock; // @[package.scala 93:22:@25079.4]
  wire  RetimeWrapper_157_reset; // @[package.scala 93:22:@25079.4]
  wire  RetimeWrapper_157_io_flow; // @[package.scala 93:22:@25079.4]
  wire  RetimeWrapper_157_io_in; // @[package.scala 93:22:@25079.4]
  wire  RetimeWrapper_157_io_out; // @[package.scala 93:22:@25079.4]
  wire  RetimeWrapper_158_clock; // @[package.scala 93:22:@25087.4]
  wire  RetimeWrapper_158_reset; // @[package.scala 93:22:@25087.4]
  wire  RetimeWrapper_158_io_flow; // @[package.scala 93:22:@25087.4]
  wire  RetimeWrapper_158_io_in; // @[package.scala 93:22:@25087.4]
  wire  RetimeWrapper_158_io_out; // @[package.scala 93:22:@25087.4]
  wire  RetimeWrapper_159_clock; // @[package.scala 93:22:@25095.4]
  wire  RetimeWrapper_159_reset; // @[package.scala 93:22:@25095.4]
  wire  RetimeWrapper_159_io_flow; // @[package.scala 93:22:@25095.4]
  wire  RetimeWrapper_159_io_in; // @[package.scala 93:22:@25095.4]
  wire  RetimeWrapper_159_io_out; // @[package.scala 93:22:@25095.4]
  wire  RetimeWrapper_160_clock; // @[package.scala 93:22:@25103.4]
  wire  RetimeWrapper_160_reset; // @[package.scala 93:22:@25103.4]
  wire  RetimeWrapper_160_io_flow; // @[package.scala 93:22:@25103.4]
  wire  RetimeWrapper_160_io_in; // @[package.scala 93:22:@25103.4]
  wire  RetimeWrapper_160_io_out; // @[package.scala 93:22:@25103.4]
  wire  RetimeWrapper_161_clock; // @[package.scala 93:22:@25111.4]
  wire  RetimeWrapper_161_reset; // @[package.scala 93:22:@25111.4]
  wire  RetimeWrapper_161_io_flow; // @[package.scala 93:22:@25111.4]
  wire  RetimeWrapper_161_io_in; // @[package.scala 93:22:@25111.4]
  wire  RetimeWrapper_161_io_out; // @[package.scala 93:22:@25111.4]
  wire  RetimeWrapper_162_clock; // @[package.scala 93:22:@25119.4]
  wire  RetimeWrapper_162_reset; // @[package.scala 93:22:@25119.4]
  wire  RetimeWrapper_162_io_flow; // @[package.scala 93:22:@25119.4]
  wire  RetimeWrapper_162_io_in; // @[package.scala 93:22:@25119.4]
  wire  RetimeWrapper_162_io_out; // @[package.scala 93:22:@25119.4]
  wire  RetimeWrapper_163_clock; // @[package.scala 93:22:@25127.4]
  wire  RetimeWrapper_163_reset; // @[package.scala 93:22:@25127.4]
  wire  RetimeWrapper_163_io_flow; // @[package.scala 93:22:@25127.4]
  wire  RetimeWrapper_163_io_in; // @[package.scala 93:22:@25127.4]
  wire  RetimeWrapper_163_io_out; // @[package.scala 93:22:@25127.4]
  wire  RetimeWrapper_164_clock; // @[package.scala 93:22:@25135.4]
  wire  RetimeWrapper_164_reset; // @[package.scala 93:22:@25135.4]
  wire  RetimeWrapper_164_io_flow; // @[package.scala 93:22:@25135.4]
  wire  RetimeWrapper_164_io_in; // @[package.scala 93:22:@25135.4]
  wire  RetimeWrapper_164_io_out; // @[package.scala 93:22:@25135.4]
  wire  RetimeWrapper_165_clock; // @[package.scala 93:22:@25143.4]
  wire  RetimeWrapper_165_reset; // @[package.scala 93:22:@25143.4]
  wire  RetimeWrapper_165_io_flow; // @[package.scala 93:22:@25143.4]
  wire  RetimeWrapper_165_io_in; // @[package.scala 93:22:@25143.4]
  wire  RetimeWrapper_165_io_out; // @[package.scala 93:22:@25143.4]
  wire  RetimeWrapper_166_clock; // @[package.scala 93:22:@25151.4]
  wire  RetimeWrapper_166_reset; // @[package.scala 93:22:@25151.4]
  wire  RetimeWrapper_166_io_flow; // @[package.scala 93:22:@25151.4]
  wire  RetimeWrapper_166_io_in; // @[package.scala 93:22:@25151.4]
  wire  RetimeWrapper_166_io_out; // @[package.scala 93:22:@25151.4]
  wire  RetimeWrapper_167_clock; // @[package.scala 93:22:@25159.4]
  wire  RetimeWrapper_167_reset; // @[package.scala 93:22:@25159.4]
  wire  RetimeWrapper_167_io_flow; // @[package.scala 93:22:@25159.4]
  wire  RetimeWrapper_167_io_in; // @[package.scala 93:22:@25159.4]
  wire  RetimeWrapper_167_io_out; // @[package.scala 93:22:@25159.4]
  wire  RetimeWrapper_168_clock; // @[package.scala 93:22:@25215.4]
  wire  RetimeWrapper_168_reset; // @[package.scala 93:22:@25215.4]
  wire  RetimeWrapper_168_io_flow; // @[package.scala 93:22:@25215.4]
  wire  RetimeWrapper_168_io_in; // @[package.scala 93:22:@25215.4]
  wire  RetimeWrapper_168_io_out; // @[package.scala 93:22:@25215.4]
  wire  RetimeWrapper_169_clock; // @[package.scala 93:22:@25223.4]
  wire  RetimeWrapper_169_reset; // @[package.scala 93:22:@25223.4]
  wire  RetimeWrapper_169_io_flow; // @[package.scala 93:22:@25223.4]
  wire  RetimeWrapper_169_io_in; // @[package.scala 93:22:@25223.4]
  wire  RetimeWrapper_169_io_out; // @[package.scala 93:22:@25223.4]
  wire  RetimeWrapper_170_clock; // @[package.scala 93:22:@25231.4]
  wire  RetimeWrapper_170_reset; // @[package.scala 93:22:@25231.4]
  wire  RetimeWrapper_170_io_flow; // @[package.scala 93:22:@25231.4]
  wire  RetimeWrapper_170_io_in; // @[package.scala 93:22:@25231.4]
  wire  RetimeWrapper_170_io_out; // @[package.scala 93:22:@25231.4]
  wire  RetimeWrapper_171_clock; // @[package.scala 93:22:@25239.4]
  wire  RetimeWrapper_171_reset; // @[package.scala 93:22:@25239.4]
  wire  RetimeWrapper_171_io_flow; // @[package.scala 93:22:@25239.4]
  wire  RetimeWrapper_171_io_in; // @[package.scala 93:22:@25239.4]
  wire  RetimeWrapper_171_io_out; // @[package.scala 93:22:@25239.4]
  wire  RetimeWrapper_172_clock; // @[package.scala 93:22:@25247.4]
  wire  RetimeWrapper_172_reset; // @[package.scala 93:22:@25247.4]
  wire  RetimeWrapper_172_io_flow; // @[package.scala 93:22:@25247.4]
  wire  RetimeWrapper_172_io_in; // @[package.scala 93:22:@25247.4]
  wire  RetimeWrapper_172_io_out; // @[package.scala 93:22:@25247.4]
  wire  RetimeWrapper_173_clock; // @[package.scala 93:22:@25255.4]
  wire  RetimeWrapper_173_reset; // @[package.scala 93:22:@25255.4]
  wire  RetimeWrapper_173_io_flow; // @[package.scala 93:22:@25255.4]
  wire  RetimeWrapper_173_io_in; // @[package.scala 93:22:@25255.4]
  wire  RetimeWrapper_173_io_out; // @[package.scala 93:22:@25255.4]
  wire  RetimeWrapper_174_clock; // @[package.scala 93:22:@25263.4]
  wire  RetimeWrapper_174_reset; // @[package.scala 93:22:@25263.4]
  wire  RetimeWrapper_174_io_flow; // @[package.scala 93:22:@25263.4]
  wire  RetimeWrapper_174_io_in; // @[package.scala 93:22:@25263.4]
  wire  RetimeWrapper_174_io_out; // @[package.scala 93:22:@25263.4]
  wire  RetimeWrapper_175_clock; // @[package.scala 93:22:@25271.4]
  wire  RetimeWrapper_175_reset; // @[package.scala 93:22:@25271.4]
  wire  RetimeWrapper_175_io_flow; // @[package.scala 93:22:@25271.4]
  wire  RetimeWrapper_175_io_in; // @[package.scala 93:22:@25271.4]
  wire  RetimeWrapper_175_io_out; // @[package.scala 93:22:@25271.4]
  wire  RetimeWrapper_176_clock; // @[package.scala 93:22:@25279.4]
  wire  RetimeWrapper_176_reset; // @[package.scala 93:22:@25279.4]
  wire  RetimeWrapper_176_io_flow; // @[package.scala 93:22:@25279.4]
  wire  RetimeWrapper_176_io_in; // @[package.scala 93:22:@25279.4]
  wire  RetimeWrapper_176_io_out; // @[package.scala 93:22:@25279.4]
  wire  RetimeWrapper_177_clock; // @[package.scala 93:22:@25287.4]
  wire  RetimeWrapper_177_reset; // @[package.scala 93:22:@25287.4]
  wire  RetimeWrapper_177_io_flow; // @[package.scala 93:22:@25287.4]
  wire  RetimeWrapper_177_io_in; // @[package.scala 93:22:@25287.4]
  wire  RetimeWrapper_177_io_out; // @[package.scala 93:22:@25287.4]
  wire  RetimeWrapper_178_clock; // @[package.scala 93:22:@25295.4]
  wire  RetimeWrapper_178_reset; // @[package.scala 93:22:@25295.4]
  wire  RetimeWrapper_178_io_flow; // @[package.scala 93:22:@25295.4]
  wire  RetimeWrapper_178_io_in; // @[package.scala 93:22:@25295.4]
  wire  RetimeWrapper_178_io_out; // @[package.scala 93:22:@25295.4]
  wire  RetimeWrapper_179_clock; // @[package.scala 93:22:@25303.4]
  wire  RetimeWrapper_179_reset; // @[package.scala 93:22:@25303.4]
  wire  RetimeWrapper_179_io_flow; // @[package.scala 93:22:@25303.4]
  wire  RetimeWrapper_179_io_in; // @[package.scala 93:22:@25303.4]
  wire  RetimeWrapper_179_io_out; // @[package.scala 93:22:@25303.4]
  wire  RetimeWrapper_180_clock; // @[package.scala 93:22:@25359.4]
  wire  RetimeWrapper_180_reset; // @[package.scala 93:22:@25359.4]
  wire  RetimeWrapper_180_io_flow; // @[package.scala 93:22:@25359.4]
  wire  RetimeWrapper_180_io_in; // @[package.scala 93:22:@25359.4]
  wire  RetimeWrapper_180_io_out; // @[package.scala 93:22:@25359.4]
  wire  RetimeWrapper_181_clock; // @[package.scala 93:22:@25367.4]
  wire  RetimeWrapper_181_reset; // @[package.scala 93:22:@25367.4]
  wire  RetimeWrapper_181_io_flow; // @[package.scala 93:22:@25367.4]
  wire  RetimeWrapper_181_io_in; // @[package.scala 93:22:@25367.4]
  wire  RetimeWrapper_181_io_out; // @[package.scala 93:22:@25367.4]
  wire  RetimeWrapper_182_clock; // @[package.scala 93:22:@25375.4]
  wire  RetimeWrapper_182_reset; // @[package.scala 93:22:@25375.4]
  wire  RetimeWrapper_182_io_flow; // @[package.scala 93:22:@25375.4]
  wire  RetimeWrapper_182_io_in; // @[package.scala 93:22:@25375.4]
  wire  RetimeWrapper_182_io_out; // @[package.scala 93:22:@25375.4]
  wire  RetimeWrapper_183_clock; // @[package.scala 93:22:@25383.4]
  wire  RetimeWrapper_183_reset; // @[package.scala 93:22:@25383.4]
  wire  RetimeWrapper_183_io_flow; // @[package.scala 93:22:@25383.4]
  wire  RetimeWrapper_183_io_in; // @[package.scala 93:22:@25383.4]
  wire  RetimeWrapper_183_io_out; // @[package.scala 93:22:@25383.4]
  wire  RetimeWrapper_184_clock; // @[package.scala 93:22:@25391.4]
  wire  RetimeWrapper_184_reset; // @[package.scala 93:22:@25391.4]
  wire  RetimeWrapper_184_io_flow; // @[package.scala 93:22:@25391.4]
  wire  RetimeWrapper_184_io_in; // @[package.scala 93:22:@25391.4]
  wire  RetimeWrapper_184_io_out; // @[package.scala 93:22:@25391.4]
  wire  RetimeWrapper_185_clock; // @[package.scala 93:22:@25399.4]
  wire  RetimeWrapper_185_reset; // @[package.scala 93:22:@25399.4]
  wire  RetimeWrapper_185_io_flow; // @[package.scala 93:22:@25399.4]
  wire  RetimeWrapper_185_io_in; // @[package.scala 93:22:@25399.4]
  wire  RetimeWrapper_185_io_out; // @[package.scala 93:22:@25399.4]
  wire  RetimeWrapper_186_clock; // @[package.scala 93:22:@25407.4]
  wire  RetimeWrapper_186_reset; // @[package.scala 93:22:@25407.4]
  wire  RetimeWrapper_186_io_flow; // @[package.scala 93:22:@25407.4]
  wire  RetimeWrapper_186_io_in; // @[package.scala 93:22:@25407.4]
  wire  RetimeWrapper_186_io_out; // @[package.scala 93:22:@25407.4]
  wire  RetimeWrapper_187_clock; // @[package.scala 93:22:@25415.4]
  wire  RetimeWrapper_187_reset; // @[package.scala 93:22:@25415.4]
  wire  RetimeWrapper_187_io_flow; // @[package.scala 93:22:@25415.4]
  wire  RetimeWrapper_187_io_in; // @[package.scala 93:22:@25415.4]
  wire  RetimeWrapper_187_io_out; // @[package.scala 93:22:@25415.4]
  wire  RetimeWrapper_188_clock; // @[package.scala 93:22:@25423.4]
  wire  RetimeWrapper_188_reset; // @[package.scala 93:22:@25423.4]
  wire  RetimeWrapper_188_io_flow; // @[package.scala 93:22:@25423.4]
  wire  RetimeWrapper_188_io_in; // @[package.scala 93:22:@25423.4]
  wire  RetimeWrapper_188_io_out; // @[package.scala 93:22:@25423.4]
  wire  RetimeWrapper_189_clock; // @[package.scala 93:22:@25431.4]
  wire  RetimeWrapper_189_reset; // @[package.scala 93:22:@25431.4]
  wire  RetimeWrapper_189_io_flow; // @[package.scala 93:22:@25431.4]
  wire  RetimeWrapper_189_io_in; // @[package.scala 93:22:@25431.4]
  wire  RetimeWrapper_189_io_out; // @[package.scala 93:22:@25431.4]
  wire  RetimeWrapper_190_clock; // @[package.scala 93:22:@25439.4]
  wire  RetimeWrapper_190_reset; // @[package.scala 93:22:@25439.4]
  wire  RetimeWrapper_190_io_flow; // @[package.scala 93:22:@25439.4]
  wire  RetimeWrapper_190_io_in; // @[package.scala 93:22:@25439.4]
  wire  RetimeWrapper_190_io_out; // @[package.scala 93:22:@25439.4]
  wire  RetimeWrapper_191_clock; // @[package.scala 93:22:@25447.4]
  wire  RetimeWrapper_191_reset; // @[package.scala 93:22:@25447.4]
  wire  RetimeWrapper_191_io_flow; // @[package.scala 93:22:@25447.4]
  wire  RetimeWrapper_191_io_in; // @[package.scala 93:22:@25447.4]
  wire  RetimeWrapper_191_io_out; // @[package.scala 93:22:@25447.4]
  wire  RetimeWrapper_192_clock; // @[package.scala 93:22:@25503.4]
  wire  RetimeWrapper_192_reset; // @[package.scala 93:22:@25503.4]
  wire  RetimeWrapper_192_io_flow; // @[package.scala 93:22:@25503.4]
  wire  RetimeWrapper_192_io_in; // @[package.scala 93:22:@25503.4]
  wire  RetimeWrapper_192_io_out; // @[package.scala 93:22:@25503.4]
  wire  RetimeWrapper_193_clock; // @[package.scala 93:22:@25511.4]
  wire  RetimeWrapper_193_reset; // @[package.scala 93:22:@25511.4]
  wire  RetimeWrapper_193_io_flow; // @[package.scala 93:22:@25511.4]
  wire  RetimeWrapper_193_io_in; // @[package.scala 93:22:@25511.4]
  wire  RetimeWrapper_193_io_out; // @[package.scala 93:22:@25511.4]
  wire  RetimeWrapper_194_clock; // @[package.scala 93:22:@25519.4]
  wire  RetimeWrapper_194_reset; // @[package.scala 93:22:@25519.4]
  wire  RetimeWrapper_194_io_flow; // @[package.scala 93:22:@25519.4]
  wire  RetimeWrapper_194_io_in; // @[package.scala 93:22:@25519.4]
  wire  RetimeWrapper_194_io_out; // @[package.scala 93:22:@25519.4]
  wire  RetimeWrapper_195_clock; // @[package.scala 93:22:@25527.4]
  wire  RetimeWrapper_195_reset; // @[package.scala 93:22:@25527.4]
  wire  RetimeWrapper_195_io_flow; // @[package.scala 93:22:@25527.4]
  wire  RetimeWrapper_195_io_in; // @[package.scala 93:22:@25527.4]
  wire  RetimeWrapper_195_io_out; // @[package.scala 93:22:@25527.4]
  wire  RetimeWrapper_196_clock; // @[package.scala 93:22:@25535.4]
  wire  RetimeWrapper_196_reset; // @[package.scala 93:22:@25535.4]
  wire  RetimeWrapper_196_io_flow; // @[package.scala 93:22:@25535.4]
  wire  RetimeWrapper_196_io_in; // @[package.scala 93:22:@25535.4]
  wire  RetimeWrapper_196_io_out; // @[package.scala 93:22:@25535.4]
  wire  RetimeWrapper_197_clock; // @[package.scala 93:22:@25543.4]
  wire  RetimeWrapper_197_reset; // @[package.scala 93:22:@25543.4]
  wire  RetimeWrapper_197_io_flow; // @[package.scala 93:22:@25543.4]
  wire  RetimeWrapper_197_io_in; // @[package.scala 93:22:@25543.4]
  wire  RetimeWrapper_197_io_out; // @[package.scala 93:22:@25543.4]
  wire  RetimeWrapper_198_clock; // @[package.scala 93:22:@25551.4]
  wire  RetimeWrapper_198_reset; // @[package.scala 93:22:@25551.4]
  wire  RetimeWrapper_198_io_flow; // @[package.scala 93:22:@25551.4]
  wire  RetimeWrapper_198_io_in; // @[package.scala 93:22:@25551.4]
  wire  RetimeWrapper_198_io_out; // @[package.scala 93:22:@25551.4]
  wire  RetimeWrapper_199_clock; // @[package.scala 93:22:@25559.4]
  wire  RetimeWrapper_199_reset; // @[package.scala 93:22:@25559.4]
  wire  RetimeWrapper_199_io_flow; // @[package.scala 93:22:@25559.4]
  wire  RetimeWrapper_199_io_in; // @[package.scala 93:22:@25559.4]
  wire  RetimeWrapper_199_io_out; // @[package.scala 93:22:@25559.4]
  wire  RetimeWrapper_200_clock; // @[package.scala 93:22:@25567.4]
  wire  RetimeWrapper_200_reset; // @[package.scala 93:22:@25567.4]
  wire  RetimeWrapper_200_io_flow; // @[package.scala 93:22:@25567.4]
  wire  RetimeWrapper_200_io_in; // @[package.scala 93:22:@25567.4]
  wire  RetimeWrapper_200_io_out; // @[package.scala 93:22:@25567.4]
  wire  RetimeWrapper_201_clock; // @[package.scala 93:22:@25575.4]
  wire  RetimeWrapper_201_reset; // @[package.scala 93:22:@25575.4]
  wire  RetimeWrapper_201_io_flow; // @[package.scala 93:22:@25575.4]
  wire  RetimeWrapper_201_io_in; // @[package.scala 93:22:@25575.4]
  wire  RetimeWrapper_201_io_out; // @[package.scala 93:22:@25575.4]
  wire  RetimeWrapper_202_clock; // @[package.scala 93:22:@25583.4]
  wire  RetimeWrapper_202_reset; // @[package.scala 93:22:@25583.4]
  wire  RetimeWrapper_202_io_flow; // @[package.scala 93:22:@25583.4]
  wire  RetimeWrapper_202_io_in; // @[package.scala 93:22:@25583.4]
  wire  RetimeWrapper_202_io_out; // @[package.scala 93:22:@25583.4]
  wire  RetimeWrapper_203_clock; // @[package.scala 93:22:@25591.4]
  wire  RetimeWrapper_203_reset; // @[package.scala 93:22:@25591.4]
  wire  RetimeWrapper_203_io_flow; // @[package.scala 93:22:@25591.4]
  wire  RetimeWrapper_203_io_in; // @[package.scala 93:22:@25591.4]
  wire  RetimeWrapper_203_io_out; // @[package.scala 93:22:@25591.4]
  wire  RetimeWrapper_204_clock; // @[package.scala 93:22:@25647.4]
  wire  RetimeWrapper_204_reset; // @[package.scala 93:22:@25647.4]
  wire  RetimeWrapper_204_io_flow; // @[package.scala 93:22:@25647.4]
  wire  RetimeWrapper_204_io_in; // @[package.scala 93:22:@25647.4]
  wire  RetimeWrapper_204_io_out; // @[package.scala 93:22:@25647.4]
  wire  RetimeWrapper_205_clock; // @[package.scala 93:22:@25655.4]
  wire  RetimeWrapper_205_reset; // @[package.scala 93:22:@25655.4]
  wire  RetimeWrapper_205_io_flow; // @[package.scala 93:22:@25655.4]
  wire  RetimeWrapper_205_io_in; // @[package.scala 93:22:@25655.4]
  wire  RetimeWrapper_205_io_out; // @[package.scala 93:22:@25655.4]
  wire  RetimeWrapper_206_clock; // @[package.scala 93:22:@25663.4]
  wire  RetimeWrapper_206_reset; // @[package.scala 93:22:@25663.4]
  wire  RetimeWrapper_206_io_flow; // @[package.scala 93:22:@25663.4]
  wire  RetimeWrapper_206_io_in; // @[package.scala 93:22:@25663.4]
  wire  RetimeWrapper_206_io_out; // @[package.scala 93:22:@25663.4]
  wire  RetimeWrapper_207_clock; // @[package.scala 93:22:@25671.4]
  wire  RetimeWrapper_207_reset; // @[package.scala 93:22:@25671.4]
  wire  RetimeWrapper_207_io_flow; // @[package.scala 93:22:@25671.4]
  wire  RetimeWrapper_207_io_in; // @[package.scala 93:22:@25671.4]
  wire  RetimeWrapper_207_io_out; // @[package.scala 93:22:@25671.4]
  wire  RetimeWrapper_208_clock; // @[package.scala 93:22:@25679.4]
  wire  RetimeWrapper_208_reset; // @[package.scala 93:22:@25679.4]
  wire  RetimeWrapper_208_io_flow; // @[package.scala 93:22:@25679.4]
  wire  RetimeWrapper_208_io_in; // @[package.scala 93:22:@25679.4]
  wire  RetimeWrapper_208_io_out; // @[package.scala 93:22:@25679.4]
  wire  RetimeWrapper_209_clock; // @[package.scala 93:22:@25687.4]
  wire  RetimeWrapper_209_reset; // @[package.scala 93:22:@25687.4]
  wire  RetimeWrapper_209_io_flow; // @[package.scala 93:22:@25687.4]
  wire  RetimeWrapper_209_io_in; // @[package.scala 93:22:@25687.4]
  wire  RetimeWrapper_209_io_out; // @[package.scala 93:22:@25687.4]
  wire  RetimeWrapper_210_clock; // @[package.scala 93:22:@25695.4]
  wire  RetimeWrapper_210_reset; // @[package.scala 93:22:@25695.4]
  wire  RetimeWrapper_210_io_flow; // @[package.scala 93:22:@25695.4]
  wire  RetimeWrapper_210_io_in; // @[package.scala 93:22:@25695.4]
  wire  RetimeWrapper_210_io_out; // @[package.scala 93:22:@25695.4]
  wire  RetimeWrapper_211_clock; // @[package.scala 93:22:@25703.4]
  wire  RetimeWrapper_211_reset; // @[package.scala 93:22:@25703.4]
  wire  RetimeWrapper_211_io_flow; // @[package.scala 93:22:@25703.4]
  wire  RetimeWrapper_211_io_in; // @[package.scala 93:22:@25703.4]
  wire  RetimeWrapper_211_io_out; // @[package.scala 93:22:@25703.4]
  wire  RetimeWrapper_212_clock; // @[package.scala 93:22:@25711.4]
  wire  RetimeWrapper_212_reset; // @[package.scala 93:22:@25711.4]
  wire  RetimeWrapper_212_io_flow; // @[package.scala 93:22:@25711.4]
  wire  RetimeWrapper_212_io_in; // @[package.scala 93:22:@25711.4]
  wire  RetimeWrapper_212_io_out; // @[package.scala 93:22:@25711.4]
  wire  RetimeWrapper_213_clock; // @[package.scala 93:22:@25719.4]
  wire  RetimeWrapper_213_reset; // @[package.scala 93:22:@25719.4]
  wire  RetimeWrapper_213_io_flow; // @[package.scala 93:22:@25719.4]
  wire  RetimeWrapper_213_io_in; // @[package.scala 93:22:@25719.4]
  wire  RetimeWrapper_213_io_out; // @[package.scala 93:22:@25719.4]
  wire  RetimeWrapper_214_clock; // @[package.scala 93:22:@25727.4]
  wire  RetimeWrapper_214_reset; // @[package.scala 93:22:@25727.4]
  wire  RetimeWrapper_214_io_flow; // @[package.scala 93:22:@25727.4]
  wire  RetimeWrapper_214_io_in; // @[package.scala 93:22:@25727.4]
  wire  RetimeWrapper_214_io_out; // @[package.scala 93:22:@25727.4]
  wire  RetimeWrapper_215_clock; // @[package.scala 93:22:@25735.4]
  wire  RetimeWrapper_215_reset; // @[package.scala 93:22:@25735.4]
  wire  RetimeWrapper_215_io_flow; // @[package.scala 93:22:@25735.4]
  wire  RetimeWrapper_215_io_in; // @[package.scala 93:22:@25735.4]
  wire  RetimeWrapper_215_io_out; // @[package.scala 93:22:@25735.4]
  wire  _T_700; // @[MemPrimitives.scala 82:210:@20570.4]
  wire  _T_702; // @[MemPrimitives.scala 82:210:@20571.4]
  wire  _T_703; // @[MemPrimitives.scala 82:228:@20572.4]
  wire  _T_704; // @[MemPrimitives.scala 83:102:@20573.4]
  wire  _T_706; // @[MemPrimitives.scala 82:210:@20574.4]
  wire  _T_708; // @[MemPrimitives.scala 82:210:@20575.4]
  wire  _T_709; // @[MemPrimitives.scala 82:228:@20576.4]
  wire  _T_710; // @[MemPrimitives.scala 83:102:@20577.4]
  wire [41:0] _T_712; // @[Cat.scala 30:58:@20579.4]
  wire [41:0] _T_714; // @[Cat.scala 30:58:@20581.4]
  wire [41:0] _T_715; // @[Mux.scala 31:69:@20582.4]
  wire  _T_720; // @[MemPrimitives.scala 82:210:@20589.4]
  wire  _T_722; // @[MemPrimitives.scala 82:210:@20590.4]
  wire  _T_723; // @[MemPrimitives.scala 82:228:@20591.4]
  wire  _T_724; // @[MemPrimitives.scala 83:102:@20592.4]
  wire  _T_726; // @[MemPrimitives.scala 82:210:@20593.4]
  wire  _T_728; // @[MemPrimitives.scala 82:210:@20594.4]
  wire  _T_729; // @[MemPrimitives.scala 82:228:@20595.4]
  wire  _T_730; // @[MemPrimitives.scala 83:102:@20596.4]
  wire [41:0] _T_732; // @[Cat.scala 30:58:@20598.4]
  wire [41:0] _T_734; // @[Cat.scala 30:58:@20600.4]
  wire [41:0] _T_735; // @[Mux.scala 31:69:@20601.4]
  wire  _T_742; // @[MemPrimitives.scala 82:210:@20609.4]
  wire  _T_743; // @[MemPrimitives.scala 82:228:@20610.4]
  wire  _T_744; // @[MemPrimitives.scala 83:102:@20611.4]
  wire  _T_748; // @[MemPrimitives.scala 82:210:@20613.4]
  wire  _T_749; // @[MemPrimitives.scala 82:228:@20614.4]
  wire  _T_750; // @[MemPrimitives.scala 83:102:@20615.4]
  wire [41:0] _T_752; // @[Cat.scala 30:58:@20617.4]
  wire [41:0] _T_754; // @[Cat.scala 30:58:@20619.4]
  wire [41:0] _T_755; // @[Mux.scala 31:69:@20620.4]
  wire  _T_762; // @[MemPrimitives.scala 82:210:@20628.4]
  wire  _T_763; // @[MemPrimitives.scala 82:228:@20629.4]
  wire  _T_764; // @[MemPrimitives.scala 83:102:@20630.4]
  wire  _T_768; // @[MemPrimitives.scala 82:210:@20632.4]
  wire  _T_769; // @[MemPrimitives.scala 82:228:@20633.4]
  wire  _T_770; // @[MemPrimitives.scala 83:102:@20634.4]
  wire [41:0] _T_772; // @[Cat.scala 30:58:@20636.4]
  wire [41:0] _T_774; // @[Cat.scala 30:58:@20638.4]
  wire [41:0] _T_775; // @[Mux.scala 31:69:@20639.4]
  wire  _T_782; // @[MemPrimitives.scala 82:210:@20647.4]
  wire  _T_783; // @[MemPrimitives.scala 82:228:@20648.4]
  wire  _T_784; // @[MemPrimitives.scala 83:102:@20649.4]
  wire  _T_788; // @[MemPrimitives.scala 82:210:@20651.4]
  wire  _T_789; // @[MemPrimitives.scala 82:228:@20652.4]
  wire  _T_790; // @[MemPrimitives.scala 83:102:@20653.4]
  wire [41:0] _T_792; // @[Cat.scala 30:58:@20655.4]
  wire [41:0] _T_794; // @[Cat.scala 30:58:@20657.4]
  wire [41:0] _T_795; // @[Mux.scala 31:69:@20658.4]
  wire  _T_802; // @[MemPrimitives.scala 82:210:@20666.4]
  wire  _T_803; // @[MemPrimitives.scala 82:228:@20667.4]
  wire  _T_804; // @[MemPrimitives.scala 83:102:@20668.4]
  wire  _T_808; // @[MemPrimitives.scala 82:210:@20670.4]
  wire  _T_809; // @[MemPrimitives.scala 82:228:@20671.4]
  wire  _T_810; // @[MemPrimitives.scala 83:102:@20672.4]
  wire [41:0] _T_812; // @[Cat.scala 30:58:@20674.4]
  wire [41:0] _T_814; // @[Cat.scala 30:58:@20676.4]
  wire [41:0] _T_815; // @[Mux.scala 31:69:@20677.4]
  wire  _T_820; // @[MemPrimitives.scala 82:210:@20684.4]
  wire  _T_823; // @[MemPrimitives.scala 82:228:@20686.4]
  wire  _T_824; // @[MemPrimitives.scala 83:102:@20687.4]
  wire  _T_826; // @[MemPrimitives.scala 82:210:@20688.4]
  wire  _T_829; // @[MemPrimitives.scala 82:228:@20690.4]
  wire  _T_830; // @[MemPrimitives.scala 83:102:@20691.4]
  wire [41:0] _T_832; // @[Cat.scala 30:58:@20693.4]
  wire [41:0] _T_834; // @[Cat.scala 30:58:@20695.4]
  wire [41:0] _T_835; // @[Mux.scala 31:69:@20696.4]
  wire  _T_840; // @[MemPrimitives.scala 82:210:@20703.4]
  wire  _T_843; // @[MemPrimitives.scala 82:228:@20705.4]
  wire  _T_844; // @[MemPrimitives.scala 83:102:@20706.4]
  wire  _T_846; // @[MemPrimitives.scala 82:210:@20707.4]
  wire  _T_849; // @[MemPrimitives.scala 82:228:@20709.4]
  wire  _T_850; // @[MemPrimitives.scala 83:102:@20710.4]
  wire [41:0] _T_852; // @[Cat.scala 30:58:@20712.4]
  wire [41:0] _T_854; // @[Cat.scala 30:58:@20714.4]
  wire [41:0] _T_855; // @[Mux.scala 31:69:@20715.4]
  wire  _T_863; // @[MemPrimitives.scala 82:228:@20724.4]
  wire  _T_864; // @[MemPrimitives.scala 83:102:@20725.4]
  wire  _T_869; // @[MemPrimitives.scala 82:228:@20728.4]
  wire  _T_870; // @[MemPrimitives.scala 83:102:@20729.4]
  wire [41:0] _T_872; // @[Cat.scala 30:58:@20731.4]
  wire [41:0] _T_874; // @[Cat.scala 30:58:@20733.4]
  wire [41:0] _T_875; // @[Mux.scala 31:69:@20734.4]
  wire  _T_883; // @[MemPrimitives.scala 82:228:@20743.4]
  wire  _T_884; // @[MemPrimitives.scala 83:102:@20744.4]
  wire  _T_889; // @[MemPrimitives.scala 82:228:@20747.4]
  wire  _T_890; // @[MemPrimitives.scala 83:102:@20748.4]
  wire [41:0] _T_892; // @[Cat.scala 30:58:@20750.4]
  wire [41:0] _T_894; // @[Cat.scala 30:58:@20752.4]
  wire [41:0] _T_895; // @[Mux.scala 31:69:@20753.4]
  wire  _T_903; // @[MemPrimitives.scala 82:228:@20762.4]
  wire  _T_904; // @[MemPrimitives.scala 83:102:@20763.4]
  wire  _T_909; // @[MemPrimitives.scala 82:228:@20766.4]
  wire  _T_910; // @[MemPrimitives.scala 83:102:@20767.4]
  wire [41:0] _T_912; // @[Cat.scala 30:58:@20769.4]
  wire [41:0] _T_914; // @[Cat.scala 30:58:@20771.4]
  wire [41:0] _T_915; // @[Mux.scala 31:69:@20772.4]
  wire  _T_923; // @[MemPrimitives.scala 82:228:@20781.4]
  wire  _T_924; // @[MemPrimitives.scala 83:102:@20782.4]
  wire  _T_929; // @[MemPrimitives.scala 82:228:@20785.4]
  wire  _T_930; // @[MemPrimitives.scala 83:102:@20786.4]
  wire [41:0] _T_932; // @[Cat.scala 30:58:@20788.4]
  wire [41:0] _T_934; // @[Cat.scala 30:58:@20790.4]
  wire [41:0] _T_935; // @[Mux.scala 31:69:@20791.4]
  wire  _T_940; // @[MemPrimitives.scala 82:210:@20798.4]
  wire  _T_943; // @[MemPrimitives.scala 82:228:@20800.4]
  wire  _T_944; // @[MemPrimitives.scala 83:102:@20801.4]
  wire  _T_946; // @[MemPrimitives.scala 82:210:@20802.4]
  wire  _T_949; // @[MemPrimitives.scala 82:228:@20804.4]
  wire  _T_950; // @[MemPrimitives.scala 83:102:@20805.4]
  wire [41:0] _T_952; // @[Cat.scala 30:58:@20807.4]
  wire [41:0] _T_954; // @[Cat.scala 30:58:@20809.4]
  wire [41:0] _T_955; // @[Mux.scala 31:69:@20810.4]
  wire  _T_960; // @[MemPrimitives.scala 82:210:@20817.4]
  wire  _T_963; // @[MemPrimitives.scala 82:228:@20819.4]
  wire  _T_964; // @[MemPrimitives.scala 83:102:@20820.4]
  wire  _T_966; // @[MemPrimitives.scala 82:210:@20821.4]
  wire  _T_969; // @[MemPrimitives.scala 82:228:@20823.4]
  wire  _T_970; // @[MemPrimitives.scala 83:102:@20824.4]
  wire [41:0] _T_972; // @[Cat.scala 30:58:@20826.4]
  wire [41:0] _T_974; // @[Cat.scala 30:58:@20828.4]
  wire [41:0] _T_975; // @[Mux.scala 31:69:@20829.4]
  wire  _T_983; // @[MemPrimitives.scala 82:228:@20838.4]
  wire  _T_984; // @[MemPrimitives.scala 83:102:@20839.4]
  wire  _T_989; // @[MemPrimitives.scala 82:228:@20842.4]
  wire  _T_990; // @[MemPrimitives.scala 83:102:@20843.4]
  wire [41:0] _T_992; // @[Cat.scala 30:58:@20845.4]
  wire [41:0] _T_994; // @[Cat.scala 30:58:@20847.4]
  wire [41:0] _T_995; // @[Mux.scala 31:69:@20848.4]
  wire  _T_1003; // @[MemPrimitives.scala 82:228:@20857.4]
  wire  _T_1004; // @[MemPrimitives.scala 83:102:@20858.4]
  wire  _T_1009; // @[MemPrimitives.scala 82:228:@20861.4]
  wire  _T_1010; // @[MemPrimitives.scala 83:102:@20862.4]
  wire [41:0] _T_1012; // @[Cat.scala 30:58:@20864.4]
  wire [41:0] _T_1014; // @[Cat.scala 30:58:@20866.4]
  wire [41:0] _T_1015; // @[Mux.scala 31:69:@20867.4]
  wire  _T_1023; // @[MemPrimitives.scala 82:228:@20876.4]
  wire  _T_1024; // @[MemPrimitives.scala 83:102:@20877.4]
  wire  _T_1029; // @[MemPrimitives.scala 82:228:@20880.4]
  wire  _T_1030; // @[MemPrimitives.scala 83:102:@20881.4]
  wire [41:0] _T_1032; // @[Cat.scala 30:58:@20883.4]
  wire [41:0] _T_1034; // @[Cat.scala 30:58:@20885.4]
  wire [41:0] _T_1035; // @[Mux.scala 31:69:@20886.4]
  wire  _T_1043; // @[MemPrimitives.scala 82:228:@20895.4]
  wire  _T_1044; // @[MemPrimitives.scala 83:102:@20896.4]
  wire  _T_1049; // @[MemPrimitives.scala 82:228:@20899.4]
  wire  _T_1050; // @[MemPrimitives.scala 83:102:@20900.4]
  wire [41:0] _T_1052; // @[Cat.scala 30:58:@20902.4]
  wire [41:0] _T_1054; // @[Cat.scala 30:58:@20904.4]
  wire [41:0] _T_1055; // @[Mux.scala 31:69:@20905.4]
  wire  _T_1060; // @[MemPrimitives.scala 82:210:@20912.4]
  wire  _T_1063; // @[MemPrimitives.scala 82:228:@20914.4]
  wire  _T_1064; // @[MemPrimitives.scala 83:102:@20915.4]
  wire  _T_1066; // @[MemPrimitives.scala 82:210:@20916.4]
  wire  _T_1069; // @[MemPrimitives.scala 82:228:@20918.4]
  wire  _T_1070; // @[MemPrimitives.scala 83:102:@20919.4]
  wire [41:0] _T_1072; // @[Cat.scala 30:58:@20921.4]
  wire [41:0] _T_1074; // @[Cat.scala 30:58:@20923.4]
  wire [41:0] _T_1075; // @[Mux.scala 31:69:@20924.4]
  wire  _T_1080; // @[MemPrimitives.scala 82:210:@20931.4]
  wire  _T_1083; // @[MemPrimitives.scala 82:228:@20933.4]
  wire  _T_1084; // @[MemPrimitives.scala 83:102:@20934.4]
  wire  _T_1086; // @[MemPrimitives.scala 82:210:@20935.4]
  wire  _T_1089; // @[MemPrimitives.scala 82:228:@20937.4]
  wire  _T_1090; // @[MemPrimitives.scala 83:102:@20938.4]
  wire [41:0] _T_1092; // @[Cat.scala 30:58:@20940.4]
  wire [41:0] _T_1094; // @[Cat.scala 30:58:@20942.4]
  wire [41:0] _T_1095; // @[Mux.scala 31:69:@20943.4]
  wire  _T_1103; // @[MemPrimitives.scala 82:228:@20952.4]
  wire  _T_1104; // @[MemPrimitives.scala 83:102:@20953.4]
  wire  _T_1109; // @[MemPrimitives.scala 82:228:@20956.4]
  wire  _T_1110; // @[MemPrimitives.scala 83:102:@20957.4]
  wire [41:0] _T_1112; // @[Cat.scala 30:58:@20959.4]
  wire [41:0] _T_1114; // @[Cat.scala 30:58:@20961.4]
  wire [41:0] _T_1115; // @[Mux.scala 31:69:@20962.4]
  wire  _T_1123; // @[MemPrimitives.scala 82:228:@20971.4]
  wire  _T_1124; // @[MemPrimitives.scala 83:102:@20972.4]
  wire  _T_1129; // @[MemPrimitives.scala 82:228:@20975.4]
  wire  _T_1130; // @[MemPrimitives.scala 83:102:@20976.4]
  wire [41:0] _T_1132; // @[Cat.scala 30:58:@20978.4]
  wire [41:0] _T_1134; // @[Cat.scala 30:58:@20980.4]
  wire [41:0] _T_1135; // @[Mux.scala 31:69:@20981.4]
  wire  _T_1143; // @[MemPrimitives.scala 82:228:@20990.4]
  wire  _T_1144; // @[MemPrimitives.scala 83:102:@20991.4]
  wire  _T_1149; // @[MemPrimitives.scala 82:228:@20994.4]
  wire  _T_1150; // @[MemPrimitives.scala 83:102:@20995.4]
  wire [41:0] _T_1152; // @[Cat.scala 30:58:@20997.4]
  wire [41:0] _T_1154; // @[Cat.scala 30:58:@20999.4]
  wire [41:0] _T_1155; // @[Mux.scala 31:69:@21000.4]
  wire  _T_1163; // @[MemPrimitives.scala 82:228:@21009.4]
  wire  _T_1164; // @[MemPrimitives.scala 83:102:@21010.4]
  wire  _T_1169; // @[MemPrimitives.scala 82:228:@21013.4]
  wire  _T_1170; // @[MemPrimitives.scala 83:102:@21014.4]
  wire [41:0] _T_1172; // @[Cat.scala 30:58:@21016.4]
  wire [41:0] _T_1174; // @[Cat.scala 30:58:@21018.4]
  wire [41:0] _T_1175; // @[Mux.scala 31:69:@21019.4]
  wire  _T_1180; // @[MemPrimitives.scala 110:210:@21026.4]
  wire  _T_1182; // @[MemPrimitives.scala 110:210:@21027.4]
  wire  _T_1183; // @[MemPrimitives.scala 110:228:@21028.4]
  wire  _T_1186; // @[MemPrimitives.scala 110:210:@21030.4]
  wire  _T_1188; // @[MemPrimitives.scala 110:210:@21031.4]
  wire  _T_1189; // @[MemPrimitives.scala 110:228:@21032.4]
  wire  _T_1192; // @[MemPrimitives.scala 110:210:@21034.4]
  wire  _T_1194; // @[MemPrimitives.scala 110:210:@21035.4]
  wire  _T_1195; // @[MemPrimitives.scala 110:228:@21036.4]
  wire  _T_1198; // @[MemPrimitives.scala 110:210:@21038.4]
  wire  _T_1200; // @[MemPrimitives.scala 110:210:@21039.4]
  wire  _T_1201; // @[MemPrimitives.scala 110:228:@21040.4]
  wire  _T_1204; // @[MemPrimitives.scala 110:210:@21042.4]
  wire  _T_1206; // @[MemPrimitives.scala 110:210:@21043.4]
  wire  _T_1207; // @[MemPrimitives.scala 110:228:@21044.4]
  wire  _T_1210; // @[MemPrimitives.scala 110:210:@21046.4]
  wire  _T_1212; // @[MemPrimitives.scala 110:210:@21047.4]
  wire  _T_1213; // @[MemPrimitives.scala 110:228:@21048.4]
  wire  _T_1216; // @[MemPrimitives.scala 110:210:@21050.4]
  wire  _T_1218; // @[MemPrimitives.scala 110:210:@21051.4]
  wire  _T_1219; // @[MemPrimitives.scala 110:228:@21052.4]
  wire  _T_1222; // @[MemPrimitives.scala 110:210:@21054.4]
  wire  _T_1224; // @[MemPrimitives.scala 110:210:@21055.4]
  wire  _T_1225; // @[MemPrimitives.scala 110:228:@21056.4]
  wire  _T_1228; // @[MemPrimitives.scala 110:210:@21058.4]
  wire  _T_1230; // @[MemPrimitives.scala 110:210:@21059.4]
  wire  _T_1231; // @[MemPrimitives.scala 110:228:@21060.4]
  wire  _T_1233; // @[MemPrimitives.scala 126:35:@21074.4]
  wire  _T_1234; // @[MemPrimitives.scala 126:35:@21075.4]
  wire  _T_1235; // @[MemPrimitives.scala 126:35:@21076.4]
  wire  _T_1236; // @[MemPrimitives.scala 126:35:@21077.4]
  wire  _T_1237; // @[MemPrimitives.scala 126:35:@21078.4]
  wire  _T_1238; // @[MemPrimitives.scala 126:35:@21079.4]
  wire  _T_1239; // @[MemPrimitives.scala 126:35:@21080.4]
  wire  _T_1240; // @[MemPrimitives.scala 126:35:@21081.4]
  wire  _T_1241; // @[MemPrimitives.scala 126:35:@21082.4]
  wire [10:0] _T_1243; // @[Cat.scala 30:58:@21084.4]
  wire [10:0] _T_1245; // @[Cat.scala 30:58:@21086.4]
  wire [10:0] _T_1247; // @[Cat.scala 30:58:@21088.4]
  wire [10:0] _T_1249; // @[Cat.scala 30:58:@21090.4]
  wire [10:0] _T_1251; // @[Cat.scala 30:58:@21092.4]
  wire [10:0] _T_1253; // @[Cat.scala 30:58:@21094.4]
  wire [10:0] _T_1255; // @[Cat.scala 30:58:@21096.4]
  wire [10:0] _T_1257; // @[Cat.scala 30:58:@21098.4]
  wire [10:0] _T_1259; // @[Cat.scala 30:58:@21100.4]
  wire [10:0] _T_1260; // @[Mux.scala 31:69:@21101.4]
  wire [10:0] _T_1261; // @[Mux.scala 31:69:@21102.4]
  wire [10:0] _T_1262; // @[Mux.scala 31:69:@21103.4]
  wire [10:0] _T_1263; // @[Mux.scala 31:69:@21104.4]
  wire [10:0] _T_1264; // @[Mux.scala 31:69:@21105.4]
  wire [10:0] _T_1265; // @[Mux.scala 31:69:@21106.4]
  wire [10:0] _T_1266; // @[Mux.scala 31:69:@21107.4]
  wire [10:0] _T_1267; // @[Mux.scala 31:69:@21108.4]
  wire  _T_1272; // @[MemPrimitives.scala 110:210:@21115.4]
  wire  _T_1274; // @[MemPrimitives.scala 110:210:@21116.4]
  wire  _T_1275; // @[MemPrimitives.scala 110:228:@21117.4]
  wire  _T_1278; // @[MemPrimitives.scala 110:210:@21119.4]
  wire  _T_1280; // @[MemPrimitives.scala 110:210:@21120.4]
  wire  _T_1281; // @[MemPrimitives.scala 110:228:@21121.4]
  wire  _T_1284; // @[MemPrimitives.scala 110:210:@21123.4]
  wire  _T_1286; // @[MemPrimitives.scala 110:210:@21124.4]
  wire  _T_1287; // @[MemPrimitives.scala 110:228:@21125.4]
  wire  _T_1290; // @[MemPrimitives.scala 110:210:@21127.4]
  wire  _T_1292; // @[MemPrimitives.scala 110:210:@21128.4]
  wire  _T_1293; // @[MemPrimitives.scala 110:228:@21129.4]
  wire  _T_1296; // @[MemPrimitives.scala 110:210:@21131.4]
  wire  _T_1298; // @[MemPrimitives.scala 110:210:@21132.4]
  wire  _T_1299; // @[MemPrimitives.scala 110:228:@21133.4]
  wire  _T_1302; // @[MemPrimitives.scala 110:210:@21135.4]
  wire  _T_1304; // @[MemPrimitives.scala 110:210:@21136.4]
  wire  _T_1305; // @[MemPrimitives.scala 110:228:@21137.4]
  wire  _T_1308; // @[MemPrimitives.scala 110:210:@21139.4]
  wire  _T_1310; // @[MemPrimitives.scala 110:210:@21140.4]
  wire  _T_1311; // @[MemPrimitives.scala 110:228:@21141.4]
  wire  _T_1314; // @[MemPrimitives.scala 110:210:@21143.4]
  wire  _T_1316; // @[MemPrimitives.scala 110:210:@21144.4]
  wire  _T_1317; // @[MemPrimitives.scala 110:228:@21145.4]
  wire  _T_1320; // @[MemPrimitives.scala 110:210:@21147.4]
  wire  _T_1322; // @[MemPrimitives.scala 110:210:@21148.4]
  wire  _T_1323; // @[MemPrimitives.scala 110:228:@21149.4]
  wire  _T_1325; // @[MemPrimitives.scala 126:35:@21163.4]
  wire  _T_1326; // @[MemPrimitives.scala 126:35:@21164.4]
  wire  _T_1327; // @[MemPrimitives.scala 126:35:@21165.4]
  wire  _T_1328; // @[MemPrimitives.scala 126:35:@21166.4]
  wire  _T_1329; // @[MemPrimitives.scala 126:35:@21167.4]
  wire  _T_1330; // @[MemPrimitives.scala 126:35:@21168.4]
  wire  _T_1331; // @[MemPrimitives.scala 126:35:@21169.4]
  wire  _T_1332; // @[MemPrimitives.scala 126:35:@21170.4]
  wire  _T_1333; // @[MemPrimitives.scala 126:35:@21171.4]
  wire [10:0] _T_1335; // @[Cat.scala 30:58:@21173.4]
  wire [10:0] _T_1337; // @[Cat.scala 30:58:@21175.4]
  wire [10:0] _T_1339; // @[Cat.scala 30:58:@21177.4]
  wire [10:0] _T_1341; // @[Cat.scala 30:58:@21179.4]
  wire [10:0] _T_1343; // @[Cat.scala 30:58:@21181.4]
  wire [10:0] _T_1345; // @[Cat.scala 30:58:@21183.4]
  wire [10:0] _T_1347; // @[Cat.scala 30:58:@21185.4]
  wire [10:0] _T_1349; // @[Cat.scala 30:58:@21187.4]
  wire [10:0] _T_1351; // @[Cat.scala 30:58:@21189.4]
  wire [10:0] _T_1352; // @[Mux.scala 31:69:@21190.4]
  wire [10:0] _T_1353; // @[Mux.scala 31:69:@21191.4]
  wire [10:0] _T_1354; // @[Mux.scala 31:69:@21192.4]
  wire [10:0] _T_1355; // @[Mux.scala 31:69:@21193.4]
  wire [10:0] _T_1356; // @[Mux.scala 31:69:@21194.4]
  wire [10:0] _T_1357; // @[Mux.scala 31:69:@21195.4]
  wire [10:0] _T_1358; // @[Mux.scala 31:69:@21196.4]
  wire [10:0] _T_1359; // @[Mux.scala 31:69:@21197.4]
  wire  _T_1366; // @[MemPrimitives.scala 110:210:@21205.4]
  wire  _T_1367; // @[MemPrimitives.scala 110:228:@21206.4]
  wire  _T_1372; // @[MemPrimitives.scala 110:210:@21209.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:228:@21210.4]
  wire  _T_1378; // @[MemPrimitives.scala 110:210:@21213.4]
  wire  _T_1379; // @[MemPrimitives.scala 110:228:@21214.4]
  wire  _T_1384; // @[MemPrimitives.scala 110:210:@21217.4]
  wire  _T_1385; // @[MemPrimitives.scala 110:228:@21218.4]
  wire  _T_1390; // @[MemPrimitives.scala 110:210:@21221.4]
  wire  _T_1391; // @[MemPrimitives.scala 110:228:@21222.4]
  wire  _T_1396; // @[MemPrimitives.scala 110:210:@21225.4]
  wire  _T_1397; // @[MemPrimitives.scala 110:228:@21226.4]
  wire  _T_1402; // @[MemPrimitives.scala 110:210:@21229.4]
  wire  _T_1403; // @[MemPrimitives.scala 110:228:@21230.4]
  wire  _T_1408; // @[MemPrimitives.scala 110:210:@21233.4]
  wire  _T_1409; // @[MemPrimitives.scala 110:228:@21234.4]
  wire  _T_1414; // @[MemPrimitives.scala 110:210:@21237.4]
  wire  _T_1415; // @[MemPrimitives.scala 110:228:@21238.4]
  wire  _T_1417; // @[MemPrimitives.scala 126:35:@21252.4]
  wire  _T_1418; // @[MemPrimitives.scala 126:35:@21253.4]
  wire  _T_1419; // @[MemPrimitives.scala 126:35:@21254.4]
  wire  _T_1420; // @[MemPrimitives.scala 126:35:@21255.4]
  wire  _T_1421; // @[MemPrimitives.scala 126:35:@21256.4]
  wire  _T_1422; // @[MemPrimitives.scala 126:35:@21257.4]
  wire  _T_1423; // @[MemPrimitives.scala 126:35:@21258.4]
  wire  _T_1424; // @[MemPrimitives.scala 126:35:@21259.4]
  wire  _T_1425; // @[MemPrimitives.scala 126:35:@21260.4]
  wire [10:0] _T_1427; // @[Cat.scala 30:58:@21262.4]
  wire [10:0] _T_1429; // @[Cat.scala 30:58:@21264.4]
  wire [10:0] _T_1431; // @[Cat.scala 30:58:@21266.4]
  wire [10:0] _T_1433; // @[Cat.scala 30:58:@21268.4]
  wire [10:0] _T_1435; // @[Cat.scala 30:58:@21270.4]
  wire [10:0] _T_1437; // @[Cat.scala 30:58:@21272.4]
  wire [10:0] _T_1439; // @[Cat.scala 30:58:@21274.4]
  wire [10:0] _T_1441; // @[Cat.scala 30:58:@21276.4]
  wire [10:0] _T_1443; // @[Cat.scala 30:58:@21278.4]
  wire [10:0] _T_1444; // @[Mux.scala 31:69:@21279.4]
  wire [10:0] _T_1445; // @[Mux.scala 31:69:@21280.4]
  wire [10:0] _T_1446; // @[Mux.scala 31:69:@21281.4]
  wire [10:0] _T_1447; // @[Mux.scala 31:69:@21282.4]
  wire [10:0] _T_1448; // @[Mux.scala 31:69:@21283.4]
  wire [10:0] _T_1449; // @[Mux.scala 31:69:@21284.4]
  wire [10:0] _T_1450; // @[Mux.scala 31:69:@21285.4]
  wire [10:0] _T_1451; // @[Mux.scala 31:69:@21286.4]
  wire  _T_1458; // @[MemPrimitives.scala 110:210:@21294.4]
  wire  _T_1459; // @[MemPrimitives.scala 110:228:@21295.4]
  wire  _T_1464; // @[MemPrimitives.scala 110:210:@21298.4]
  wire  _T_1465; // @[MemPrimitives.scala 110:228:@21299.4]
  wire  _T_1470; // @[MemPrimitives.scala 110:210:@21302.4]
  wire  _T_1471; // @[MemPrimitives.scala 110:228:@21303.4]
  wire  _T_1476; // @[MemPrimitives.scala 110:210:@21306.4]
  wire  _T_1477; // @[MemPrimitives.scala 110:228:@21307.4]
  wire  _T_1482; // @[MemPrimitives.scala 110:210:@21310.4]
  wire  _T_1483; // @[MemPrimitives.scala 110:228:@21311.4]
  wire  _T_1488; // @[MemPrimitives.scala 110:210:@21314.4]
  wire  _T_1489; // @[MemPrimitives.scala 110:228:@21315.4]
  wire  _T_1494; // @[MemPrimitives.scala 110:210:@21318.4]
  wire  _T_1495; // @[MemPrimitives.scala 110:228:@21319.4]
  wire  _T_1500; // @[MemPrimitives.scala 110:210:@21322.4]
  wire  _T_1501; // @[MemPrimitives.scala 110:228:@21323.4]
  wire  _T_1506; // @[MemPrimitives.scala 110:210:@21326.4]
  wire  _T_1507; // @[MemPrimitives.scala 110:228:@21327.4]
  wire  _T_1509; // @[MemPrimitives.scala 126:35:@21341.4]
  wire  _T_1510; // @[MemPrimitives.scala 126:35:@21342.4]
  wire  _T_1511; // @[MemPrimitives.scala 126:35:@21343.4]
  wire  _T_1512; // @[MemPrimitives.scala 126:35:@21344.4]
  wire  _T_1513; // @[MemPrimitives.scala 126:35:@21345.4]
  wire  _T_1514; // @[MemPrimitives.scala 126:35:@21346.4]
  wire  _T_1515; // @[MemPrimitives.scala 126:35:@21347.4]
  wire  _T_1516; // @[MemPrimitives.scala 126:35:@21348.4]
  wire  _T_1517; // @[MemPrimitives.scala 126:35:@21349.4]
  wire [10:0] _T_1519; // @[Cat.scala 30:58:@21351.4]
  wire [10:0] _T_1521; // @[Cat.scala 30:58:@21353.4]
  wire [10:0] _T_1523; // @[Cat.scala 30:58:@21355.4]
  wire [10:0] _T_1525; // @[Cat.scala 30:58:@21357.4]
  wire [10:0] _T_1527; // @[Cat.scala 30:58:@21359.4]
  wire [10:0] _T_1529; // @[Cat.scala 30:58:@21361.4]
  wire [10:0] _T_1531; // @[Cat.scala 30:58:@21363.4]
  wire [10:0] _T_1533; // @[Cat.scala 30:58:@21365.4]
  wire [10:0] _T_1535; // @[Cat.scala 30:58:@21367.4]
  wire [10:0] _T_1536; // @[Mux.scala 31:69:@21368.4]
  wire [10:0] _T_1537; // @[Mux.scala 31:69:@21369.4]
  wire [10:0] _T_1538; // @[Mux.scala 31:69:@21370.4]
  wire [10:0] _T_1539; // @[Mux.scala 31:69:@21371.4]
  wire [10:0] _T_1540; // @[Mux.scala 31:69:@21372.4]
  wire [10:0] _T_1541; // @[Mux.scala 31:69:@21373.4]
  wire [10:0] _T_1542; // @[Mux.scala 31:69:@21374.4]
  wire [10:0] _T_1543; // @[Mux.scala 31:69:@21375.4]
  wire  _T_1550; // @[MemPrimitives.scala 110:210:@21383.4]
  wire  _T_1551; // @[MemPrimitives.scala 110:228:@21384.4]
  wire  _T_1556; // @[MemPrimitives.scala 110:210:@21387.4]
  wire  _T_1557; // @[MemPrimitives.scala 110:228:@21388.4]
  wire  _T_1562; // @[MemPrimitives.scala 110:210:@21391.4]
  wire  _T_1563; // @[MemPrimitives.scala 110:228:@21392.4]
  wire  _T_1568; // @[MemPrimitives.scala 110:210:@21395.4]
  wire  _T_1569; // @[MemPrimitives.scala 110:228:@21396.4]
  wire  _T_1574; // @[MemPrimitives.scala 110:210:@21399.4]
  wire  _T_1575; // @[MemPrimitives.scala 110:228:@21400.4]
  wire  _T_1580; // @[MemPrimitives.scala 110:210:@21403.4]
  wire  _T_1581; // @[MemPrimitives.scala 110:228:@21404.4]
  wire  _T_1586; // @[MemPrimitives.scala 110:210:@21407.4]
  wire  _T_1587; // @[MemPrimitives.scala 110:228:@21408.4]
  wire  _T_1592; // @[MemPrimitives.scala 110:210:@21411.4]
  wire  _T_1593; // @[MemPrimitives.scala 110:228:@21412.4]
  wire  _T_1598; // @[MemPrimitives.scala 110:210:@21415.4]
  wire  _T_1599; // @[MemPrimitives.scala 110:228:@21416.4]
  wire  _T_1601; // @[MemPrimitives.scala 126:35:@21430.4]
  wire  _T_1602; // @[MemPrimitives.scala 126:35:@21431.4]
  wire  _T_1603; // @[MemPrimitives.scala 126:35:@21432.4]
  wire  _T_1604; // @[MemPrimitives.scala 126:35:@21433.4]
  wire  _T_1605; // @[MemPrimitives.scala 126:35:@21434.4]
  wire  _T_1606; // @[MemPrimitives.scala 126:35:@21435.4]
  wire  _T_1607; // @[MemPrimitives.scala 126:35:@21436.4]
  wire  _T_1608; // @[MemPrimitives.scala 126:35:@21437.4]
  wire  _T_1609; // @[MemPrimitives.scala 126:35:@21438.4]
  wire [10:0] _T_1611; // @[Cat.scala 30:58:@21440.4]
  wire [10:0] _T_1613; // @[Cat.scala 30:58:@21442.4]
  wire [10:0] _T_1615; // @[Cat.scala 30:58:@21444.4]
  wire [10:0] _T_1617; // @[Cat.scala 30:58:@21446.4]
  wire [10:0] _T_1619; // @[Cat.scala 30:58:@21448.4]
  wire [10:0] _T_1621; // @[Cat.scala 30:58:@21450.4]
  wire [10:0] _T_1623; // @[Cat.scala 30:58:@21452.4]
  wire [10:0] _T_1625; // @[Cat.scala 30:58:@21454.4]
  wire [10:0] _T_1627; // @[Cat.scala 30:58:@21456.4]
  wire [10:0] _T_1628; // @[Mux.scala 31:69:@21457.4]
  wire [10:0] _T_1629; // @[Mux.scala 31:69:@21458.4]
  wire [10:0] _T_1630; // @[Mux.scala 31:69:@21459.4]
  wire [10:0] _T_1631; // @[Mux.scala 31:69:@21460.4]
  wire [10:0] _T_1632; // @[Mux.scala 31:69:@21461.4]
  wire [10:0] _T_1633; // @[Mux.scala 31:69:@21462.4]
  wire [10:0] _T_1634; // @[Mux.scala 31:69:@21463.4]
  wire [10:0] _T_1635; // @[Mux.scala 31:69:@21464.4]
  wire  _T_1642; // @[MemPrimitives.scala 110:210:@21472.4]
  wire  _T_1643; // @[MemPrimitives.scala 110:228:@21473.4]
  wire  _T_1648; // @[MemPrimitives.scala 110:210:@21476.4]
  wire  _T_1649; // @[MemPrimitives.scala 110:228:@21477.4]
  wire  _T_1654; // @[MemPrimitives.scala 110:210:@21480.4]
  wire  _T_1655; // @[MemPrimitives.scala 110:228:@21481.4]
  wire  _T_1660; // @[MemPrimitives.scala 110:210:@21484.4]
  wire  _T_1661; // @[MemPrimitives.scala 110:228:@21485.4]
  wire  _T_1666; // @[MemPrimitives.scala 110:210:@21488.4]
  wire  _T_1667; // @[MemPrimitives.scala 110:228:@21489.4]
  wire  _T_1672; // @[MemPrimitives.scala 110:210:@21492.4]
  wire  _T_1673; // @[MemPrimitives.scala 110:228:@21493.4]
  wire  _T_1678; // @[MemPrimitives.scala 110:210:@21496.4]
  wire  _T_1679; // @[MemPrimitives.scala 110:228:@21497.4]
  wire  _T_1684; // @[MemPrimitives.scala 110:210:@21500.4]
  wire  _T_1685; // @[MemPrimitives.scala 110:228:@21501.4]
  wire  _T_1690; // @[MemPrimitives.scala 110:210:@21504.4]
  wire  _T_1691; // @[MemPrimitives.scala 110:228:@21505.4]
  wire  _T_1693; // @[MemPrimitives.scala 126:35:@21519.4]
  wire  _T_1694; // @[MemPrimitives.scala 126:35:@21520.4]
  wire  _T_1695; // @[MemPrimitives.scala 126:35:@21521.4]
  wire  _T_1696; // @[MemPrimitives.scala 126:35:@21522.4]
  wire  _T_1697; // @[MemPrimitives.scala 126:35:@21523.4]
  wire  _T_1698; // @[MemPrimitives.scala 126:35:@21524.4]
  wire  _T_1699; // @[MemPrimitives.scala 126:35:@21525.4]
  wire  _T_1700; // @[MemPrimitives.scala 126:35:@21526.4]
  wire  _T_1701; // @[MemPrimitives.scala 126:35:@21527.4]
  wire [10:0] _T_1703; // @[Cat.scala 30:58:@21529.4]
  wire [10:0] _T_1705; // @[Cat.scala 30:58:@21531.4]
  wire [10:0] _T_1707; // @[Cat.scala 30:58:@21533.4]
  wire [10:0] _T_1709; // @[Cat.scala 30:58:@21535.4]
  wire [10:0] _T_1711; // @[Cat.scala 30:58:@21537.4]
  wire [10:0] _T_1713; // @[Cat.scala 30:58:@21539.4]
  wire [10:0] _T_1715; // @[Cat.scala 30:58:@21541.4]
  wire [10:0] _T_1717; // @[Cat.scala 30:58:@21543.4]
  wire [10:0] _T_1719; // @[Cat.scala 30:58:@21545.4]
  wire [10:0] _T_1720; // @[Mux.scala 31:69:@21546.4]
  wire [10:0] _T_1721; // @[Mux.scala 31:69:@21547.4]
  wire [10:0] _T_1722; // @[Mux.scala 31:69:@21548.4]
  wire [10:0] _T_1723; // @[Mux.scala 31:69:@21549.4]
  wire [10:0] _T_1724; // @[Mux.scala 31:69:@21550.4]
  wire [10:0] _T_1725; // @[Mux.scala 31:69:@21551.4]
  wire [10:0] _T_1726; // @[Mux.scala 31:69:@21552.4]
  wire [10:0] _T_1727; // @[Mux.scala 31:69:@21553.4]
  wire  _T_1732; // @[MemPrimitives.scala 110:210:@21560.4]
  wire  _T_1735; // @[MemPrimitives.scala 110:228:@21562.4]
  wire  _T_1738; // @[MemPrimitives.scala 110:210:@21564.4]
  wire  _T_1741; // @[MemPrimitives.scala 110:228:@21566.4]
  wire  _T_1744; // @[MemPrimitives.scala 110:210:@21568.4]
  wire  _T_1747; // @[MemPrimitives.scala 110:228:@21570.4]
  wire  _T_1750; // @[MemPrimitives.scala 110:210:@21572.4]
  wire  _T_1753; // @[MemPrimitives.scala 110:228:@21574.4]
  wire  _T_1756; // @[MemPrimitives.scala 110:210:@21576.4]
  wire  _T_1759; // @[MemPrimitives.scala 110:228:@21578.4]
  wire  _T_1762; // @[MemPrimitives.scala 110:210:@21580.4]
  wire  _T_1765; // @[MemPrimitives.scala 110:228:@21582.4]
  wire  _T_1768; // @[MemPrimitives.scala 110:210:@21584.4]
  wire  _T_1771; // @[MemPrimitives.scala 110:228:@21586.4]
  wire  _T_1774; // @[MemPrimitives.scala 110:210:@21588.4]
  wire  _T_1777; // @[MemPrimitives.scala 110:228:@21590.4]
  wire  _T_1780; // @[MemPrimitives.scala 110:210:@21592.4]
  wire  _T_1783; // @[MemPrimitives.scala 110:228:@21594.4]
  wire  _T_1785; // @[MemPrimitives.scala 126:35:@21608.4]
  wire  _T_1786; // @[MemPrimitives.scala 126:35:@21609.4]
  wire  _T_1787; // @[MemPrimitives.scala 126:35:@21610.4]
  wire  _T_1788; // @[MemPrimitives.scala 126:35:@21611.4]
  wire  _T_1789; // @[MemPrimitives.scala 126:35:@21612.4]
  wire  _T_1790; // @[MemPrimitives.scala 126:35:@21613.4]
  wire  _T_1791; // @[MemPrimitives.scala 126:35:@21614.4]
  wire  _T_1792; // @[MemPrimitives.scala 126:35:@21615.4]
  wire  _T_1793; // @[MemPrimitives.scala 126:35:@21616.4]
  wire [10:0] _T_1795; // @[Cat.scala 30:58:@21618.4]
  wire [10:0] _T_1797; // @[Cat.scala 30:58:@21620.4]
  wire [10:0] _T_1799; // @[Cat.scala 30:58:@21622.4]
  wire [10:0] _T_1801; // @[Cat.scala 30:58:@21624.4]
  wire [10:0] _T_1803; // @[Cat.scala 30:58:@21626.4]
  wire [10:0] _T_1805; // @[Cat.scala 30:58:@21628.4]
  wire [10:0] _T_1807; // @[Cat.scala 30:58:@21630.4]
  wire [10:0] _T_1809; // @[Cat.scala 30:58:@21632.4]
  wire [10:0] _T_1811; // @[Cat.scala 30:58:@21634.4]
  wire [10:0] _T_1812; // @[Mux.scala 31:69:@21635.4]
  wire [10:0] _T_1813; // @[Mux.scala 31:69:@21636.4]
  wire [10:0] _T_1814; // @[Mux.scala 31:69:@21637.4]
  wire [10:0] _T_1815; // @[Mux.scala 31:69:@21638.4]
  wire [10:0] _T_1816; // @[Mux.scala 31:69:@21639.4]
  wire [10:0] _T_1817; // @[Mux.scala 31:69:@21640.4]
  wire [10:0] _T_1818; // @[Mux.scala 31:69:@21641.4]
  wire [10:0] _T_1819; // @[Mux.scala 31:69:@21642.4]
  wire  _T_1824; // @[MemPrimitives.scala 110:210:@21649.4]
  wire  _T_1827; // @[MemPrimitives.scala 110:228:@21651.4]
  wire  _T_1830; // @[MemPrimitives.scala 110:210:@21653.4]
  wire  _T_1833; // @[MemPrimitives.scala 110:228:@21655.4]
  wire  _T_1836; // @[MemPrimitives.scala 110:210:@21657.4]
  wire  _T_1839; // @[MemPrimitives.scala 110:228:@21659.4]
  wire  _T_1842; // @[MemPrimitives.scala 110:210:@21661.4]
  wire  _T_1845; // @[MemPrimitives.scala 110:228:@21663.4]
  wire  _T_1848; // @[MemPrimitives.scala 110:210:@21665.4]
  wire  _T_1851; // @[MemPrimitives.scala 110:228:@21667.4]
  wire  _T_1854; // @[MemPrimitives.scala 110:210:@21669.4]
  wire  _T_1857; // @[MemPrimitives.scala 110:228:@21671.4]
  wire  _T_1860; // @[MemPrimitives.scala 110:210:@21673.4]
  wire  _T_1863; // @[MemPrimitives.scala 110:228:@21675.4]
  wire  _T_1866; // @[MemPrimitives.scala 110:210:@21677.4]
  wire  _T_1869; // @[MemPrimitives.scala 110:228:@21679.4]
  wire  _T_1872; // @[MemPrimitives.scala 110:210:@21681.4]
  wire  _T_1875; // @[MemPrimitives.scala 110:228:@21683.4]
  wire  _T_1877; // @[MemPrimitives.scala 126:35:@21697.4]
  wire  _T_1878; // @[MemPrimitives.scala 126:35:@21698.4]
  wire  _T_1879; // @[MemPrimitives.scala 126:35:@21699.4]
  wire  _T_1880; // @[MemPrimitives.scala 126:35:@21700.4]
  wire  _T_1881; // @[MemPrimitives.scala 126:35:@21701.4]
  wire  _T_1882; // @[MemPrimitives.scala 126:35:@21702.4]
  wire  _T_1883; // @[MemPrimitives.scala 126:35:@21703.4]
  wire  _T_1884; // @[MemPrimitives.scala 126:35:@21704.4]
  wire  _T_1885; // @[MemPrimitives.scala 126:35:@21705.4]
  wire [10:0] _T_1887; // @[Cat.scala 30:58:@21707.4]
  wire [10:0] _T_1889; // @[Cat.scala 30:58:@21709.4]
  wire [10:0] _T_1891; // @[Cat.scala 30:58:@21711.4]
  wire [10:0] _T_1893; // @[Cat.scala 30:58:@21713.4]
  wire [10:0] _T_1895; // @[Cat.scala 30:58:@21715.4]
  wire [10:0] _T_1897; // @[Cat.scala 30:58:@21717.4]
  wire [10:0] _T_1899; // @[Cat.scala 30:58:@21719.4]
  wire [10:0] _T_1901; // @[Cat.scala 30:58:@21721.4]
  wire [10:0] _T_1903; // @[Cat.scala 30:58:@21723.4]
  wire [10:0] _T_1904; // @[Mux.scala 31:69:@21724.4]
  wire [10:0] _T_1905; // @[Mux.scala 31:69:@21725.4]
  wire [10:0] _T_1906; // @[Mux.scala 31:69:@21726.4]
  wire [10:0] _T_1907; // @[Mux.scala 31:69:@21727.4]
  wire [10:0] _T_1908; // @[Mux.scala 31:69:@21728.4]
  wire [10:0] _T_1909; // @[Mux.scala 31:69:@21729.4]
  wire [10:0] _T_1910; // @[Mux.scala 31:69:@21730.4]
  wire [10:0] _T_1911; // @[Mux.scala 31:69:@21731.4]
  wire  _T_1919; // @[MemPrimitives.scala 110:228:@21740.4]
  wire  _T_1925; // @[MemPrimitives.scala 110:228:@21744.4]
  wire  _T_1931; // @[MemPrimitives.scala 110:228:@21748.4]
  wire  _T_1937; // @[MemPrimitives.scala 110:228:@21752.4]
  wire  _T_1943; // @[MemPrimitives.scala 110:228:@21756.4]
  wire  _T_1949; // @[MemPrimitives.scala 110:228:@21760.4]
  wire  _T_1955; // @[MemPrimitives.scala 110:228:@21764.4]
  wire  _T_1961; // @[MemPrimitives.scala 110:228:@21768.4]
  wire  _T_1967; // @[MemPrimitives.scala 110:228:@21772.4]
  wire  _T_1969; // @[MemPrimitives.scala 126:35:@21786.4]
  wire  _T_1970; // @[MemPrimitives.scala 126:35:@21787.4]
  wire  _T_1971; // @[MemPrimitives.scala 126:35:@21788.4]
  wire  _T_1972; // @[MemPrimitives.scala 126:35:@21789.4]
  wire  _T_1973; // @[MemPrimitives.scala 126:35:@21790.4]
  wire  _T_1974; // @[MemPrimitives.scala 126:35:@21791.4]
  wire  _T_1975; // @[MemPrimitives.scala 126:35:@21792.4]
  wire  _T_1976; // @[MemPrimitives.scala 126:35:@21793.4]
  wire  _T_1977; // @[MemPrimitives.scala 126:35:@21794.4]
  wire [10:0] _T_1979; // @[Cat.scala 30:58:@21796.4]
  wire [10:0] _T_1981; // @[Cat.scala 30:58:@21798.4]
  wire [10:0] _T_1983; // @[Cat.scala 30:58:@21800.4]
  wire [10:0] _T_1985; // @[Cat.scala 30:58:@21802.4]
  wire [10:0] _T_1987; // @[Cat.scala 30:58:@21804.4]
  wire [10:0] _T_1989; // @[Cat.scala 30:58:@21806.4]
  wire [10:0] _T_1991; // @[Cat.scala 30:58:@21808.4]
  wire [10:0] _T_1993; // @[Cat.scala 30:58:@21810.4]
  wire [10:0] _T_1995; // @[Cat.scala 30:58:@21812.4]
  wire [10:0] _T_1996; // @[Mux.scala 31:69:@21813.4]
  wire [10:0] _T_1997; // @[Mux.scala 31:69:@21814.4]
  wire [10:0] _T_1998; // @[Mux.scala 31:69:@21815.4]
  wire [10:0] _T_1999; // @[Mux.scala 31:69:@21816.4]
  wire [10:0] _T_2000; // @[Mux.scala 31:69:@21817.4]
  wire [10:0] _T_2001; // @[Mux.scala 31:69:@21818.4]
  wire [10:0] _T_2002; // @[Mux.scala 31:69:@21819.4]
  wire [10:0] _T_2003; // @[Mux.scala 31:69:@21820.4]
  wire  _T_2011; // @[MemPrimitives.scala 110:228:@21829.4]
  wire  _T_2017; // @[MemPrimitives.scala 110:228:@21833.4]
  wire  _T_2023; // @[MemPrimitives.scala 110:228:@21837.4]
  wire  _T_2029; // @[MemPrimitives.scala 110:228:@21841.4]
  wire  _T_2035; // @[MemPrimitives.scala 110:228:@21845.4]
  wire  _T_2041; // @[MemPrimitives.scala 110:228:@21849.4]
  wire  _T_2047; // @[MemPrimitives.scala 110:228:@21853.4]
  wire  _T_2053; // @[MemPrimitives.scala 110:228:@21857.4]
  wire  _T_2059; // @[MemPrimitives.scala 110:228:@21861.4]
  wire  _T_2061; // @[MemPrimitives.scala 126:35:@21875.4]
  wire  _T_2062; // @[MemPrimitives.scala 126:35:@21876.4]
  wire  _T_2063; // @[MemPrimitives.scala 126:35:@21877.4]
  wire  _T_2064; // @[MemPrimitives.scala 126:35:@21878.4]
  wire  _T_2065; // @[MemPrimitives.scala 126:35:@21879.4]
  wire  _T_2066; // @[MemPrimitives.scala 126:35:@21880.4]
  wire  _T_2067; // @[MemPrimitives.scala 126:35:@21881.4]
  wire  _T_2068; // @[MemPrimitives.scala 126:35:@21882.4]
  wire  _T_2069; // @[MemPrimitives.scala 126:35:@21883.4]
  wire [10:0] _T_2071; // @[Cat.scala 30:58:@21885.4]
  wire [10:0] _T_2073; // @[Cat.scala 30:58:@21887.4]
  wire [10:0] _T_2075; // @[Cat.scala 30:58:@21889.4]
  wire [10:0] _T_2077; // @[Cat.scala 30:58:@21891.4]
  wire [10:0] _T_2079; // @[Cat.scala 30:58:@21893.4]
  wire [10:0] _T_2081; // @[Cat.scala 30:58:@21895.4]
  wire [10:0] _T_2083; // @[Cat.scala 30:58:@21897.4]
  wire [10:0] _T_2085; // @[Cat.scala 30:58:@21899.4]
  wire [10:0] _T_2087; // @[Cat.scala 30:58:@21901.4]
  wire [10:0] _T_2088; // @[Mux.scala 31:69:@21902.4]
  wire [10:0] _T_2089; // @[Mux.scala 31:69:@21903.4]
  wire [10:0] _T_2090; // @[Mux.scala 31:69:@21904.4]
  wire [10:0] _T_2091; // @[Mux.scala 31:69:@21905.4]
  wire [10:0] _T_2092; // @[Mux.scala 31:69:@21906.4]
  wire [10:0] _T_2093; // @[Mux.scala 31:69:@21907.4]
  wire [10:0] _T_2094; // @[Mux.scala 31:69:@21908.4]
  wire [10:0] _T_2095; // @[Mux.scala 31:69:@21909.4]
  wire  _T_2103; // @[MemPrimitives.scala 110:228:@21918.4]
  wire  _T_2109; // @[MemPrimitives.scala 110:228:@21922.4]
  wire  _T_2115; // @[MemPrimitives.scala 110:228:@21926.4]
  wire  _T_2121; // @[MemPrimitives.scala 110:228:@21930.4]
  wire  _T_2127; // @[MemPrimitives.scala 110:228:@21934.4]
  wire  _T_2133; // @[MemPrimitives.scala 110:228:@21938.4]
  wire  _T_2139; // @[MemPrimitives.scala 110:228:@21942.4]
  wire  _T_2145; // @[MemPrimitives.scala 110:228:@21946.4]
  wire  _T_2151; // @[MemPrimitives.scala 110:228:@21950.4]
  wire  _T_2153; // @[MemPrimitives.scala 126:35:@21964.4]
  wire  _T_2154; // @[MemPrimitives.scala 126:35:@21965.4]
  wire  _T_2155; // @[MemPrimitives.scala 126:35:@21966.4]
  wire  _T_2156; // @[MemPrimitives.scala 126:35:@21967.4]
  wire  _T_2157; // @[MemPrimitives.scala 126:35:@21968.4]
  wire  _T_2158; // @[MemPrimitives.scala 126:35:@21969.4]
  wire  _T_2159; // @[MemPrimitives.scala 126:35:@21970.4]
  wire  _T_2160; // @[MemPrimitives.scala 126:35:@21971.4]
  wire  _T_2161; // @[MemPrimitives.scala 126:35:@21972.4]
  wire [10:0] _T_2163; // @[Cat.scala 30:58:@21974.4]
  wire [10:0] _T_2165; // @[Cat.scala 30:58:@21976.4]
  wire [10:0] _T_2167; // @[Cat.scala 30:58:@21978.4]
  wire [10:0] _T_2169; // @[Cat.scala 30:58:@21980.4]
  wire [10:0] _T_2171; // @[Cat.scala 30:58:@21982.4]
  wire [10:0] _T_2173; // @[Cat.scala 30:58:@21984.4]
  wire [10:0] _T_2175; // @[Cat.scala 30:58:@21986.4]
  wire [10:0] _T_2177; // @[Cat.scala 30:58:@21988.4]
  wire [10:0] _T_2179; // @[Cat.scala 30:58:@21990.4]
  wire [10:0] _T_2180; // @[Mux.scala 31:69:@21991.4]
  wire [10:0] _T_2181; // @[Mux.scala 31:69:@21992.4]
  wire [10:0] _T_2182; // @[Mux.scala 31:69:@21993.4]
  wire [10:0] _T_2183; // @[Mux.scala 31:69:@21994.4]
  wire [10:0] _T_2184; // @[Mux.scala 31:69:@21995.4]
  wire [10:0] _T_2185; // @[Mux.scala 31:69:@21996.4]
  wire [10:0] _T_2186; // @[Mux.scala 31:69:@21997.4]
  wire [10:0] _T_2187; // @[Mux.scala 31:69:@21998.4]
  wire  _T_2195; // @[MemPrimitives.scala 110:228:@22007.4]
  wire  _T_2201; // @[MemPrimitives.scala 110:228:@22011.4]
  wire  _T_2207; // @[MemPrimitives.scala 110:228:@22015.4]
  wire  _T_2213; // @[MemPrimitives.scala 110:228:@22019.4]
  wire  _T_2219; // @[MemPrimitives.scala 110:228:@22023.4]
  wire  _T_2225; // @[MemPrimitives.scala 110:228:@22027.4]
  wire  _T_2231; // @[MemPrimitives.scala 110:228:@22031.4]
  wire  _T_2237; // @[MemPrimitives.scala 110:228:@22035.4]
  wire  _T_2243; // @[MemPrimitives.scala 110:228:@22039.4]
  wire  _T_2245; // @[MemPrimitives.scala 126:35:@22053.4]
  wire  _T_2246; // @[MemPrimitives.scala 126:35:@22054.4]
  wire  _T_2247; // @[MemPrimitives.scala 126:35:@22055.4]
  wire  _T_2248; // @[MemPrimitives.scala 126:35:@22056.4]
  wire  _T_2249; // @[MemPrimitives.scala 126:35:@22057.4]
  wire  _T_2250; // @[MemPrimitives.scala 126:35:@22058.4]
  wire  _T_2251; // @[MemPrimitives.scala 126:35:@22059.4]
  wire  _T_2252; // @[MemPrimitives.scala 126:35:@22060.4]
  wire  _T_2253; // @[MemPrimitives.scala 126:35:@22061.4]
  wire [10:0] _T_2255; // @[Cat.scala 30:58:@22063.4]
  wire [10:0] _T_2257; // @[Cat.scala 30:58:@22065.4]
  wire [10:0] _T_2259; // @[Cat.scala 30:58:@22067.4]
  wire [10:0] _T_2261; // @[Cat.scala 30:58:@22069.4]
  wire [10:0] _T_2263; // @[Cat.scala 30:58:@22071.4]
  wire [10:0] _T_2265; // @[Cat.scala 30:58:@22073.4]
  wire [10:0] _T_2267; // @[Cat.scala 30:58:@22075.4]
  wire [10:0] _T_2269; // @[Cat.scala 30:58:@22077.4]
  wire [10:0] _T_2271; // @[Cat.scala 30:58:@22079.4]
  wire [10:0] _T_2272; // @[Mux.scala 31:69:@22080.4]
  wire [10:0] _T_2273; // @[Mux.scala 31:69:@22081.4]
  wire [10:0] _T_2274; // @[Mux.scala 31:69:@22082.4]
  wire [10:0] _T_2275; // @[Mux.scala 31:69:@22083.4]
  wire [10:0] _T_2276; // @[Mux.scala 31:69:@22084.4]
  wire [10:0] _T_2277; // @[Mux.scala 31:69:@22085.4]
  wire [10:0] _T_2278; // @[Mux.scala 31:69:@22086.4]
  wire [10:0] _T_2279; // @[Mux.scala 31:69:@22087.4]
  wire  _T_2284; // @[MemPrimitives.scala 110:210:@22094.4]
  wire  _T_2287; // @[MemPrimitives.scala 110:228:@22096.4]
  wire  _T_2290; // @[MemPrimitives.scala 110:210:@22098.4]
  wire  _T_2293; // @[MemPrimitives.scala 110:228:@22100.4]
  wire  _T_2296; // @[MemPrimitives.scala 110:210:@22102.4]
  wire  _T_2299; // @[MemPrimitives.scala 110:228:@22104.4]
  wire  _T_2302; // @[MemPrimitives.scala 110:210:@22106.4]
  wire  _T_2305; // @[MemPrimitives.scala 110:228:@22108.4]
  wire  _T_2308; // @[MemPrimitives.scala 110:210:@22110.4]
  wire  _T_2311; // @[MemPrimitives.scala 110:228:@22112.4]
  wire  _T_2314; // @[MemPrimitives.scala 110:210:@22114.4]
  wire  _T_2317; // @[MemPrimitives.scala 110:228:@22116.4]
  wire  _T_2320; // @[MemPrimitives.scala 110:210:@22118.4]
  wire  _T_2323; // @[MemPrimitives.scala 110:228:@22120.4]
  wire  _T_2326; // @[MemPrimitives.scala 110:210:@22122.4]
  wire  _T_2329; // @[MemPrimitives.scala 110:228:@22124.4]
  wire  _T_2332; // @[MemPrimitives.scala 110:210:@22126.4]
  wire  _T_2335; // @[MemPrimitives.scala 110:228:@22128.4]
  wire  _T_2337; // @[MemPrimitives.scala 126:35:@22142.4]
  wire  _T_2338; // @[MemPrimitives.scala 126:35:@22143.4]
  wire  _T_2339; // @[MemPrimitives.scala 126:35:@22144.4]
  wire  _T_2340; // @[MemPrimitives.scala 126:35:@22145.4]
  wire  _T_2341; // @[MemPrimitives.scala 126:35:@22146.4]
  wire  _T_2342; // @[MemPrimitives.scala 126:35:@22147.4]
  wire  _T_2343; // @[MemPrimitives.scala 126:35:@22148.4]
  wire  _T_2344; // @[MemPrimitives.scala 126:35:@22149.4]
  wire  _T_2345; // @[MemPrimitives.scala 126:35:@22150.4]
  wire [10:0] _T_2347; // @[Cat.scala 30:58:@22152.4]
  wire [10:0] _T_2349; // @[Cat.scala 30:58:@22154.4]
  wire [10:0] _T_2351; // @[Cat.scala 30:58:@22156.4]
  wire [10:0] _T_2353; // @[Cat.scala 30:58:@22158.4]
  wire [10:0] _T_2355; // @[Cat.scala 30:58:@22160.4]
  wire [10:0] _T_2357; // @[Cat.scala 30:58:@22162.4]
  wire [10:0] _T_2359; // @[Cat.scala 30:58:@22164.4]
  wire [10:0] _T_2361; // @[Cat.scala 30:58:@22166.4]
  wire [10:0] _T_2363; // @[Cat.scala 30:58:@22168.4]
  wire [10:0] _T_2364; // @[Mux.scala 31:69:@22169.4]
  wire [10:0] _T_2365; // @[Mux.scala 31:69:@22170.4]
  wire [10:0] _T_2366; // @[Mux.scala 31:69:@22171.4]
  wire [10:0] _T_2367; // @[Mux.scala 31:69:@22172.4]
  wire [10:0] _T_2368; // @[Mux.scala 31:69:@22173.4]
  wire [10:0] _T_2369; // @[Mux.scala 31:69:@22174.4]
  wire [10:0] _T_2370; // @[Mux.scala 31:69:@22175.4]
  wire [10:0] _T_2371; // @[Mux.scala 31:69:@22176.4]
  wire  _T_2376; // @[MemPrimitives.scala 110:210:@22183.4]
  wire  _T_2379; // @[MemPrimitives.scala 110:228:@22185.4]
  wire  _T_2382; // @[MemPrimitives.scala 110:210:@22187.4]
  wire  _T_2385; // @[MemPrimitives.scala 110:228:@22189.4]
  wire  _T_2388; // @[MemPrimitives.scala 110:210:@22191.4]
  wire  _T_2391; // @[MemPrimitives.scala 110:228:@22193.4]
  wire  _T_2394; // @[MemPrimitives.scala 110:210:@22195.4]
  wire  _T_2397; // @[MemPrimitives.scala 110:228:@22197.4]
  wire  _T_2400; // @[MemPrimitives.scala 110:210:@22199.4]
  wire  _T_2403; // @[MemPrimitives.scala 110:228:@22201.4]
  wire  _T_2406; // @[MemPrimitives.scala 110:210:@22203.4]
  wire  _T_2409; // @[MemPrimitives.scala 110:228:@22205.4]
  wire  _T_2412; // @[MemPrimitives.scala 110:210:@22207.4]
  wire  _T_2415; // @[MemPrimitives.scala 110:228:@22209.4]
  wire  _T_2418; // @[MemPrimitives.scala 110:210:@22211.4]
  wire  _T_2421; // @[MemPrimitives.scala 110:228:@22213.4]
  wire  _T_2424; // @[MemPrimitives.scala 110:210:@22215.4]
  wire  _T_2427; // @[MemPrimitives.scala 110:228:@22217.4]
  wire  _T_2429; // @[MemPrimitives.scala 126:35:@22231.4]
  wire  _T_2430; // @[MemPrimitives.scala 126:35:@22232.4]
  wire  _T_2431; // @[MemPrimitives.scala 126:35:@22233.4]
  wire  _T_2432; // @[MemPrimitives.scala 126:35:@22234.4]
  wire  _T_2433; // @[MemPrimitives.scala 126:35:@22235.4]
  wire  _T_2434; // @[MemPrimitives.scala 126:35:@22236.4]
  wire  _T_2435; // @[MemPrimitives.scala 126:35:@22237.4]
  wire  _T_2436; // @[MemPrimitives.scala 126:35:@22238.4]
  wire  _T_2437; // @[MemPrimitives.scala 126:35:@22239.4]
  wire [10:0] _T_2439; // @[Cat.scala 30:58:@22241.4]
  wire [10:0] _T_2441; // @[Cat.scala 30:58:@22243.4]
  wire [10:0] _T_2443; // @[Cat.scala 30:58:@22245.4]
  wire [10:0] _T_2445; // @[Cat.scala 30:58:@22247.4]
  wire [10:0] _T_2447; // @[Cat.scala 30:58:@22249.4]
  wire [10:0] _T_2449; // @[Cat.scala 30:58:@22251.4]
  wire [10:0] _T_2451; // @[Cat.scala 30:58:@22253.4]
  wire [10:0] _T_2453; // @[Cat.scala 30:58:@22255.4]
  wire [10:0] _T_2455; // @[Cat.scala 30:58:@22257.4]
  wire [10:0] _T_2456; // @[Mux.scala 31:69:@22258.4]
  wire [10:0] _T_2457; // @[Mux.scala 31:69:@22259.4]
  wire [10:0] _T_2458; // @[Mux.scala 31:69:@22260.4]
  wire [10:0] _T_2459; // @[Mux.scala 31:69:@22261.4]
  wire [10:0] _T_2460; // @[Mux.scala 31:69:@22262.4]
  wire [10:0] _T_2461; // @[Mux.scala 31:69:@22263.4]
  wire [10:0] _T_2462; // @[Mux.scala 31:69:@22264.4]
  wire [10:0] _T_2463; // @[Mux.scala 31:69:@22265.4]
  wire  _T_2471; // @[MemPrimitives.scala 110:228:@22274.4]
  wire  _T_2477; // @[MemPrimitives.scala 110:228:@22278.4]
  wire  _T_2483; // @[MemPrimitives.scala 110:228:@22282.4]
  wire  _T_2489; // @[MemPrimitives.scala 110:228:@22286.4]
  wire  _T_2495; // @[MemPrimitives.scala 110:228:@22290.4]
  wire  _T_2501; // @[MemPrimitives.scala 110:228:@22294.4]
  wire  _T_2507; // @[MemPrimitives.scala 110:228:@22298.4]
  wire  _T_2513; // @[MemPrimitives.scala 110:228:@22302.4]
  wire  _T_2519; // @[MemPrimitives.scala 110:228:@22306.4]
  wire  _T_2521; // @[MemPrimitives.scala 126:35:@22320.4]
  wire  _T_2522; // @[MemPrimitives.scala 126:35:@22321.4]
  wire  _T_2523; // @[MemPrimitives.scala 126:35:@22322.4]
  wire  _T_2524; // @[MemPrimitives.scala 126:35:@22323.4]
  wire  _T_2525; // @[MemPrimitives.scala 126:35:@22324.4]
  wire  _T_2526; // @[MemPrimitives.scala 126:35:@22325.4]
  wire  _T_2527; // @[MemPrimitives.scala 126:35:@22326.4]
  wire  _T_2528; // @[MemPrimitives.scala 126:35:@22327.4]
  wire  _T_2529; // @[MemPrimitives.scala 126:35:@22328.4]
  wire [10:0] _T_2531; // @[Cat.scala 30:58:@22330.4]
  wire [10:0] _T_2533; // @[Cat.scala 30:58:@22332.4]
  wire [10:0] _T_2535; // @[Cat.scala 30:58:@22334.4]
  wire [10:0] _T_2537; // @[Cat.scala 30:58:@22336.4]
  wire [10:0] _T_2539; // @[Cat.scala 30:58:@22338.4]
  wire [10:0] _T_2541; // @[Cat.scala 30:58:@22340.4]
  wire [10:0] _T_2543; // @[Cat.scala 30:58:@22342.4]
  wire [10:0] _T_2545; // @[Cat.scala 30:58:@22344.4]
  wire [10:0] _T_2547; // @[Cat.scala 30:58:@22346.4]
  wire [10:0] _T_2548; // @[Mux.scala 31:69:@22347.4]
  wire [10:0] _T_2549; // @[Mux.scala 31:69:@22348.4]
  wire [10:0] _T_2550; // @[Mux.scala 31:69:@22349.4]
  wire [10:0] _T_2551; // @[Mux.scala 31:69:@22350.4]
  wire [10:0] _T_2552; // @[Mux.scala 31:69:@22351.4]
  wire [10:0] _T_2553; // @[Mux.scala 31:69:@22352.4]
  wire [10:0] _T_2554; // @[Mux.scala 31:69:@22353.4]
  wire [10:0] _T_2555; // @[Mux.scala 31:69:@22354.4]
  wire  _T_2563; // @[MemPrimitives.scala 110:228:@22363.4]
  wire  _T_2569; // @[MemPrimitives.scala 110:228:@22367.4]
  wire  _T_2575; // @[MemPrimitives.scala 110:228:@22371.4]
  wire  _T_2581; // @[MemPrimitives.scala 110:228:@22375.4]
  wire  _T_2587; // @[MemPrimitives.scala 110:228:@22379.4]
  wire  _T_2593; // @[MemPrimitives.scala 110:228:@22383.4]
  wire  _T_2599; // @[MemPrimitives.scala 110:228:@22387.4]
  wire  _T_2605; // @[MemPrimitives.scala 110:228:@22391.4]
  wire  _T_2611; // @[MemPrimitives.scala 110:228:@22395.4]
  wire  _T_2613; // @[MemPrimitives.scala 126:35:@22409.4]
  wire  _T_2614; // @[MemPrimitives.scala 126:35:@22410.4]
  wire  _T_2615; // @[MemPrimitives.scala 126:35:@22411.4]
  wire  _T_2616; // @[MemPrimitives.scala 126:35:@22412.4]
  wire  _T_2617; // @[MemPrimitives.scala 126:35:@22413.4]
  wire  _T_2618; // @[MemPrimitives.scala 126:35:@22414.4]
  wire  _T_2619; // @[MemPrimitives.scala 126:35:@22415.4]
  wire  _T_2620; // @[MemPrimitives.scala 126:35:@22416.4]
  wire  _T_2621; // @[MemPrimitives.scala 126:35:@22417.4]
  wire [10:0] _T_2623; // @[Cat.scala 30:58:@22419.4]
  wire [10:0] _T_2625; // @[Cat.scala 30:58:@22421.4]
  wire [10:0] _T_2627; // @[Cat.scala 30:58:@22423.4]
  wire [10:0] _T_2629; // @[Cat.scala 30:58:@22425.4]
  wire [10:0] _T_2631; // @[Cat.scala 30:58:@22427.4]
  wire [10:0] _T_2633; // @[Cat.scala 30:58:@22429.4]
  wire [10:0] _T_2635; // @[Cat.scala 30:58:@22431.4]
  wire [10:0] _T_2637; // @[Cat.scala 30:58:@22433.4]
  wire [10:0] _T_2639; // @[Cat.scala 30:58:@22435.4]
  wire [10:0] _T_2640; // @[Mux.scala 31:69:@22436.4]
  wire [10:0] _T_2641; // @[Mux.scala 31:69:@22437.4]
  wire [10:0] _T_2642; // @[Mux.scala 31:69:@22438.4]
  wire [10:0] _T_2643; // @[Mux.scala 31:69:@22439.4]
  wire [10:0] _T_2644; // @[Mux.scala 31:69:@22440.4]
  wire [10:0] _T_2645; // @[Mux.scala 31:69:@22441.4]
  wire [10:0] _T_2646; // @[Mux.scala 31:69:@22442.4]
  wire [10:0] _T_2647; // @[Mux.scala 31:69:@22443.4]
  wire  _T_2655; // @[MemPrimitives.scala 110:228:@22452.4]
  wire  _T_2661; // @[MemPrimitives.scala 110:228:@22456.4]
  wire  _T_2667; // @[MemPrimitives.scala 110:228:@22460.4]
  wire  _T_2673; // @[MemPrimitives.scala 110:228:@22464.4]
  wire  _T_2679; // @[MemPrimitives.scala 110:228:@22468.4]
  wire  _T_2685; // @[MemPrimitives.scala 110:228:@22472.4]
  wire  _T_2691; // @[MemPrimitives.scala 110:228:@22476.4]
  wire  _T_2697; // @[MemPrimitives.scala 110:228:@22480.4]
  wire  _T_2703; // @[MemPrimitives.scala 110:228:@22484.4]
  wire  _T_2705; // @[MemPrimitives.scala 126:35:@22498.4]
  wire  _T_2706; // @[MemPrimitives.scala 126:35:@22499.4]
  wire  _T_2707; // @[MemPrimitives.scala 126:35:@22500.4]
  wire  _T_2708; // @[MemPrimitives.scala 126:35:@22501.4]
  wire  _T_2709; // @[MemPrimitives.scala 126:35:@22502.4]
  wire  _T_2710; // @[MemPrimitives.scala 126:35:@22503.4]
  wire  _T_2711; // @[MemPrimitives.scala 126:35:@22504.4]
  wire  _T_2712; // @[MemPrimitives.scala 126:35:@22505.4]
  wire  _T_2713; // @[MemPrimitives.scala 126:35:@22506.4]
  wire [10:0] _T_2715; // @[Cat.scala 30:58:@22508.4]
  wire [10:0] _T_2717; // @[Cat.scala 30:58:@22510.4]
  wire [10:0] _T_2719; // @[Cat.scala 30:58:@22512.4]
  wire [10:0] _T_2721; // @[Cat.scala 30:58:@22514.4]
  wire [10:0] _T_2723; // @[Cat.scala 30:58:@22516.4]
  wire [10:0] _T_2725; // @[Cat.scala 30:58:@22518.4]
  wire [10:0] _T_2727; // @[Cat.scala 30:58:@22520.4]
  wire [10:0] _T_2729; // @[Cat.scala 30:58:@22522.4]
  wire [10:0] _T_2731; // @[Cat.scala 30:58:@22524.4]
  wire [10:0] _T_2732; // @[Mux.scala 31:69:@22525.4]
  wire [10:0] _T_2733; // @[Mux.scala 31:69:@22526.4]
  wire [10:0] _T_2734; // @[Mux.scala 31:69:@22527.4]
  wire [10:0] _T_2735; // @[Mux.scala 31:69:@22528.4]
  wire [10:0] _T_2736; // @[Mux.scala 31:69:@22529.4]
  wire [10:0] _T_2737; // @[Mux.scala 31:69:@22530.4]
  wire [10:0] _T_2738; // @[Mux.scala 31:69:@22531.4]
  wire [10:0] _T_2739; // @[Mux.scala 31:69:@22532.4]
  wire  _T_2747; // @[MemPrimitives.scala 110:228:@22541.4]
  wire  _T_2753; // @[MemPrimitives.scala 110:228:@22545.4]
  wire  _T_2759; // @[MemPrimitives.scala 110:228:@22549.4]
  wire  _T_2765; // @[MemPrimitives.scala 110:228:@22553.4]
  wire  _T_2771; // @[MemPrimitives.scala 110:228:@22557.4]
  wire  _T_2777; // @[MemPrimitives.scala 110:228:@22561.4]
  wire  _T_2783; // @[MemPrimitives.scala 110:228:@22565.4]
  wire  _T_2789; // @[MemPrimitives.scala 110:228:@22569.4]
  wire  _T_2795; // @[MemPrimitives.scala 110:228:@22573.4]
  wire  _T_2797; // @[MemPrimitives.scala 126:35:@22587.4]
  wire  _T_2798; // @[MemPrimitives.scala 126:35:@22588.4]
  wire  _T_2799; // @[MemPrimitives.scala 126:35:@22589.4]
  wire  _T_2800; // @[MemPrimitives.scala 126:35:@22590.4]
  wire  _T_2801; // @[MemPrimitives.scala 126:35:@22591.4]
  wire  _T_2802; // @[MemPrimitives.scala 126:35:@22592.4]
  wire  _T_2803; // @[MemPrimitives.scala 126:35:@22593.4]
  wire  _T_2804; // @[MemPrimitives.scala 126:35:@22594.4]
  wire  _T_2805; // @[MemPrimitives.scala 126:35:@22595.4]
  wire [10:0] _T_2807; // @[Cat.scala 30:58:@22597.4]
  wire [10:0] _T_2809; // @[Cat.scala 30:58:@22599.4]
  wire [10:0] _T_2811; // @[Cat.scala 30:58:@22601.4]
  wire [10:0] _T_2813; // @[Cat.scala 30:58:@22603.4]
  wire [10:0] _T_2815; // @[Cat.scala 30:58:@22605.4]
  wire [10:0] _T_2817; // @[Cat.scala 30:58:@22607.4]
  wire [10:0] _T_2819; // @[Cat.scala 30:58:@22609.4]
  wire [10:0] _T_2821; // @[Cat.scala 30:58:@22611.4]
  wire [10:0] _T_2823; // @[Cat.scala 30:58:@22613.4]
  wire [10:0] _T_2824; // @[Mux.scala 31:69:@22614.4]
  wire [10:0] _T_2825; // @[Mux.scala 31:69:@22615.4]
  wire [10:0] _T_2826; // @[Mux.scala 31:69:@22616.4]
  wire [10:0] _T_2827; // @[Mux.scala 31:69:@22617.4]
  wire [10:0] _T_2828; // @[Mux.scala 31:69:@22618.4]
  wire [10:0] _T_2829; // @[Mux.scala 31:69:@22619.4]
  wire [10:0] _T_2830; // @[Mux.scala 31:69:@22620.4]
  wire [10:0] _T_2831; // @[Mux.scala 31:69:@22621.4]
  wire  _T_2836; // @[MemPrimitives.scala 110:210:@22628.4]
  wire  _T_2839; // @[MemPrimitives.scala 110:228:@22630.4]
  wire  _T_2842; // @[MemPrimitives.scala 110:210:@22632.4]
  wire  _T_2845; // @[MemPrimitives.scala 110:228:@22634.4]
  wire  _T_2848; // @[MemPrimitives.scala 110:210:@22636.4]
  wire  _T_2851; // @[MemPrimitives.scala 110:228:@22638.4]
  wire  _T_2854; // @[MemPrimitives.scala 110:210:@22640.4]
  wire  _T_2857; // @[MemPrimitives.scala 110:228:@22642.4]
  wire  _T_2860; // @[MemPrimitives.scala 110:210:@22644.4]
  wire  _T_2863; // @[MemPrimitives.scala 110:228:@22646.4]
  wire  _T_2866; // @[MemPrimitives.scala 110:210:@22648.4]
  wire  _T_2869; // @[MemPrimitives.scala 110:228:@22650.4]
  wire  _T_2872; // @[MemPrimitives.scala 110:210:@22652.4]
  wire  _T_2875; // @[MemPrimitives.scala 110:228:@22654.4]
  wire  _T_2878; // @[MemPrimitives.scala 110:210:@22656.4]
  wire  _T_2881; // @[MemPrimitives.scala 110:228:@22658.4]
  wire  _T_2884; // @[MemPrimitives.scala 110:210:@22660.4]
  wire  _T_2887; // @[MemPrimitives.scala 110:228:@22662.4]
  wire  _T_2889; // @[MemPrimitives.scala 126:35:@22676.4]
  wire  _T_2890; // @[MemPrimitives.scala 126:35:@22677.4]
  wire  _T_2891; // @[MemPrimitives.scala 126:35:@22678.4]
  wire  _T_2892; // @[MemPrimitives.scala 126:35:@22679.4]
  wire  _T_2893; // @[MemPrimitives.scala 126:35:@22680.4]
  wire  _T_2894; // @[MemPrimitives.scala 126:35:@22681.4]
  wire  _T_2895; // @[MemPrimitives.scala 126:35:@22682.4]
  wire  _T_2896; // @[MemPrimitives.scala 126:35:@22683.4]
  wire  _T_2897; // @[MemPrimitives.scala 126:35:@22684.4]
  wire [10:0] _T_2899; // @[Cat.scala 30:58:@22686.4]
  wire [10:0] _T_2901; // @[Cat.scala 30:58:@22688.4]
  wire [10:0] _T_2903; // @[Cat.scala 30:58:@22690.4]
  wire [10:0] _T_2905; // @[Cat.scala 30:58:@22692.4]
  wire [10:0] _T_2907; // @[Cat.scala 30:58:@22694.4]
  wire [10:0] _T_2909; // @[Cat.scala 30:58:@22696.4]
  wire [10:0] _T_2911; // @[Cat.scala 30:58:@22698.4]
  wire [10:0] _T_2913; // @[Cat.scala 30:58:@22700.4]
  wire [10:0] _T_2915; // @[Cat.scala 30:58:@22702.4]
  wire [10:0] _T_2916; // @[Mux.scala 31:69:@22703.4]
  wire [10:0] _T_2917; // @[Mux.scala 31:69:@22704.4]
  wire [10:0] _T_2918; // @[Mux.scala 31:69:@22705.4]
  wire [10:0] _T_2919; // @[Mux.scala 31:69:@22706.4]
  wire [10:0] _T_2920; // @[Mux.scala 31:69:@22707.4]
  wire [10:0] _T_2921; // @[Mux.scala 31:69:@22708.4]
  wire [10:0] _T_2922; // @[Mux.scala 31:69:@22709.4]
  wire [10:0] _T_2923; // @[Mux.scala 31:69:@22710.4]
  wire  _T_2928; // @[MemPrimitives.scala 110:210:@22717.4]
  wire  _T_2931; // @[MemPrimitives.scala 110:228:@22719.4]
  wire  _T_2934; // @[MemPrimitives.scala 110:210:@22721.4]
  wire  _T_2937; // @[MemPrimitives.scala 110:228:@22723.4]
  wire  _T_2940; // @[MemPrimitives.scala 110:210:@22725.4]
  wire  _T_2943; // @[MemPrimitives.scala 110:228:@22727.4]
  wire  _T_2946; // @[MemPrimitives.scala 110:210:@22729.4]
  wire  _T_2949; // @[MemPrimitives.scala 110:228:@22731.4]
  wire  _T_2952; // @[MemPrimitives.scala 110:210:@22733.4]
  wire  _T_2955; // @[MemPrimitives.scala 110:228:@22735.4]
  wire  _T_2958; // @[MemPrimitives.scala 110:210:@22737.4]
  wire  _T_2961; // @[MemPrimitives.scala 110:228:@22739.4]
  wire  _T_2964; // @[MemPrimitives.scala 110:210:@22741.4]
  wire  _T_2967; // @[MemPrimitives.scala 110:228:@22743.4]
  wire  _T_2970; // @[MemPrimitives.scala 110:210:@22745.4]
  wire  _T_2973; // @[MemPrimitives.scala 110:228:@22747.4]
  wire  _T_2976; // @[MemPrimitives.scala 110:210:@22749.4]
  wire  _T_2979; // @[MemPrimitives.scala 110:228:@22751.4]
  wire  _T_2981; // @[MemPrimitives.scala 126:35:@22765.4]
  wire  _T_2982; // @[MemPrimitives.scala 126:35:@22766.4]
  wire  _T_2983; // @[MemPrimitives.scala 126:35:@22767.4]
  wire  _T_2984; // @[MemPrimitives.scala 126:35:@22768.4]
  wire  _T_2985; // @[MemPrimitives.scala 126:35:@22769.4]
  wire  _T_2986; // @[MemPrimitives.scala 126:35:@22770.4]
  wire  _T_2987; // @[MemPrimitives.scala 126:35:@22771.4]
  wire  _T_2988; // @[MemPrimitives.scala 126:35:@22772.4]
  wire  _T_2989; // @[MemPrimitives.scala 126:35:@22773.4]
  wire [10:0] _T_2991; // @[Cat.scala 30:58:@22775.4]
  wire [10:0] _T_2993; // @[Cat.scala 30:58:@22777.4]
  wire [10:0] _T_2995; // @[Cat.scala 30:58:@22779.4]
  wire [10:0] _T_2997; // @[Cat.scala 30:58:@22781.4]
  wire [10:0] _T_2999; // @[Cat.scala 30:58:@22783.4]
  wire [10:0] _T_3001; // @[Cat.scala 30:58:@22785.4]
  wire [10:0] _T_3003; // @[Cat.scala 30:58:@22787.4]
  wire [10:0] _T_3005; // @[Cat.scala 30:58:@22789.4]
  wire [10:0] _T_3007; // @[Cat.scala 30:58:@22791.4]
  wire [10:0] _T_3008; // @[Mux.scala 31:69:@22792.4]
  wire [10:0] _T_3009; // @[Mux.scala 31:69:@22793.4]
  wire [10:0] _T_3010; // @[Mux.scala 31:69:@22794.4]
  wire [10:0] _T_3011; // @[Mux.scala 31:69:@22795.4]
  wire [10:0] _T_3012; // @[Mux.scala 31:69:@22796.4]
  wire [10:0] _T_3013; // @[Mux.scala 31:69:@22797.4]
  wire [10:0] _T_3014; // @[Mux.scala 31:69:@22798.4]
  wire [10:0] _T_3015; // @[Mux.scala 31:69:@22799.4]
  wire  _T_3023; // @[MemPrimitives.scala 110:228:@22808.4]
  wire  _T_3029; // @[MemPrimitives.scala 110:228:@22812.4]
  wire  _T_3035; // @[MemPrimitives.scala 110:228:@22816.4]
  wire  _T_3041; // @[MemPrimitives.scala 110:228:@22820.4]
  wire  _T_3047; // @[MemPrimitives.scala 110:228:@22824.4]
  wire  _T_3053; // @[MemPrimitives.scala 110:228:@22828.4]
  wire  _T_3059; // @[MemPrimitives.scala 110:228:@22832.4]
  wire  _T_3065; // @[MemPrimitives.scala 110:228:@22836.4]
  wire  _T_3071; // @[MemPrimitives.scala 110:228:@22840.4]
  wire  _T_3073; // @[MemPrimitives.scala 126:35:@22854.4]
  wire  _T_3074; // @[MemPrimitives.scala 126:35:@22855.4]
  wire  _T_3075; // @[MemPrimitives.scala 126:35:@22856.4]
  wire  _T_3076; // @[MemPrimitives.scala 126:35:@22857.4]
  wire  _T_3077; // @[MemPrimitives.scala 126:35:@22858.4]
  wire  _T_3078; // @[MemPrimitives.scala 126:35:@22859.4]
  wire  _T_3079; // @[MemPrimitives.scala 126:35:@22860.4]
  wire  _T_3080; // @[MemPrimitives.scala 126:35:@22861.4]
  wire  _T_3081; // @[MemPrimitives.scala 126:35:@22862.4]
  wire [10:0] _T_3083; // @[Cat.scala 30:58:@22864.4]
  wire [10:0] _T_3085; // @[Cat.scala 30:58:@22866.4]
  wire [10:0] _T_3087; // @[Cat.scala 30:58:@22868.4]
  wire [10:0] _T_3089; // @[Cat.scala 30:58:@22870.4]
  wire [10:0] _T_3091; // @[Cat.scala 30:58:@22872.4]
  wire [10:0] _T_3093; // @[Cat.scala 30:58:@22874.4]
  wire [10:0] _T_3095; // @[Cat.scala 30:58:@22876.4]
  wire [10:0] _T_3097; // @[Cat.scala 30:58:@22878.4]
  wire [10:0] _T_3099; // @[Cat.scala 30:58:@22880.4]
  wire [10:0] _T_3100; // @[Mux.scala 31:69:@22881.4]
  wire [10:0] _T_3101; // @[Mux.scala 31:69:@22882.4]
  wire [10:0] _T_3102; // @[Mux.scala 31:69:@22883.4]
  wire [10:0] _T_3103; // @[Mux.scala 31:69:@22884.4]
  wire [10:0] _T_3104; // @[Mux.scala 31:69:@22885.4]
  wire [10:0] _T_3105; // @[Mux.scala 31:69:@22886.4]
  wire [10:0] _T_3106; // @[Mux.scala 31:69:@22887.4]
  wire [10:0] _T_3107; // @[Mux.scala 31:69:@22888.4]
  wire  _T_3115; // @[MemPrimitives.scala 110:228:@22897.4]
  wire  _T_3121; // @[MemPrimitives.scala 110:228:@22901.4]
  wire  _T_3127; // @[MemPrimitives.scala 110:228:@22905.4]
  wire  _T_3133; // @[MemPrimitives.scala 110:228:@22909.4]
  wire  _T_3139; // @[MemPrimitives.scala 110:228:@22913.4]
  wire  _T_3145; // @[MemPrimitives.scala 110:228:@22917.4]
  wire  _T_3151; // @[MemPrimitives.scala 110:228:@22921.4]
  wire  _T_3157; // @[MemPrimitives.scala 110:228:@22925.4]
  wire  _T_3163; // @[MemPrimitives.scala 110:228:@22929.4]
  wire  _T_3165; // @[MemPrimitives.scala 126:35:@22943.4]
  wire  _T_3166; // @[MemPrimitives.scala 126:35:@22944.4]
  wire  _T_3167; // @[MemPrimitives.scala 126:35:@22945.4]
  wire  _T_3168; // @[MemPrimitives.scala 126:35:@22946.4]
  wire  _T_3169; // @[MemPrimitives.scala 126:35:@22947.4]
  wire  _T_3170; // @[MemPrimitives.scala 126:35:@22948.4]
  wire  _T_3171; // @[MemPrimitives.scala 126:35:@22949.4]
  wire  _T_3172; // @[MemPrimitives.scala 126:35:@22950.4]
  wire  _T_3173; // @[MemPrimitives.scala 126:35:@22951.4]
  wire [10:0] _T_3175; // @[Cat.scala 30:58:@22953.4]
  wire [10:0] _T_3177; // @[Cat.scala 30:58:@22955.4]
  wire [10:0] _T_3179; // @[Cat.scala 30:58:@22957.4]
  wire [10:0] _T_3181; // @[Cat.scala 30:58:@22959.4]
  wire [10:0] _T_3183; // @[Cat.scala 30:58:@22961.4]
  wire [10:0] _T_3185; // @[Cat.scala 30:58:@22963.4]
  wire [10:0] _T_3187; // @[Cat.scala 30:58:@22965.4]
  wire [10:0] _T_3189; // @[Cat.scala 30:58:@22967.4]
  wire [10:0] _T_3191; // @[Cat.scala 30:58:@22969.4]
  wire [10:0] _T_3192; // @[Mux.scala 31:69:@22970.4]
  wire [10:0] _T_3193; // @[Mux.scala 31:69:@22971.4]
  wire [10:0] _T_3194; // @[Mux.scala 31:69:@22972.4]
  wire [10:0] _T_3195; // @[Mux.scala 31:69:@22973.4]
  wire [10:0] _T_3196; // @[Mux.scala 31:69:@22974.4]
  wire [10:0] _T_3197; // @[Mux.scala 31:69:@22975.4]
  wire [10:0] _T_3198; // @[Mux.scala 31:69:@22976.4]
  wire [10:0] _T_3199; // @[Mux.scala 31:69:@22977.4]
  wire  _T_3207; // @[MemPrimitives.scala 110:228:@22986.4]
  wire  _T_3213; // @[MemPrimitives.scala 110:228:@22990.4]
  wire  _T_3219; // @[MemPrimitives.scala 110:228:@22994.4]
  wire  _T_3225; // @[MemPrimitives.scala 110:228:@22998.4]
  wire  _T_3231; // @[MemPrimitives.scala 110:228:@23002.4]
  wire  _T_3237; // @[MemPrimitives.scala 110:228:@23006.4]
  wire  _T_3243; // @[MemPrimitives.scala 110:228:@23010.4]
  wire  _T_3249; // @[MemPrimitives.scala 110:228:@23014.4]
  wire  _T_3255; // @[MemPrimitives.scala 110:228:@23018.4]
  wire  _T_3257; // @[MemPrimitives.scala 126:35:@23032.4]
  wire  _T_3258; // @[MemPrimitives.scala 126:35:@23033.4]
  wire  _T_3259; // @[MemPrimitives.scala 126:35:@23034.4]
  wire  _T_3260; // @[MemPrimitives.scala 126:35:@23035.4]
  wire  _T_3261; // @[MemPrimitives.scala 126:35:@23036.4]
  wire  _T_3262; // @[MemPrimitives.scala 126:35:@23037.4]
  wire  _T_3263; // @[MemPrimitives.scala 126:35:@23038.4]
  wire  _T_3264; // @[MemPrimitives.scala 126:35:@23039.4]
  wire  _T_3265; // @[MemPrimitives.scala 126:35:@23040.4]
  wire [10:0] _T_3267; // @[Cat.scala 30:58:@23042.4]
  wire [10:0] _T_3269; // @[Cat.scala 30:58:@23044.4]
  wire [10:0] _T_3271; // @[Cat.scala 30:58:@23046.4]
  wire [10:0] _T_3273; // @[Cat.scala 30:58:@23048.4]
  wire [10:0] _T_3275; // @[Cat.scala 30:58:@23050.4]
  wire [10:0] _T_3277; // @[Cat.scala 30:58:@23052.4]
  wire [10:0] _T_3279; // @[Cat.scala 30:58:@23054.4]
  wire [10:0] _T_3281; // @[Cat.scala 30:58:@23056.4]
  wire [10:0] _T_3283; // @[Cat.scala 30:58:@23058.4]
  wire [10:0] _T_3284; // @[Mux.scala 31:69:@23059.4]
  wire [10:0] _T_3285; // @[Mux.scala 31:69:@23060.4]
  wire [10:0] _T_3286; // @[Mux.scala 31:69:@23061.4]
  wire [10:0] _T_3287; // @[Mux.scala 31:69:@23062.4]
  wire [10:0] _T_3288; // @[Mux.scala 31:69:@23063.4]
  wire [10:0] _T_3289; // @[Mux.scala 31:69:@23064.4]
  wire [10:0] _T_3290; // @[Mux.scala 31:69:@23065.4]
  wire [10:0] _T_3291; // @[Mux.scala 31:69:@23066.4]
  wire  _T_3299; // @[MemPrimitives.scala 110:228:@23075.4]
  wire  _T_3305; // @[MemPrimitives.scala 110:228:@23079.4]
  wire  _T_3311; // @[MemPrimitives.scala 110:228:@23083.4]
  wire  _T_3317; // @[MemPrimitives.scala 110:228:@23087.4]
  wire  _T_3323; // @[MemPrimitives.scala 110:228:@23091.4]
  wire  _T_3329; // @[MemPrimitives.scala 110:228:@23095.4]
  wire  _T_3335; // @[MemPrimitives.scala 110:228:@23099.4]
  wire  _T_3341; // @[MemPrimitives.scala 110:228:@23103.4]
  wire  _T_3347; // @[MemPrimitives.scala 110:228:@23107.4]
  wire  _T_3349; // @[MemPrimitives.scala 126:35:@23121.4]
  wire  _T_3350; // @[MemPrimitives.scala 126:35:@23122.4]
  wire  _T_3351; // @[MemPrimitives.scala 126:35:@23123.4]
  wire  _T_3352; // @[MemPrimitives.scala 126:35:@23124.4]
  wire  _T_3353; // @[MemPrimitives.scala 126:35:@23125.4]
  wire  _T_3354; // @[MemPrimitives.scala 126:35:@23126.4]
  wire  _T_3355; // @[MemPrimitives.scala 126:35:@23127.4]
  wire  _T_3356; // @[MemPrimitives.scala 126:35:@23128.4]
  wire  _T_3357; // @[MemPrimitives.scala 126:35:@23129.4]
  wire [10:0] _T_3359; // @[Cat.scala 30:58:@23131.4]
  wire [10:0] _T_3361; // @[Cat.scala 30:58:@23133.4]
  wire [10:0] _T_3363; // @[Cat.scala 30:58:@23135.4]
  wire [10:0] _T_3365; // @[Cat.scala 30:58:@23137.4]
  wire [10:0] _T_3367; // @[Cat.scala 30:58:@23139.4]
  wire [10:0] _T_3369; // @[Cat.scala 30:58:@23141.4]
  wire [10:0] _T_3371; // @[Cat.scala 30:58:@23143.4]
  wire [10:0] _T_3373; // @[Cat.scala 30:58:@23145.4]
  wire [10:0] _T_3375; // @[Cat.scala 30:58:@23147.4]
  wire [10:0] _T_3376; // @[Mux.scala 31:69:@23148.4]
  wire [10:0] _T_3377; // @[Mux.scala 31:69:@23149.4]
  wire [10:0] _T_3378; // @[Mux.scala 31:69:@23150.4]
  wire [10:0] _T_3379; // @[Mux.scala 31:69:@23151.4]
  wire [10:0] _T_3380; // @[Mux.scala 31:69:@23152.4]
  wire [10:0] _T_3381; // @[Mux.scala 31:69:@23153.4]
  wire [10:0] _T_3382; // @[Mux.scala 31:69:@23154.4]
  wire [10:0] _T_3383; // @[Mux.scala 31:69:@23155.4]
  wire  _T_3479; // @[package.scala 96:25:@23284.4 package.scala 96:25:@23285.4]
  wire [31:0] _T_3483; // @[Mux.scala 31:69:@23294.4]
  wire  _T_3476; // @[package.scala 96:25:@23276.4 package.scala 96:25:@23277.4]
  wire [31:0] _T_3484; // @[Mux.scala 31:69:@23295.4]
  wire  _T_3473; // @[package.scala 96:25:@23268.4 package.scala 96:25:@23269.4]
  wire [31:0] _T_3485; // @[Mux.scala 31:69:@23296.4]
  wire  _T_3470; // @[package.scala 96:25:@23260.4 package.scala 96:25:@23261.4]
  wire [31:0] _T_3486; // @[Mux.scala 31:69:@23297.4]
  wire  _T_3467; // @[package.scala 96:25:@23252.4 package.scala 96:25:@23253.4]
  wire [31:0] _T_3487; // @[Mux.scala 31:69:@23298.4]
  wire  _T_3464; // @[package.scala 96:25:@23244.4 package.scala 96:25:@23245.4]
  wire [31:0] _T_3488; // @[Mux.scala 31:69:@23299.4]
  wire  _T_3461; // @[package.scala 96:25:@23236.4 package.scala 96:25:@23237.4]
  wire [31:0] _T_3489; // @[Mux.scala 31:69:@23300.4]
  wire  _T_3458; // @[package.scala 96:25:@23228.4 package.scala 96:25:@23229.4]
  wire [31:0] _T_3490; // @[Mux.scala 31:69:@23301.4]
  wire  _T_3455; // @[package.scala 96:25:@23220.4 package.scala 96:25:@23221.4]
  wire [31:0] _T_3491; // @[Mux.scala 31:69:@23302.4]
  wire  _T_3452; // @[package.scala 96:25:@23212.4 package.scala 96:25:@23213.4]
  wire [31:0] _T_3492; // @[Mux.scala 31:69:@23303.4]
  wire  _T_3449; // @[package.scala 96:25:@23204.4 package.scala 96:25:@23205.4]
  wire  _T_3586; // @[package.scala 96:25:@23428.4 package.scala 96:25:@23429.4]
  wire [31:0] _T_3590; // @[Mux.scala 31:69:@23438.4]
  wire  _T_3583; // @[package.scala 96:25:@23420.4 package.scala 96:25:@23421.4]
  wire [31:0] _T_3591; // @[Mux.scala 31:69:@23439.4]
  wire  _T_3580; // @[package.scala 96:25:@23412.4 package.scala 96:25:@23413.4]
  wire [31:0] _T_3592; // @[Mux.scala 31:69:@23440.4]
  wire  _T_3577; // @[package.scala 96:25:@23404.4 package.scala 96:25:@23405.4]
  wire [31:0] _T_3593; // @[Mux.scala 31:69:@23441.4]
  wire  _T_3574; // @[package.scala 96:25:@23396.4 package.scala 96:25:@23397.4]
  wire [31:0] _T_3594; // @[Mux.scala 31:69:@23442.4]
  wire  _T_3571; // @[package.scala 96:25:@23388.4 package.scala 96:25:@23389.4]
  wire [31:0] _T_3595; // @[Mux.scala 31:69:@23443.4]
  wire  _T_3568; // @[package.scala 96:25:@23380.4 package.scala 96:25:@23381.4]
  wire [31:0] _T_3596; // @[Mux.scala 31:69:@23444.4]
  wire  _T_3565; // @[package.scala 96:25:@23372.4 package.scala 96:25:@23373.4]
  wire [31:0] _T_3597; // @[Mux.scala 31:69:@23445.4]
  wire  _T_3562; // @[package.scala 96:25:@23364.4 package.scala 96:25:@23365.4]
  wire [31:0] _T_3598; // @[Mux.scala 31:69:@23446.4]
  wire  _T_3559; // @[package.scala 96:25:@23356.4 package.scala 96:25:@23357.4]
  wire [31:0] _T_3599; // @[Mux.scala 31:69:@23447.4]
  wire  _T_3556; // @[package.scala 96:25:@23348.4 package.scala 96:25:@23349.4]
  wire  _T_3693; // @[package.scala 96:25:@23572.4 package.scala 96:25:@23573.4]
  wire [31:0] _T_3697; // @[Mux.scala 31:69:@23582.4]
  wire  _T_3690; // @[package.scala 96:25:@23564.4 package.scala 96:25:@23565.4]
  wire [31:0] _T_3698; // @[Mux.scala 31:69:@23583.4]
  wire  _T_3687; // @[package.scala 96:25:@23556.4 package.scala 96:25:@23557.4]
  wire [31:0] _T_3699; // @[Mux.scala 31:69:@23584.4]
  wire  _T_3684; // @[package.scala 96:25:@23548.4 package.scala 96:25:@23549.4]
  wire [31:0] _T_3700; // @[Mux.scala 31:69:@23585.4]
  wire  _T_3681; // @[package.scala 96:25:@23540.4 package.scala 96:25:@23541.4]
  wire [31:0] _T_3701; // @[Mux.scala 31:69:@23586.4]
  wire  _T_3678; // @[package.scala 96:25:@23532.4 package.scala 96:25:@23533.4]
  wire [31:0] _T_3702; // @[Mux.scala 31:69:@23587.4]
  wire  _T_3675; // @[package.scala 96:25:@23524.4 package.scala 96:25:@23525.4]
  wire [31:0] _T_3703; // @[Mux.scala 31:69:@23588.4]
  wire  _T_3672; // @[package.scala 96:25:@23516.4 package.scala 96:25:@23517.4]
  wire [31:0] _T_3704; // @[Mux.scala 31:69:@23589.4]
  wire  _T_3669; // @[package.scala 96:25:@23508.4 package.scala 96:25:@23509.4]
  wire [31:0] _T_3705; // @[Mux.scala 31:69:@23590.4]
  wire  _T_3666; // @[package.scala 96:25:@23500.4 package.scala 96:25:@23501.4]
  wire [31:0] _T_3706; // @[Mux.scala 31:69:@23591.4]
  wire  _T_3663; // @[package.scala 96:25:@23492.4 package.scala 96:25:@23493.4]
  wire  _T_3800; // @[package.scala 96:25:@23716.4 package.scala 96:25:@23717.4]
  wire [31:0] _T_3804; // @[Mux.scala 31:69:@23726.4]
  wire  _T_3797; // @[package.scala 96:25:@23708.4 package.scala 96:25:@23709.4]
  wire [31:0] _T_3805; // @[Mux.scala 31:69:@23727.4]
  wire  _T_3794; // @[package.scala 96:25:@23700.4 package.scala 96:25:@23701.4]
  wire [31:0] _T_3806; // @[Mux.scala 31:69:@23728.4]
  wire  _T_3791; // @[package.scala 96:25:@23692.4 package.scala 96:25:@23693.4]
  wire [31:0] _T_3807; // @[Mux.scala 31:69:@23729.4]
  wire  _T_3788; // @[package.scala 96:25:@23684.4 package.scala 96:25:@23685.4]
  wire [31:0] _T_3808; // @[Mux.scala 31:69:@23730.4]
  wire  _T_3785; // @[package.scala 96:25:@23676.4 package.scala 96:25:@23677.4]
  wire [31:0] _T_3809; // @[Mux.scala 31:69:@23731.4]
  wire  _T_3782; // @[package.scala 96:25:@23668.4 package.scala 96:25:@23669.4]
  wire [31:0] _T_3810; // @[Mux.scala 31:69:@23732.4]
  wire  _T_3779; // @[package.scala 96:25:@23660.4 package.scala 96:25:@23661.4]
  wire [31:0] _T_3811; // @[Mux.scala 31:69:@23733.4]
  wire  _T_3776; // @[package.scala 96:25:@23652.4 package.scala 96:25:@23653.4]
  wire [31:0] _T_3812; // @[Mux.scala 31:69:@23734.4]
  wire  _T_3773; // @[package.scala 96:25:@23644.4 package.scala 96:25:@23645.4]
  wire [31:0] _T_3813; // @[Mux.scala 31:69:@23735.4]
  wire  _T_3770; // @[package.scala 96:25:@23636.4 package.scala 96:25:@23637.4]
  wire  _T_3907; // @[package.scala 96:25:@23860.4 package.scala 96:25:@23861.4]
  wire [31:0] _T_3911; // @[Mux.scala 31:69:@23870.4]
  wire  _T_3904; // @[package.scala 96:25:@23852.4 package.scala 96:25:@23853.4]
  wire [31:0] _T_3912; // @[Mux.scala 31:69:@23871.4]
  wire  _T_3901; // @[package.scala 96:25:@23844.4 package.scala 96:25:@23845.4]
  wire [31:0] _T_3913; // @[Mux.scala 31:69:@23872.4]
  wire  _T_3898; // @[package.scala 96:25:@23836.4 package.scala 96:25:@23837.4]
  wire [31:0] _T_3914; // @[Mux.scala 31:69:@23873.4]
  wire  _T_3895; // @[package.scala 96:25:@23828.4 package.scala 96:25:@23829.4]
  wire [31:0] _T_3915; // @[Mux.scala 31:69:@23874.4]
  wire  _T_3892; // @[package.scala 96:25:@23820.4 package.scala 96:25:@23821.4]
  wire [31:0] _T_3916; // @[Mux.scala 31:69:@23875.4]
  wire  _T_3889; // @[package.scala 96:25:@23812.4 package.scala 96:25:@23813.4]
  wire [31:0] _T_3917; // @[Mux.scala 31:69:@23876.4]
  wire  _T_3886; // @[package.scala 96:25:@23804.4 package.scala 96:25:@23805.4]
  wire [31:0] _T_3918; // @[Mux.scala 31:69:@23877.4]
  wire  _T_3883; // @[package.scala 96:25:@23796.4 package.scala 96:25:@23797.4]
  wire [31:0] _T_3919; // @[Mux.scala 31:69:@23878.4]
  wire  _T_3880; // @[package.scala 96:25:@23788.4 package.scala 96:25:@23789.4]
  wire [31:0] _T_3920; // @[Mux.scala 31:69:@23879.4]
  wire  _T_3877; // @[package.scala 96:25:@23780.4 package.scala 96:25:@23781.4]
  wire  _T_4014; // @[package.scala 96:25:@24004.4 package.scala 96:25:@24005.4]
  wire [31:0] _T_4018; // @[Mux.scala 31:69:@24014.4]
  wire  _T_4011; // @[package.scala 96:25:@23996.4 package.scala 96:25:@23997.4]
  wire [31:0] _T_4019; // @[Mux.scala 31:69:@24015.4]
  wire  _T_4008; // @[package.scala 96:25:@23988.4 package.scala 96:25:@23989.4]
  wire [31:0] _T_4020; // @[Mux.scala 31:69:@24016.4]
  wire  _T_4005; // @[package.scala 96:25:@23980.4 package.scala 96:25:@23981.4]
  wire [31:0] _T_4021; // @[Mux.scala 31:69:@24017.4]
  wire  _T_4002; // @[package.scala 96:25:@23972.4 package.scala 96:25:@23973.4]
  wire [31:0] _T_4022; // @[Mux.scala 31:69:@24018.4]
  wire  _T_3999; // @[package.scala 96:25:@23964.4 package.scala 96:25:@23965.4]
  wire [31:0] _T_4023; // @[Mux.scala 31:69:@24019.4]
  wire  _T_3996; // @[package.scala 96:25:@23956.4 package.scala 96:25:@23957.4]
  wire [31:0] _T_4024; // @[Mux.scala 31:69:@24020.4]
  wire  _T_3993; // @[package.scala 96:25:@23948.4 package.scala 96:25:@23949.4]
  wire [31:0] _T_4025; // @[Mux.scala 31:69:@24021.4]
  wire  _T_3990; // @[package.scala 96:25:@23940.4 package.scala 96:25:@23941.4]
  wire [31:0] _T_4026; // @[Mux.scala 31:69:@24022.4]
  wire  _T_3987; // @[package.scala 96:25:@23932.4 package.scala 96:25:@23933.4]
  wire [31:0] _T_4027; // @[Mux.scala 31:69:@24023.4]
  wire  _T_3984; // @[package.scala 96:25:@23924.4 package.scala 96:25:@23925.4]
  wire  _T_4121; // @[package.scala 96:25:@24148.4 package.scala 96:25:@24149.4]
  wire [31:0] _T_4125; // @[Mux.scala 31:69:@24158.4]
  wire  _T_4118; // @[package.scala 96:25:@24140.4 package.scala 96:25:@24141.4]
  wire [31:0] _T_4126; // @[Mux.scala 31:69:@24159.4]
  wire  _T_4115; // @[package.scala 96:25:@24132.4 package.scala 96:25:@24133.4]
  wire [31:0] _T_4127; // @[Mux.scala 31:69:@24160.4]
  wire  _T_4112; // @[package.scala 96:25:@24124.4 package.scala 96:25:@24125.4]
  wire [31:0] _T_4128; // @[Mux.scala 31:69:@24161.4]
  wire  _T_4109; // @[package.scala 96:25:@24116.4 package.scala 96:25:@24117.4]
  wire [31:0] _T_4129; // @[Mux.scala 31:69:@24162.4]
  wire  _T_4106; // @[package.scala 96:25:@24108.4 package.scala 96:25:@24109.4]
  wire [31:0] _T_4130; // @[Mux.scala 31:69:@24163.4]
  wire  _T_4103; // @[package.scala 96:25:@24100.4 package.scala 96:25:@24101.4]
  wire [31:0] _T_4131; // @[Mux.scala 31:69:@24164.4]
  wire  _T_4100; // @[package.scala 96:25:@24092.4 package.scala 96:25:@24093.4]
  wire [31:0] _T_4132; // @[Mux.scala 31:69:@24165.4]
  wire  _T_4097; // @[package.scala 96:25:@24084.4 package.scala 96:25:@24085.4]
  wire [31:0] _T_4133; // @[Mux.scala 31:69:@24166.4]
  wire  _T_4094; // @[package.scala 96:25:@24076.4 package.scala 96:25:@24077.4]
  wire [31:0] _T_4134; // @[Mux.scala 31:69:@24167.4]
  wire  _T_4091; // @[package.scala 96:25:@24068.4 package.scala 96:25:@24069.4]
  wire  _T_4228; // @[package.scala 96:25:@24292.4 package.scala 96:25:@24293.4]
  wire [31:0] _T_4232; // @[Mux.scala 31:69:@24302.4]
  wire  _T_4225; // @[package.scala 96:25:@24284.4 package.scala 96:25:@24285.4]
  wire [31:0] _T_4233; // @[Mux.scala 31:69:@24303.4]
  wire  _T_4222; // @[package.scala 96:25:@24276.4 package.scala 96:25:@24277.4]
  wire [31:0] _T_4234; // @[Mux.scala 31:69:@24304.4]
  wire  _T_4219; // @[package.scala 96:25:@24268.4 package.scala 96:25:@24269.4]
  wire [31:0] _T_4235; // @[Mux.scala 31:69:@24305.4]
  wire  _T_4216; // @[package.scala 96:25:@24260.4 package.scala 96:25:@24261.4]
  wire [31:0] _T_4236; // @[Mux.scala 31:69:@24306.4]
  wire  _T_4213; // @[package.scala 96:25:@24252.4 package.scala 96:25:@24253.4]
  wire [31:0] _T_4237; // @[Mux.scala 31:69:@24307.4]
  wire  _T_4210; // @[package.scala 96:25:@24244.4 package.scala 96:25:@24245.4]
  wire [31:0] _T_4238; // @[Mux.scala 31:69:@24308.4]
  wire  _T_4207; // @[package.scala 96:25:@24236.4 package.scala 96:25:@24237.4]
  wire [31:0] _T_4239; // @[Mux.scala 31:69:@24309.4]
  wire  _T_4204; // @[package.scala 96:25:@24228.4 package.scala 96:25:@24229.4]
  wire [31:0] _T_4240; // @[Mux.scala 31:69:@24310.4]
  wire  _T_4201; // @[package.scala 96:25:@24220.4 package.scala 96:25:@24221.4]
  wire [31:0] _T_4241; // @[Mux.scala 31:69:@24311.4]
  wire  _T_4198; // @[package.scala 96:25:@24212.4 package.scala 96:25:@24213.4]
  wire  _T_4335; // @[package.scala 96:25:@24436.4 package.scala 96:25:@24437.4]
  wire [31:0] _T_4339; // @[Mux.scala 31:69:@24446.4]
  wire  _T_4332; // @[package.scala 96:25:@24428.4 package.scala 96:25:@24429.4]
  wire [31:0] _T_4340; // @[Mux.scala 31:69:@24447.4]
  wire  _T_4329; // @[package.scala 96:25:@24420.4 package.scala 96:25:@24421.4]
  wire [31:0] _T_4341; // @[Mux.scala 31:69:@24448.4]
  wire  _T_4326; // @[package.scala 96:25:@24412.4 package.scala 96:25:@24413.4]
  wire [31:0] _T_4342; // @[Mux.scala 31:69:@24449.4]
  wire  _T_4323; // @[package.scala 96:25:@24404.4 package.scala 96:25:@24405.4]
  wire [31:0] _T_4343; // @[Mux.scala 31:69:@24450.4]
  wire  _T_4320; // @[package.scala 96:25:@24396.4 package.scala 96:25:@24397.4]
  wire [31:0] _T_4344; // @[Mux.scala 31:69:@24451.4]
  wire  _T_4317; // @[package.scala 96:25:@24388.4 package.scala 96:25:@24389.4]
  wire [31:0] _T_4345; // @[Mux.scala 31:69:@24452.4]
  wire  _T_4314; // @[package.scala 96:25:@24380.4 package.scala 96:25:@24381.4]
  wire [31:0] _T_4346; // @[Mux.scala 31:69:@24453.4]
  wire  _T_4311; // @[package.scala 96:25:@24372.4 package.scala 96:25:@24373.4]
  wire [31:0] _T_4347; // @[Mux.scala 31:69:@24454.4]
  wire  _T_4308; // @[package.scala 96:25:@24364.4 package.scala 96:25:@24365.4]
  wire [31:0] _T_4348; // @[Mux.scala 31:69:@24455.4]
  wire  _T_4305; // @[package.scala 96:25:@24356.4 package.scala 96:25:@24357.4]
  wire  _T_4442; // @[package.scala 96:25:@24580.4 package.scala 96:25:@24581.4]
  wire [31:0] _T_4446; // @[Mux.scala 31:69:@24590.4]
  wire  _T_4439; // @[package.scala 96:25:@24572.4 package.scala 96:25:@24573.4]
  wire [31:0] _T_4447; // @[Mux.scala 31:69:@24591.4]
  wire  _T_4436; // @[package.scala 96:25:@24564.4 package.scala 96:25:@24565.4]
  wire [31:0] _T_4448; // @[Mux.scala 31:69:@24592.4]
  wire  _T_4433; // @[package.scala 96:25:@24556.4 package.scala 96:25:@24557.4]
  wire [31:0] _T_4449; // @[Mux.scala 31:69:@24593.4]
  wire  _T_4430; // @[package.scala 96:25:@24548.4 package.scala 96:25:@24549.4]
  wire [31:0] _T_4450; // @[Mux.scala 31:69:@24594.4]
  wire  _T_4427; // @[package.scala 96:25:@24540.4 package.scala 96:25:@24541.4]
  wire [31:0] _T_4451; // @[Mux.scala 31:69:@24595.4]
  wire  _T_4424; // @[package.scala 96:25:@24532.4 package.scala 96:25:@24533.4]
  wire [31:0] _T_4452; // @[Mux.scala 31:69:@24596.4]
  wire  _T_4421; // @[package.scala 96:25:@24524.4 package.scala 96:25:@24525.4]
  wire [31:0] _T_4453; // @[Mux.scala 31:69:@24597.4]
  wire  _T_4418; // @[package.scala 96:25:@24516.4 package.scala 96:25:@24517.4]
  wire [31:0] _T_4454; // @[Mux.scala 31:69:@24598.4]
  wire  _T_4415; // @[package.scala 96:25:@24508.4 package.scala 96:25:@24509.4]
  wire [31:0] _T_4455; // @[Mux.scala 31:69:@24599.4]
  wire  _T_4412; // @[package.scala 96:25:@24500.4 package.scala 96:25:@24501.4]
  wire  _T_4549; // @[package.scala 96:25:@24724.4 package.scala 96:25:@24725.4]
  wire [31:0] _T_4553; // @[Mux.scala 31:69:@24734.4]
  wire  _T_4546; // @[package.scala 96:25:@24716.4 package.scala 96:25:@24717.4]
  wire [31:0] _T_4554; // @[Mux.scala 31:69:@24735.4]
  wire  _T_4543; // @[package.scala 96:25:@24708.4 package.scala 96:25:@24709.4]
  wire [31:0] _T_4555; // @[Mux.scala 31:69:@24736.4]
  wire  _T_4540; // @[package.scala 96:25:@24700.4 package.scala 96:25:@24701.4]
  wire [31:0] _T_4556; // @[Mux.scala 31:69:@24737.4]
  wire  _T_4537; // @[package.scala 96:25:@24692.4 package.scala 96:25:@24693.4]
  wire [31:0] _T_4557; // @[Mux.scala 31:69:@24738.4]
  wire  _T_4534; // @[package.scala 96:25:@24684.4 package.scala 96:25:@24685.4]
  wire [31:0] _T_4558; // @[Mux.scala 31:69:@24739.4]
  wire  _T_4531; // @[package.scala 96:25:@24676.4 package.scala 96:25:@24677.4]
  wire [31:0] _T_4559; // @[Mux.scala 31:69:@24740.4]
  wire  _T_4528; // @[package.scala 96:25:@24668.4 package.scala 96:25:@24669.4]
  wire [31:0] _T_4560; // @[Mux.scala 31:69:@24741.4]
  wire  _T_4525; // @[package.scala 96:25:@24660.4 package.scala 96:25:@24661.4]
  wire [31:0] _T_4561; // @[Mux.scala 31:69:@24742.4]
  wire  _T_4522; // @[package.scala 96:25:@24652.4 package.scala 96:25:@24653.4]
  wire [31:0] _T_4562; // @[Mux.scala 31:69:@24743.4]
  wire  _T_4519; // @[package.scala 96:25:@24644.4 package.scala 96:25:@24645.4]
  wire  _T_4656; // @[package.scala 96:25:@24868.4 package.scala 96:25:@24869.4]
  wire [31:0] _T_4660; // @[Mux.scala 31:69:@24878.4]
  wire  _T_4653; // @[package.scala 96:25:@24860.4 package.scala 96:25:@24861.4]
  wire [31:0] _T_4661; // @[Mux.scala 31:69:@24879.4]
  wire  _T_4650; // @[package.scala 96:25:@24852.4 package.scala 96:25:@24853.4]
  wire [31:0] _T_4662; // @[Mux.scala 31:69:@24880.4]
  wire  _T_4647; // @[package.scala 96:25:@24844.4 package.scala 96:25:@24845.4]
  wire [31:0] _T_4663; // @[Mux.scala 31:69:@24881.4]
  wire  _T_4644; // @[package.scala 96:25:@24836.4 package.scala 96:25:@24837.4]
  wire [31:0] _T_4664; // @[Mux.scala 31:69:@24882.4]
  wire  _T_4641; // @[package.scala 96:25:@24828.4 package.scala 96:25:@24829.4]
  wire [31:0] _T_4665; // @[Mux.scala 31:69:@24883.4]
  wire  _T_4638; // @[package.scala 96:25:@24820.4 package.scala 96:25:@24821.4]
  wire [31:0] _T_4666; // @[Mux.scala 31:69:@24884.4]
  wire  _T_4635; // @[package.scala 96:25:@24812.4 package.scala 96:25:@24813.4]
  wire [31:0] _T_4667; // @[Mux.scala 31:69:@24885.4]
  wire  _T_4632; // @[package.scala 96:25:@24804.4 package.scala 96:25:@24805.4]
  wire [31:0] _T_4668; // @[Mux.scala 31:69:@24886.4]
  wire  _T_4629; // @[package.scala 96:25:@24796.4 package.scala 96:25:@24797.4]
  wire [31:0] _T_4669; // @[Mux.scala 31:69:@24887.4]
  wire  _T_4626; // @[package.scala 96:25:@24788.4 package.scala 96:25:@24789.4]
  wire  _T_4763; // @[package.scala 96:25:@25012.4 package.scala 96:25:@25013.4]
  wire [31:0] _T_4767; // @[Mux.scala 31:69:@25022.4]
  wire  _T_4760; // @[package.scala 96:25:@25004.4 package.scala 96:25:@25005.4]
  wire [31:0] _T_4768; // @[Mux.scala 31:69:@25023.4]
  wire  _T_4757; // @[package.scala 96:25:@24996.4 package.scala 96:25:@24997.4]
  wire [31:0] _T_4769; // @[Mux.scala 31:69:@25024.4]
  wire  _T_4754; // @[package.scala 96:25:@24988.4 package.scala 96:25:@24989.4]
  wire [31:0] _T_4770; // @[Mux.scala 31:69:@25025.4]
  wire  _T_4751; // @[package.scala 96:25:@24980.4 package.scala 96:25:@24981.4]
  wire [31:0] _T_4771; // @[Mux.scala 31:69:@25026.4]
  wire  _T_4748; // @[package.scala 96:25:@24972.4 package.scala 96:25:@24973.4]
  wire [31:0] _T_4772; // @[Mux.scala 31:69:@25027.4]
  wire  _T_4745; // @[package.scala 96:25:@24964.4 package.scala 96:25:@24965.4]
  wire [31:0] _T_4773; // @[Mux.scala 31:69:@25028.4]
  wire  _T_4742; // @[package.scala 96:25:@24956.4 package.scala 96:25:@24957.4]
  wire [31:0] _T_4774; // @[Mux.scala 31:69:@25029.4]
  wire  _T_4739; // @[package.scala 96:25:@24948.4 package.scala 96:25:@24949.4]
  wire [31:0] _T_4775; // @[Mux.scala 31:69:@25030.4]
  wire  _T_4736; // @[package.scala 96:25:@24940.4 package.scala 96:25:@24941.4]
  wire [31:0] _T_4776; // @[Mux.scala 31:69:@25031.4]
  wire  _T_4733; // @[package.scala 96:25:@24932.4 package.scala 96:25:@24933.4]
  wire  _T_4870; // @[package.scala 96:25:@25156.4 package.scala 96:25:@25157.4]
  wire [31:0] _T_4874; // @[Mux.scala 31:69:@25166.4]
  wire  _T_4867; // @[package.scala 96:25:@25148.4 package.scala 96:25:@25149.4]
  wire [31:0] _T_4875; // @[Mux.scala 31:69:@25167.4]
  wire  _T_4864; // @[package.scala 96:25:@25140.4 package.scala 96:25:@25141.4]
  wire [31:0] _T_4876; // @[Mux.scala 31:69:@25168.4]
  wire  _T_4861; // @[package.scala 96:25:@25132.4 package.scala 96:25:@25133.4]
  wire [31:0] _T_4877; // @[Mux.scala 31:69:@25169.4]
  wire  _T_4858; // @[package.scala 96:25:@25124.4 package.scala 96:25:@25125.4]
  wire [31:0] _T_4878; // @[Mux.scala 31:69:@25170.4]
  wire  _T_4855; // @[package.scala 96:25:@25116.4 package.scala 96:25:@25117.4]
  wire [31:0] _T_4879; // @[Mux.scala 31:69:@25171.4]
  wire  _T_4852; // @[package.scala 96:25:@25108.4 package.scala 96:25:@25109.4]
  wire [31:0] _T_4880; // @[Mux.scala 31:69:@25172.4]
  wire  _T_4849; // @[package.scala 96:25:@25100.4 package.scala 96:25:@25101.4]
  wire [31:0] _T_4881; // @[Mux.scala 31:69:@25173.4]
  wire  _T_4846; // @[package.scala 96:25:@25092.4 package.scala 96:25:@25093.4]
  wire [31:0] _T_4882; // @[Mux.scala 31:69:@25174.4]
  wire  _T_4843; // @[package.scala 96:25:@25084.4 package.scala 96:25:@25085.4]
  wire [31:0] _T_4883; // @[Mux.scala 31:69:@25175.4]
  wire  _T_4840; // @[package.scala 96:25:@25076.4 package.scala 96:25:@25077.4]
  wire  _T_4977; // @[package.scala 96:25:@25300.4 package.scala 96:25:@25301.4]
  wire [31:0] _T_4981; // @[Mux.scala 31:69:@25310.4]
  wire  _T_4974; // @[package.scala 96:25:@25292.4 package.scala 96:25:@25293.4]
  wire [31:0] _T_4982; // @[Mux.scala 31:69:@25311.4]
  wire  _T_4971; // @[package.scala 96:25:@25284.4 package.scala 96:25:@25285.4]
  wire [31:0] _T_4983; // @[Mux.scala 31:69:@25312.4]
  wire  _T_4968; // @[package.scala 96:25:@25276.4 package.scala 96:25:@25277.4]
  wire [31:0] _T_4984; // @[Mux.scala 31:69:@25313.4]
  wire  _T_4965; // @[package.scala 96:25:@25268.4 package.scala 96:25:@25269.4]
  wire [31:0] _T_4985; // @[Mux.scala 31:69:@25314.4]
  wire  _T_4962; // @[package.scala 96:25:@25260.4 package.scala 96:25:@25261.4]
  wire [31:0] _T_4986; // @[Mux.scala 31:69:@25315.4]
  wire  _T_4959; // @[package.scala 96:25:@25252.4 package.scala 96:25:@25253.4]
  wire [31:0] _T_4987; // @[Mux.scala 31:69:@25316.4]
  wire  _T_4956; // @[package.scala 96:25:@25244.4 package.scala 96:25:@25245.4]
  wire [31:0] _T_4988; // @[Mux.scala 31:69:@25317.4]
  wire  _T_4953; // @[package.scala 96:25:@25236.4 package.scala 96:25:@25237.4]
  wire [31:0] _T_4989; // @[Mux.scala 31:69:@25318.4]
  wire  _T_4950; // @[package.scala 96:25:@25228.4 package.scala 96:25:@25229.4]
  wire [31:0] _T_4990; // @[Mux.scala 31:69:@25319.4]
  wire  _T_4947; // @[package.scala 96:25:@25220.4 package.scala 96:25:@25221.4]
  wire  _T_5084; // @[package.scala 96:25:@25444.4 package.scala 96:25:@25445.4]
  wire [31:0] _T_5088; // @[Mux.scala 31:69:@25454.4]
  wire  _T_5081; // @[package.scala 96:25:@25436.4 package.scala 96:25:@25437.4]
  wire [31:0] _T_5089; // @[Mux.scala 31:69:@25455.4]
  wire  _T_5078; // @[package.scala 96:25:@25428.4 package.scala 96:25:@25429.4]
  wire [31:0] _T_5090; // @[Mux.scala 31:69:@25456.4]
  wire  _T_5075; // @[package.scala 96:25:@25420.4 package.scala 96:25:@25421.4]
  wire [31:0] _T_5091; // @[Mux.scala 31:69:@25457.4]
  wire  _T_5072; // @[package.scala 96:25:@25412.4 package.scala 96:25:@25413.4]
  wire [31:0] _T_5092; // @[Mux.scala 31:69:@25458.4]
  wire  _T_5069; // @[package.scala 96:25:@25404.4 package.scala 96:25:@25405.4]
  wire [31:0] _T_5093; // @[Mux.scala 31:69:@25459.4]
  wire  _T_5066; // @[package.scala 96:25:@25396.4 package.scala 96:25:@25397.4]
  wire [31:0] _T_5094; // @[Mux.scala 31:69:@25460.4]
  wire  _T_5063; // @[package.scala 96:25:@25388.4 package.scala 96:25:@25389.4]
  wire [31:0] _T_5095; // @[Mux.scala 31:69:@25461.4]
  wire  _T_5060; // @[package.scala 96:25:@25380.4 package.scala 96:25:@25381.4]
  wire [31:0] _T_5096; // @[Mux.scala 31:69:@25462.4]
  wire  _T_5057; // @[package.scala 96:25:@25372.4 package.scala 96:25:@25373.4]
  wire [31:0] _T_5097; // @[Mux.scala 31:69:@25463.4]
  wire  _T_5054; // @[package.scala 96:25:@25364.4 package.scala 96:25:@25365.4]
  wire  _T_5191; // @[package.scala 96:25:@25588.4 package.scala 96:25:@25589.4]
  wire [31:0] _T_5195; // @[Mux.scala 31:69:@25598.4]
  wire  _T_5188; // @[package.scala 96:25:@25580.4 package.scala 96:25:@25581.4]
  wire [31:0] _T_5196; // @[Mux.scala 31:69:@25599.4]
  wire  _T_5185; // @[package.scala 96:25:@25572.4 package.scala 96:25:@25573.4]
  wire [31:0] _T_5197; // @[Mux.scala 31:69:@25600.4]
  wire  _T_5182; // @[package.scala 96:25:@25564.4 package.scala 96:25:@25565.4]
  wire [31:0] _T_5198; // @[Mux.scala 31:69:@25601.4]
  wire  _T_5179; // @[package.scala 96:25:@25556.4 package.scala 96:25:@25557.4]
  wire [31:0] _T_5199; // @[Mux.scala 31:69:@25602.4]
  wire  _T_5176; // @[package.scala 96:25:@25548.4 package.scala 96:25:@25549.4]
  wire [31:0] _T_5200; // @[Mux.scala 31:69:@25603.4]
  wire  _T_5173; // @[package.scala 96:25:@25540.4 package.scala 96:25:@25541.4]
  wire [31:0] _T_5201; // @[Mux.scala 31:69:@25604.4]
  wire  _T_5170; // @[package.scala 96:25:@25532.4 package.scala 96:25:@25533.4]
  wire [31:0] _T_5202; // @[Mux.scala 31:69:@25605.4]
  wire  _T_5167; // @[package.scala 96:25:@25524.4 package.scala 96:25:@25525.4]
  wire [31:0] _T_5203; // @[Mux.scala 31:69:@25606.4]
  wire  _T_5164; // @[package.scala 96:25:@25516.4 package.scala 96:25:@25517.4]
  wire [31:0] _T_5204; // @[Mux.scala 31:69:@25607.4]
  wire  _T_5161; // @[package.scala 96:25:@25508.4 package.scala 96:25:@25509.4]
  wire  _T_5298; // @[package.scala 96:25:@25732.4 package.scala 96:25:@25733.4]
  wire [31:0] _T_5302; // @[Mux.scala 31:69:@25742.4]
  wire  _T_5295; // @[package.scala 96:25:@25724.4 package.scala 96:25:@25725.4]
  wire [31:0] _T_5303; // @[Mux.scala 31:69:@25743.4]
  wire  _T_5292; // @[package.scala 96:25:@25716.4 package.scala 96:25:@25717.4]
  wire [31:0] _T_5304; // @[Mux.scala 31:69:@25744.4]
  wire  _T_5289; // @[package.scala 96:25:@25708.4 package.scala 96:25:@25709.4]
  wire [31:0] _T_5305; // @[Mux.scala 31:69:@25745.4]
  wire  _T_5286; // @[package.scala 96:25:@25700.4 package.scala 96:25:@25701.4]
  wire [31:0] _T_5306; // @[Mux.scala 31:69:@25746.4]
  wire  _T_5283; // @[package.scala 96:25:@25692.4 package.scala 96:25:@25693.4]
  wire [31:0] _T_5307; // @[Mux.scala 31:69:@25747.4]
  wire  _T_5280; // @[package.scala 96:25:@25684.4 package.scala 96:25:@25685.4]
  wire [31:0] _T_5308; // @[Mux.scala 31:69:@25748.4]
  wire  _T_5277; // @[package.scala 96:25:@25676.4 package.scala 96:25:@25677.4]
  wire [31:0] _T_5309; // @[Mux.scala 31:69:@25749.4]
  wire  _T_5274; // @[package.scala 96:25:@25668.4 package.scala 96:25:@25669.4]
  wire [31:0] _T_5310; // @[Mux.scala 31:69:@25750.4]
  wire  _T_5271; // @[package.scala 96:25:@25660.4 package.scala 96:25:@25661.4]
  wire [31:0] _T_5311; // @[Mux.scala 31:69:@25751.4]
  wire  _T_5268; // @[package.scala 96:25:@25652.4 package.scala 96:25:@25653.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@20186.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@20202.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@20218.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@20234.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@20250.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@20266.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@20282.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@20298.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@20314.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@20330.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@20346.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@20362.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_5 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@20378.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_5 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@20394.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_5 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@20410.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_5 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@20426.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  Mem1D_5 Mem1D_16 ( // @[MemPrimitives.scala 64:21:@20442.4]
    .clock(Mem1D_16_clock),
    .reset(Mem1D_16_reset),
    .io_r_ofs_0(Mem1D_16_io_r_ofs_0),
    .io_r_backpressure(Mem1D_16_io_r_backpressure),
    .io_w_ofs_0(Mem1D_16_io_w_ofs_0),
    .io_w_data_0(Mem1D_16_io_w_data_0),
    .io_w_en_0(Mem1D_16_io_w_en_0),
    .io_output(Mem1D_16_io_output)
  );
  Mem1D_5 Mem1D_17 ( // @[MemPrimitives.scala 64:21:@20458.4]
    .clock(Mem1D_17_clock),
    .reset(Mem1D_17_reset),
    .io_r_ofs_0(Mem1D_17_io_r_ofs_0),
    .io_r_backpressure(Mem1D_17_io_r_backpressure),
    .io_w_ofs_0(Mem1D_17_io_w_ofs_0),
    .io_w_data_0(Mem1D_17_io_w_data_0),
    .io_w_en_0(Mem1D_17_io_w_en_0),
    .io_output(Mem1D_17_io_output)
  );
  Mem1D_5 Mem1D_18 ( // @[MemPrimitives.scala 64:21:@20474.4]
    .clock(Mem1D_18_clock),
    .reset(Mem1D_18_reset),
    .io_r_ofs_0(Mem1D_18_io_r_ofs_0),
    .io_r_backpressure(Mem1D_18_io_r_backpressure),
    .io_w_ofs_0(Mem1D_18_io_w_ofs_0),
    .io_w_data_0(Mem1D_18_io_w_data_0),
    .io_w_en_0(Mem1D_18_io_w_en_0),
    .io_output(Mem1D_18_io_output)
  );
  Mem1D_5 Mem1D_19 ( // @[MemPrimitives.scala 64:21:@20490.4]
    .clock(Mem1D_19_clock),
    .reset(Mem1D_19_reset),
    .io_r_ofs_0(Mem1D_19_io_r_ofs_0),
    .io_r_backpressure(Mem1D_19_io_r_backpressure),
    .io_w_ofs_0(Mem1D_19_io_w_ofs_0),
    .io_w_data_0(Mem1D_19_io_w_data_0),
    .io_w_en_0(Mem1D_19_io_w_en_0),
    .io_output(Mem1D_19_io_output)
  );
  Mem1D_5 Mem1D_20 ( // @[MemPrimitives.scala 64:21:@20506.4]
    .clock(Mem1D_20_clock),
    .reset(Mem1D_20_reset),
    .io_r_ofs_0(Mem1D_20_io_r_ofs_0),
    .io_r_backpressure(Mem1D_20_io_r_backpressure),
    .io_w_ofs_0(Mem1D_20_io_w_ofs_0),
    .io_w_data_0(Mem1D_20_io_w_data_0),
    .io_w_en_0(Mem1D_20_io_w_en_0),
    .io_output(Mem1D_20_io_output)
  );
  Mem1D_5 Mem1D_21 ( // @[MemPrimitives.scala 64:21:@20522.4]
    .clock(Mem1D_21_clock),
    .reset(Mem1D_21_reset),
    .io_r_ofs_0(Mem1D_21_io_r_ofs_0),
    .io_r_backpressure(Mem1D_21_io_r_backpressure),
    .io_w_ofs_0(Mem1D_21_io_w_ofs_0),
    .io_w_data_0(Mem1D_21_io_w_data_0),
    .io_w_en_0(Mem1D_21_io_w_en_0),
    .io_output(Mem1D_21_io_output)
  );
  Mem1D_5 Mem1D_22 ( // @[MemPrimitives.scala 64:21:@20538.4]
    .clock(Mem1D_22_clock),
    .reset(Mem1D_22_reset),
    .io_r_ofs_0(Mem1D_22_io_r_ofs_0),
    .io_r_backpressure(Mem1D_22_io_r_backpressure),
    .io_w_ofs_0(Mem1D_22_io_w_ofs_0),
    .io_w_data_0(Mem1D_22_io_w_data_0),
    .io_w_en_0(Mem1D_22_io_w_en_0),
    .io_output(Mem1D_22_io_output)
  );
  Mem1D_5 Mem1D_23 ( // @[MemPrimitives.scala 64:21:@20554.4]
    .clock(Mem1D_23_clock),
    .reset(Mem1D_23_reset),
    .io_r_ofs_0(Mem1D_23_io_r_ofs_0),
    .io_r_backpressure(Mem1D_23_io_r_backpressure),
    .io_w_ofs_0(Mem1D_23_io_w_ofs_0),
    .io_w_data_0(Mem1D_23_io_w_data_0),
    .io_w_en_0(Mem1D_23_io_w_en_0),
    .io_output(Mem1D_23_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 124:33:@21062.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_ins_6(StickySelects_io_ins_6),
    .io_ins_7(StickySelects_io_ins_7),
    .io_ins_8(StickySelects_io_ins_8),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5),
    .io_outs_6(StickySelects_io_outs_6),
    .io_outs_7(StickySelects_io_outs_7),
    .io_outs_8(StickySelects_io_outs_8)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@21151.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_ins_6(StickySelects_1_io_ins_6),
    .io_ins_7(StickySelects_1_io_ins_7),
    .io_ins_8(StickySelects_1_io_ins_8),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5),
    .io_outs_6(StickySelects_1_io_outs_6),
    .io_outs_7(StickySelects_1_io_outs_7),
    .io_outs_8(StickySelects_1_io_outs_8)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@21240.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_ins_8(StickySelects_2_io_ins_8),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7),
    .io_outs_8(StickySelects_2_io_outs_8)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@21329.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_ins_8(StickySelects_3_io_ins_8),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7),
    .io_outs_8(StickySelects_3_io_outs_8)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@21418.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_ins_6(StickySelects_4_io_ins_6),
    .io_ins_7(StickySelects_4_io_ins_7),
    .io_ins_8(StickySelects_4_io_ins_8),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5),
    .io_outs_6(StickySelects_4_io_outs_6),
    .io_outs_7(StickySelects_4_io_outs_7),
    .io_outs_8(StickySelects_4_io_outs_8)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@21507.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_ins_6(StickySelects_5_io_ins_6),
    .io_ins_7(StickySelects_5_io_ins_7),
    .io_ins_8(StickySelects_5_io_ins_8),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5),
    .io_outs_6(StickySelects_5_io_outs_6),
    .io_outs_7(StickySelects_5_io_outs_7),
    .io_outs_8(StickySelects_5_io_outs_8)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@21596.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_ins_8(StickySelects_6_io_ins_8),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7),
    .io_outs_8(StickySelects_6_io_outs_8)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@21685.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_ins_8(StickySelects_7_io_ins_8),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7),
    .io_outs_8(StickySelects_7_io_outs_8)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@21774.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_ins_6(StickySelects_8_io_ins_6),
    .io_ins_7(StickySelects_8_io_ins_7),
    .io_ins_8(StickySelects_8_io_ins_8),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5),
    .io_outs_6(StickySelects_8_io_outs_6),
    .io_outs_7(StickySelects_8_io_outs_7),
    .io_outs_8(StickySelects_8_io_outs_8)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@21863.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_ins_6(StickySelects_9_io_ins_6),
    .io_ins_7(StickySelects_9_io_ins_7),
    .io_ins_8(StickySelects_9_io_ins_8),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5),
    .io_outs_6(StickySelects_9_io_outs_6),
    .io_outs_7(StickySelects_9_io_outs_7),
    .io_outs_8(StickySelects_9_io_outs_8)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@21952.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_ins_8(StickySelects_10_io_ins_8),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7),
    .io_outs_8(StickySelects_10_io_outs_8)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@22041.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_ins_8(StickySelects_11_io_ins_8),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7),
    .io_outs_8(StickySelects_11_io_outs_8)
  );
  StickySelects_1 StickySelects_12 ( // @[MemPrimitives.scala 124:33:@22130.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_ins_6(StickySelects_12_io_ins_6),
    .io_ins_7(StickySelects_12_io_ins_7),
    .io_ins_8(StickySelects_12_io_ins_8),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5),
    .io_outs_6(StickySelects_12_io_outs_6),
    .io_outs_7(StickySelects_12_io_outs_7),
    .io_outs_8(StickySelects_12_io_outs_8)
  );
  StickySelects_1 StickySelects_13 ( // @[MemPrimitives.scala 124:33:@22219.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_ins_6(StickySelects_13_io_ins_6),
    .io_ins_7(StickySelects_13_io_ins_7),
    .io_ins_8(StickySelects_13_io_ins_8),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5),
    .io_outs_6(StickySelects_13_io_outs_6),
    .io_outs_7(StickySelects_13_io_outs_7),
    .io_outs_8(StickySelects_13_io_outs_8)
  );
  StickySelects_1 StickySelects_14 ( // @[MemPrimitives.scala 124:33:@22308.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_ins_6(StickySelects_14_io_ins_6),
    .io_ins_7(StickySelects_14_io_ins_7),
    .io_ins_8(StickySelects_14_io_ins_8),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5),
    .io_outs_6(StickySelects_14_io_outs_6),
    .io_outs_7(StickySelects_14_io_outs_7),
    .io_outs_8(StickySelects_14_io_outs_8)
  );
  StickySelects_1 StickySelects_15 ( // @[MemPrimitives.scala 124:33:@22397.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_ins_6(StickySelects_15_io_ins_6),
    .io_ins_7(StickySelects_15_io_ins_7),
    .io_ins_8(StickySelects_15_io_ins_8),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5),
    .io_outs_6(StickySelects_15_io_outs_6),
    .io_outs_7(StickySelects_15_io_outs_7),
    .io_outs_8(StickySelects_15_io_outs_8)
  );
  StickySelects_1 StickySelects_16 ( // @[MemPrimitives.scala 124:33:@22486.4]
    .clock(StickySelects_16_clock),
    .reset(StickySelects_16_reset),
    .io_ins_0(StickySelects_16_io_ins_0),
    .io_ins_1(StickySelects_16_io_ins_1),
    .io_ins_2(StickySelects_16_io_ins_2),
    .io_ins_3(StickySelects_16_io_ins_3),
    .io_ins_4(StickySelects_16_io_ins_4),
    .io_ins_5(StickySelects_16_io_ins_5),
    .io_ins_6(StickySelects_16_io_ins_6),
    .io_ins_7(StickySelects_16_io_ins_7),
    .io_ins_8(StickySelects_16_io_ins_8),
    .io_outs_0(StickySelects_16_io_outs_0),
    .io_outs_1(StickySelects_16_io_outs_1),
    .io_outs_2(StickySelects_16_io_outs_2),
    .io_outs_3(StickySelects_16_io_outs_3),
    .io_outs_4(StickySelects_16_io_outs_4),
    .io_outs_5(StickySelects_16_io_outs_5),
    .io_outs_6(StickySelects_16_io_outs_6),
    .io_outs_7(StickySelects_16_io_outs_7),
    .io_outs_8(StickySelects_16_io_outs_8)
  );
  StickySelects_1 StickySelects_17 ( // @[MemPrimitives.scala 124:33:@22575.4]
    .clock(StickySelects_17_clock),
    .reset(StickySelects_17_reset),
    .io_ins_0(StickySelects_17_io_ins_0),
    .io_ins_1(StickySelects_17_io_ins_1),
    .io_ins_2(StickySelects_17_io_ins_2),
    .io_ins_3(StickySelects_17_io_ins_3),
    .io_ins_4(StickySelects_17_io_ins_4),
    .io_ins_5(StickySelects_17_io_ins_5),
    .io_ins_6(StickySelects_17_io_ins_6),
    .io_ins_7(StickySelects_17_io_ins_7),
    .io_ins_8(StickySelects_17_io_ins_8),
    .io_outs_0(StickySelects_17_io_outs_0),
    .io_outs_1(StickySelects_17_io_outs_1),
    .io_outs_2(StickySelects_17_io_outs_2),
    .io_outs_3(StickySelects_17_io_outs_3),
    .io_outs_4(StickySelects_17_io_outs_4),
    .io_outs_5(StickySelects_17_io_outs_5),
    .io_outs_6(StickySelects_17_io_outs_6),
    .io_outs_7(StickySelects_17_io_outs_7),
    .io_outs_8(StickySelects_17_io_outs_8)
  );
  StickySelects_1 StickySelects_18 ( // @[MemPrimitives.scala 124:33:@22664.4]
    .clock(StickySelects_18_clock),
    .reset(StickySelects_18_reset),
    .io_ins_0(StickySelects_18_io_ins_0),
    .io_ins_1(StickySelects_18_io_ins_1),
    .io_ins_2(StickySelects_18_io_ins_2),
    .io_ins_3(StickySelects_18_io_ins_3),
    .io_ins_4(StickySelects_18_io_ins_4),
    .io_ins_5(StickySelects_18_io_ins_5),
    .io_ins_6(StickySelects_18_io_ins_6),
    .io_ins_7(StickySelects_18_io_ins_7),
    .io_ins_8(StickySelects_18_io_ins_8),
    .io_outs_0(StickySelects_18_io_outs_0),
    .io_outs_1(StickySelects_18_io_outs_1),
    .io_outs_2(StickySelects_18_io_outs_2),
    .io_outs_3(StickySelects_18_io_outs_3),
    .io_outs_4(StickySelects_18_io_outs_4),
    .io_outs_5(StickySelects_18_io_outs_5),
    .io_outs_6(StickySelects_18_io_outs_6),
    .io_outs_7(StickySelects_18_io_outs_7),
    .io_outs_8(StickySelects_18_io_outs_8)
  );
  StickySelects_1 StickySelects_19 ( // @[MemPrimitives.scala 124:33:@22753.4]
    .clock(StickySelects_19_clock),
    .reset(StickySelects_19_reset),
    .io_ins_0(StickySelects_19_io_ins_0),
    .io_ins_1(StickySelects_19_io_ins_1),
    .io_ins_2(StickySelects_19_io_ins_2),
    .io_ins_3(StickySelects_19_io_ins_3),
    .io_ins_4(StickySelects_19_io_ins_4),
    .io_ins_5(StickySelects_19_io_ins_5),
    .io_ins_6(StickySelects_19_io_ins_6),
    .io_ins_7(StickySelects_19_io_ins_7),
    .io_ins_8(StickySelects_19_io_ins_8),
    .io_outs_0(StickySelects_19_io_outs_0),
    .io_outs_1(StickySelects_19_io_outs_1),
    .io_outs_2(StickySelects_19_io_outs_2),
    .io_outs_3(StickySelects_19_io_outs_3),
    .io_outs_4(StickySelects_19_io_outs_4),
    .io_outs_5(StickySelects_19_io_outs_5),
    .io_outs_6(StickySelects_19_io_outs_6),
    .io_outs_7(StickySelects_19_io_outs_7),
    .io_outs_8(StickySelects_19_io_outs_8)
  );
  StickySelects_1 StickySelects_20 ( // @[MemPrimitives.scala 124:33:@22842.4]
    .clock(StickySelects_20_clock),
    .reset(StickySelects_20_reset),
    .io_ins_0(StickySelects_20_io_ins_0),
    .io_ins_1(StickySelects_20_io_ins_1),
    .io_ins_2(StickySelects_20_io_ins_2),
    .io_ins_3(StickySelects_20_io_ins_3),
    .io_ins_4(StickySelects_20_io_ins_4),
    .io_ins_5(StickySelects_20_io_ins_5),
    .io_ins_6(StickySelects_20_io_ins_6),
    .io_ins_7(StickySelects_20_io_ins_7),
    .io_ins_8(StickySelects_20_io_ins_8),
    .io_outs_0(StickySelects_20_io_outs_0),
    .io_outs_1(StickySelects_20_io_outs_1),
    .io_outs_2(StickySelects_20_io_outs_2),
    .io_outs_3(StickySelects_20_io_outs_3),
    .io_outs_4(StickySelects_20_io_outs_4),
    .io_outs_5(StickySelects_20_io_outs_5),
    .io_outs_6(StickySelects_20_io_outs_6),
    .io_outs_7(StickySelects_20_io_outs_7),
    .io_outs_8(StickySelects_20_io_outs_8)
  );
  StickySelects_1 StickySelects_21 ( // @[MemPrimitives.scala 124:33:@22931.4]
    .clock(StickySelects_21_clock),
    .reset(StickySelects_21_reset),
    .io_ins_0(StickySelects_21_io_ins_0),
    .io_ins_1(StickySelects_21_io_ins_1),
    .io_ins_2(StickySelects_21_io_ins_2),
    .io_ins_3(StickySelects_21_io_ins_3),
    .io_ins_4(StickySelects_21_io_ins_4),
    .io_ins_5(StickySelects_21_io_ins_5),
    .io_ins_6(StickySelects_21_io_ins_6),
    .io_ins_7(StickySelects_21_io_ins_7),
    .io_ins_8(StickySelects_21_io_ins_8),
    .io_outs_0(StickySelects_21_io_outs_0),
    .io_outs_1(StickySelects_21_io_outs_1),
    .io_outs_2(StickySelects_21_io_outs_2),
    .io_outs_3(StickySelects_21_io_outs_3),
    .io_outs_4(StickySelects_21_io_outs_4),
    .io_outs_5(StickySelects_21_io_outs_5),
    .io_outs_6(StickySelects_21_io_outs_6),
    .io_outs_7(StickySelects_21_io_outs_7),
    .io_outs_8(StickySelects_21_io_outs_8)
  );
  StickySelects_1 StickySelects_22 ( // @[MemPrimitives.scala 124:33:@23020.4]
    .clock(StickySelects_22_clock),
    .reset(StickySelects_22_reset),
    .io_ins_0(StickySelects_22_io_ins_0),
    .io_ins_1(StickySelects_22_io_ins_1),
    .io_ins_2(StickySelects_22_io_ins_2),
    .io_ins_3(StickySelects_22_io_ins_3),
    .io_ins_4(StickySelects_22_io_ins_4),
    .io_ins_5(StickySelects_22_io_ins_5),
    .io_ins_6(StickySelects_22_io_ins_6),
    .io_ins_7(StickySelects_22_io_ins_7),
    .io_ins_8(StickySelects_22_io_ins_8),
    .io_outs_0(StickySelects_22_io_outs_0),
    .io_outs_1(StickySelects_22_io_outs_1),
    .io_outs_2(StickySelects_22_io_outs_2),
    .io_outs_3(StickySelects_22_io_outs_3),
    .io_outs_4(StickySelects_22_io_outs_4),
    .io_outs_5(StickySelects_22_io_outs_5),
    .io_outs_6(StickySelects_22_io_outs_6),
    .io_outs_7(StickySelects_22_io_outs_7),
    .io_outs_8(StickySelects_22_io_outs_8)
  );
  StickySelects_1 StickySelects_23 ( // @[MemPrimitives.scala 124:33:@23109.4]
    .clock(StickySelects_23_clock),
    .reset(StickySelects_23_reset),
    .io_ins_0(StickySelects_23_io_ins_0),
    .io_ins_1(StickySelects_23_io_ins_1),
    .io_ins_2(StickySelects_23_io_ins_2),
    .io_ins_3(StickySelects_23_io_ins_3),
    .io_ins_4(StickySelects_23_io_ins_4),
    .io_ins_5(StickySelects_23_io_ins_5),
    .io_ins_6(StickySelects_23_io_ins_6),
    .io_ins_7(StickySelects_23_io_ins_7),
    .io_ins_8(StickySelects_23_io_ins_8),
    .io_outs_0(StickySelects_23_io_outs_0),
    .io_outs_1(StickySelects_23_io_outs_1),
    .io_outs_2(StickySelects_23_io_outs_2),
    .io_outs_3(StickySelects_23_io_outs_3),
    .io_outs_4(StickySelects_23_io_outs_4),
    .io_outs_5(StickySelects_23_io_outs_5),
    .io_outs_6(StickySelects_23_io_outs_6),
    .io_outs_7(StickySelects_23_io_outs_7),
    .io_outs_8(StickySelects_23_io_outs_8)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@23199.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@23207.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@23215.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@23223.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@23231.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@23239.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@23247.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@23255.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@23263.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@23271.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@23279.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@23287.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@23343.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@23351.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@23359.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@23367.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@23375.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@23383.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@23391.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@23399.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@23407.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@23415.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@23423.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@23431.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@23487.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@23495.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@23503.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@23511.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@23519.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@23527.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@23535.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@23543.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@23551.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@23559.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@23567.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@23575.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@23631.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@23639.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@23647.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@23655.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@23663.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@23671.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@23679.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@23687.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@23695.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@23703.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@23711.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@23719.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@23775.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@23783.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@23791.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@23799.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@23807.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@23815.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@23823.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@23831.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@23839.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@23847.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@23855.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@23863.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@23919.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@23927.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@23935.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@23943.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@23951.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@23959.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@23967.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@23975.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@23983.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@23991.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@23999.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@24007.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@24063.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@24071.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@24079.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@24087.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@24095.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@24103.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@24111.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@24119.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@24127.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@24135.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@24143.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@24151.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@24207.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@24215.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@24223.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@24231.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@24239.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@24247.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@24255.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@24263.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@24271.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@24279.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@24287.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@24295.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_96 ( // @[package.scala 93:22:@24351.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_97 ( // @[package.scala 93:22:@24359.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_98 ( // @[package.scala 93:22:@24367.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_99 ( // @[package.scala 93:22:@24375.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_100 ( // @[package.scala 93:22:@24383.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_101 ( // @[package.scala 93:22:@24391.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_102 ( // @[package.scala 93:22:@24399.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_103 ( // @[package.scala 93:22:@24407.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_104 ( // @[package.scala 93:22:@24415.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_105 ( // @[package.scala 93:22:@24423.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_106 ( // @[package.scala 93:22:@24431.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_107 ( // @[package.scala 93:22:@24439.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_108 ( // @[package.scala 93:22:@24495.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_109 ( // @[package.scala 93:22:@24503.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_110 ( // @[package.scala 93:22:@24511.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_111 ( // @[package.scala 93:22:@24519.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_112 ( // @[package.scala 93:22:@24527.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_113 ( // @[package.scala 93:22:@24535.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_114 ( // @[package.scala 93:22:@24543.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_115 ( // @[package.scala 93:22:@24551.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_116 ( // @[package.scala 93:22:@24559.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_117 ( // @[package.scala 93:22:@24567.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_118 ( // @[package.scala 93:22:@24575.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_119 ( // @[package.scala 93:22:@24583.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_120 ( // @[package.scala 93:22:@24639.4]
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_121 ( // @[package.scala 93:22:@24647.4]
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_122 ( // @[package.scala 93:22:@24655.4]
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_123 ( // @[package.scala 93:22:@24663.4]
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_124 ( // @[package.scala 93:22:@24671.4]
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_125 ( // @[package.scala 93:22:@24679.4]
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_126 ( // @[package.scala 93:22:@24687.4]
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_127 ( // @[package.scala 93:22:@24695.4]
    .clock(RetimeWrapper_127_clock),
    .reset(RetimeWrapper_127_reset),
    .io_flow(RetimeWrapper_127_io_flow),
    .io_in(RetimeWrapper_127_io_in),
    .io_out(RetimeWrapper_127_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_128 ( // @[package.scala 93:22:@24703.4]
    .clock(RetimeWrapper_128_clock),
    .reset(RetimeWrapper_128_reset),
    .io_flow(RetimeWrapper_128_io_flow),
    .io_in(RetimeWrapper_128_io_in),
    .io_out(RetimeWrapper_128_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_129 ( // @[package.scala 93:22:@24711.4]
    .clock(RetimeWrapper_129_clock),
    .reset(RetimeWrapper_129_reset),
    .io_flow(RetimeWrapper_129_io_flow),
    .io_in(RetimeWrapper_129_io_in),
    .io_out(RetimeWrapper_129_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_130 ( // @[package.scala 93:22:@24719.4]
    .clock(RetimeWrapper_130_clock),
    .reset(RetimeWrapper_130_reset),
    .io_flow(RetimeWrapper_130_io_flow),
    .io_in(RetimeWrapper_130_io_in),
    .io_out(RetimeWrapper_130_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_131 ( // @[package.scala 93:22:@24727.4]
    .clock(RetimeWrapper_131_clock),
    .reset(RetimeWrapper_131_reset),
    .io_flow(RetimeWrapper_131_io_flow),
    .io_in(RetimeWrapper_131_io_in),
    .io_out(RetimeWrapper_131_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_132 ( // @[package.scala 93:22:@24783.4]
    .clock(RetimeWrapper_132_clock),
    .reset(RetimeWrapper_132_reset),
    .io_flow(RetimeWrapper_132_io_flow),
    .io_in(RetimeWrapper_132_io_in),
    .io_out(RetimeWrapper_132_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_133 ( // @[package.scala 93:22:@24791.4]
    .clock(RetimeWrapper_133_clock),
    .reset(RetimeWrapper_133_reset),
    .io_flow(RetimeWrapper_133_io_flow),
    .io_in(RetimeWrapper_133_io_in),
    .io_out(RetimeWrapper_133_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_134 ( // @[package.scala 93:22:@24799.4]
    .clock(RetimeWrapper_134_clock),
    .reset(RetimeWrapper_134_reset),
    .io_flow(RetimeWrapper_134_io_flow),
    .io_in(RetimeWrapper_134_io_in),
    .io_out(RetimeWrapper_134_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_135 ( // @[package.scala 93:22:@24807.4]
    .clock(RetimeWrapper_135_clock),
    .reset(RetimeWrapper_135_reset),
    .io_flow(RetimeWrapper_135_io_flow),
    .io_in(RetimeWrapper_135_io_in),
    .io_out(RetimeWrapper_135_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_136 ( // @[package.scala 93:22:@24815.4]
    .clock(RetimeWrapper_136_clock),
    .reset(RetimeWrapper_136_reset),
    .io_flow(RetimeWrapper_136_io_flow),
    .io_in(RetimeWrapper_136_io_in),
    .io_out(RetimeWrapper_136_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_137 ( // @[package.scala 93:22:@24823.4]
    .clock(RetimeWrapper_137_clock),
    .reset(RetimeWrapper_137_reset),
    .io_flow(RetimeWrapper_137_io_flow),
    .io_in(RetimeWrapper_137_io_in),
    .io_out(RetimeWrapper_137_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_138 ( // @[package.scala 93:22:@24831.4]
    .clock(RetimeWrapper_138_clock),
    .reset(RetimeWrapper_138_reset),
    .io_flow(RetimeWrapper_138_io_flow),
    .io_in(RetimeWrapper_138_io_in),
    .io_out(RetimeWrapper_138_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_139 ( // @[package.scala 93:22:@24839.4]
    .clock(RetimeWrapper_139_clock),
    .reset(RetimeWrapper_139_reset),
    .io_flow(RetimeWrapper_139_io_flow),
    .io_in(RetimeWrapper_139_io_in),
    .io_out(RetimeWrapper_139_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_140 ( // @[package.scala 93:22:@24847.4]
    .clock(RetimeWrapper_140_clock),
    .reset(RetimeWrapper_140_reset),
    .io_flow(RetimeWrapper_140_io_flow),
    .io_in(RetimeWrapper_140_io_in),
    .io_out(RetimeWrapper_140_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_141 ( // @[package.scala 93:22:@24855.4]
    .clock(RetimeWrapper_141_clock),
    .reset(RetimeWrapper_141_reset),
    .io_flow(RetimeWrapper_141_io_flow),
    .io_in(RetimeWrapper_141_io_in),
    .io_out(RetimeWrapper_141_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_142 ( // @[package.scala 93:22:@24863.4]
    .clock(RetimeWrapper_142_clock),
    .reset(RetimeWrapper_142_reset),
    .io_flow(RetimeWrapper_142_io_flow),
    .io_in(RetimeWrapper_142_io_in),
    .io_out(RetimeWrapper_142_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_143 ( // @[package.scala 93:22:@24871.4]
    .clock(RetimeWrapper_143_clock),
    .reset(RetimeWrapper_143_reset),
    .io_flow(RetimeWrapper_143_io_flow),
    .io_in(RetimeWrapper_143_io_in),
    .io_out(RetimeWrapper_143_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_144 ( // @[package.scala 93:22:@24927.4]
    .clock(RetimeWrapper_144_clock),
    .reset(RetimeWrapper_144_reset),
    .io_flow(RetimeWrapper_144_io_flow),
    .io_in(RetimeWrapper_144_io_in),
    .io_out(RetimeWrapper_144_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_145 ( // @[package.scala 93:22:@24935.4]
    .clock(RetimeWrapper_145_clock),
    .reset(RetimeWrapper_145_reset),
    .io_flow(RetimeWrapper_145_io_flow),
    .io_in(RetimeWrapper_145_io_in),
    .io_out(RetimeWrapper_145_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_146 ( // @[package.scala 93:22:@24943.4]
    .clock(RetimeWrapper_146_clock),
    .reset(RetimeWrapper_146_reset),
    .io_flow(RetimeWrapper_146_io_flow),
    .io_in(RetimeWrapper_146_io_in),
    .io_out(RetimeWrapper_146_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_147 ( // @[package.scala 93:22:@24951.4]
    .clock(RetimeWrapper_147_clock),
    .reset(RetimeWrapper_147_reset),
    .io_flow(RetimeWrapper_147_io_flow),
    .io_in(RetimeWrapper_147_io_in),
    .io_out(RetimeWrapper_147_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_148 ( // @[package.scala 93:22:@24959.4]
    .clock(RetimeWrapper_148_clock),
    .reset(RetimeWrapper_148_reset),
    .io_flow(RetimeWrapper_148_io_flow),
    .io_in(RetimeWrapper_148_io_in),
    .io_out(RetimeWrapper_148_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_149 ( // @[package.scala 93:22:@24967.4]
    .clock(RetimeWrapper_149_clock),
    .reset(RetimeWrapper_149_reset),
    .io_flow(RetimeWrapper_149_io_flow),
    .io_in(RetimeWrapper_149_io_in),
    .io_out(RetimeWrapper_149_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_150 ( // @[package.scala 93:22:@24975.4]
    .clock(RetimeWrapper_150_clock),
    .reset(RetimeWrapper_150_reset),
    .io_flow(RetimeWrapper_150_io_flow),
    .io_in(RetimeWrapper_150_io_in),
    .io_out(RetimeWrapper_150_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_151 ( // @[package.scala 93:22:@24983.4]
    .clock(RetimeWrapper_151_clock),
    .reset(RetimeWrapper_151_reset),
    .io_flow(RetimeWrapper_151_io_flow),
    .io_in(RetimeWrapper_151_io_in),
    .io_out(RetimeWrapper_151_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_152 ( // @[package.scala 93:22:@24991.4]
    .clock(RetimeWrapper_152_clock),
    .reset(RetimeWrapper_152_reset),
    .io_flow(RetimeWrapper_152_io_flow),
    .io_in(RetimeWrapper_152_io_in),
    .io_out(RetimeWrapper_152_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_153 ( // @[package.scala 93:22:@24999.4]
    .clock(RetimeWrapper_153_clock),
    .reset(RetimeWrapper_153_reset),
    .io_flow(RetimeWrapper_153_io_flow),
    .io_in(RetimeWrapper_153_io_in),
    .io_out(RetimeWrapper_153_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_154 ( // @[package.scala 93:22:@25007.4]
    .clock(RetimeWrapper_154_clock),
    .reset(RetimeWrapper_154_reset),
    .io_flow(RetimeWrapper_154_io_flow),
    .io_in(RetimeWrapper_154_io_in),
    .io_out(RetimeWrapper_154_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_155 ( // @[package.scala 93:22:@25015.4]
    .clock(RetimeWrapper_155_clock),
    .reset(RetimeWrapper_155_reset),
    .io_flow(RetimeWrapper_155_io_flow),
    .io_in(RetimeWrapper_155_io_in),
    .io_out(RetimeWrapper_155_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_156 ( // @[package.scala 93:22:@25071.4]
    .clock(RetimeWrapper_156_clock),
    .reset(RetimeWrapper_156_reset),
    .io_flow(RetimeWrapper_156_io_flow),
    .io_in(RetimeWrapper_156_io_in),
    .io_out(RetimeWrapper_156_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_157 ( // @[package.scala 93:22:@25079.4]
    .clock(RetimeWrapper_157_clock),
    .reset(RetimeWrapper_157_reset),
    .io_flow(RetimeWrapper_157_io_flow),
    .io_in(RetimeWrapper_157_io_in),
    .io_out(RetimeWrapper_157_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_158 ( // @[package.scala 93:22:@25087.4]
    .clock(RetimeWrapper_158_clock),
    .reset(RetimeWrapper_158_reset),
    .io_flow(RetimeWrapper_158_io_flow),
    .io_in(RetimeWrapper_158_io_in),
    .io_out(RetimeWrapper_158_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_159 ( // @[package.scala 93:22:@25095.4]
    .clock(RetimeWrapper_159_clock),
    .reset(RetimeWrapper_159_reset),
    .io_flow(RetimeWrapper_159_io_flow),
    .io_in(RetimeWrapper_159_io_in),
    .io_out(RetimeWrapper_159_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_160 ( // @[package.scala 93:22:@25103.4]
    .clock(RetimeWrapper_160_clock),
    .reset(RetimeWrapper_160_reset),
    .io_flow(RetimeWrapper_160_io_flow),
    .io_in(RetimeWrapper_160_io_in),
    .io_out(RetimeWrapper_160_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_161 ( // @[package.scala 93:22:@25111.4]
    .clock(RetimeWrapper_161_clock),
    .reset(RetimeWrapper_161_reset),
    .io_flow(RetimeWrapper_161_io_flow),
    .io_in(RetimeWrapper_161_io_in),
    .io_out(RetimeWrapper_161_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_162 ( // @[package.scala 93:22:@25119.4]
    .clock(RetimeWrapper_162_clock),
    .reset(RetimeWrapper_162_reset),
    .io_flow(RetimeWrapper_162_io_flow),
    .io_in(RetimeWrapper_162_io_in),
    .io_out(RetimeWrapper_162_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_163 ( // @[package.scala 93:22:@25127.4]
    .clock(RetimeWrapper_163_clock),
    .reset(RetimeWrapper_163_reset),
    .io_flow(RetimeWrapper_163_io_flow),
    .io_in(RetimeWrapper_163_io_in),
    .io_out(RetimeWrapper_163_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_164 ( // @[package.scala 93:22:@25135.4]
    .clock(RetimeWrapper_164_clock),
    .reset(RetimeWrapper_164_reset),
    .io_flow(RetimeWrapper_164_io_flow),
    .io_in(RetimeWrapper_164_io_in),
    .io_out(RetimeWrapper_164_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_165 ( // @[package.scala 93:22:@25143.4]
    .clock(RetimeWrapper_165_clock),
    .reset(RetimeWrapper_165_reset),
    .io_flow(RetimeWrapper_165_io_flow),
    .io_in(RetimeWrapper_165_io_in),
    .io_out(RetimeWrapper_165_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_166 ( // @[package.scala 93:22:@25151.4]
    .clock(RetimeWrapper_166_clock),
    .reset(RetimeWrapper_166_reset),
    .io_flow(RetimeWrapper_166_io_flow),
    .io_in(RetimeWrapper_166_io_in),
    .io_out(RetimeWrapper_166_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_167 ( // @[package.scala 93:22:@25159.4]
    .clock(RetimeWrapper_167_clock),
    .reset(RetimeWrapper_167_reset),
    .io_flow(RetimeWrapper_167_io_flow),
    .io_in(RetimeWrapper_167_io_in),
    .io_out(RetimeWrapper_167_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_168 ( // @[package.scala 93:22:@25215.4]
    .clock(RetimeWrapper_168_clock),
    .reset(RetimeWrapper_168_reset),
    .io_flow(RetimeWrapper_168_io_flow),
    .io_in(RetimeWrapper_168_io_in),
    .io_out(RetimeWrapper_168_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_169 ( // @[package.scala 93:22:@25223.4]
    .clock(RetimeWrapper_169_clock),
    .reset(RetimeWrapper_169_reset),
    .io_flow(RetimeWrapper_169_io_flow),
    .io_in(RetimeWrapper_169_io_in),
    .io_out(RetimeWrapper_169_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_170 ( // @[package.scala 93:22:@25231.4]
    .clock(RetimeWrapper_170_clock),
    .reset(RetimeWrapper_170_reset),
    .io_flow(RetimeWrapper_170_io_flow),
    .io_in(RetimeWrapper_170_io_in),
    .io_out(RetimeWrapper_170_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_171 ( // @[package.scala 93:22:@25239.4]
    .clock(RetimeWrapper_171_clock),
    .reset(RetimeWrapper_171_reset),
    .io_flow(RetimeWrapper_171_io_flow),
    .io_in(RetimeWrapper_171_io_in),
    .io_out(RetimeWrapper_171_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_172 ( // @[package.scala 93:22:@25247.4]
    .clock(RetimeWrapper_172_clock),
    .reset(RetimeWrapper_172_reset),
    .io_flow(RetimeWrapper_172_io_flow),
    .io_in(RetimeWrapper_172_io_in),
    .io_out(RetimeWrapper_172_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_173 ( // @[package.scala 93:22:@25255.4]
    .clock(RetimeWrapper_173_clock),
    .reset(RetimeWrapper_173_reset),
    .io_flow(RetimeWrapper_173_io_flow),
    .io_in(RetimeWrapper_173_io_in),
    .io_out(RetimeWrapper_173_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_174 ( // @[package.scala 93:22:@25263.4]
    .clock(RetimeWrapper_174_clock),
    .reset(RetimeWrapper_174_reset),
    .io_flow(RetimeWrapper_174_io_flow),
    .io_in(RetimeWrapper_174_io_in),
    .io_out(RetimeWrapper_174_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_175 ( // @[package.scala 93:22:@25271.4]
    .clock(RetimeWrapper_175_clock),
    .reset(RetimeWrapper_175_reset),
    .io_flow(RetimeWrapper_175_io_flow),
    .io_in(RetimeWrapper_175_io_in),
    .io_out(RetimeWrapper_175_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_176 ( // @[package.scala 93:22:@25279.4]
    .clock(RetimeWrapper_176_clock),
    .reset(RetimeWrapper_176_reset),
    .io_flow(RetimeWrapper_176_io_flow),
    .io_in(RetimeWrapper_176_io_in),
    .io_out(RetimeWrapper_176_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_177 ( // @[package.scala 93:22:@25287.4]
    .clock(RetimeWrapper_177_clock),
    .reset(RetimeWrapper_177_reset),
    .io_flow(RetimeWrapper_177_io_flow),
    .io_in(RetimeWrapper_177_io_in),
    .io_out(RetimeWrapper_177_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_178 ( // @[package.scala 93:22:@25295.4]
    .clock(RetimeWrapper_178_clock),
    .reset(RetimeWrapper_178_reset),
    .io_flow(RetimeWrapper_178_io_flow),
    .io_in(RetimeWrapper_178_io_in),
    .io_out(RetimeWrapper_178_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_179 ( // @[package.scala 93:22:@25303.4]
    .clock(RetimeWrapper_179_clock),
    .reset(RetimeWrapper_179_reset),
    .io_flow(RetimeWrapper_179_io_flow),
    .io_in(RetimeWrapper_179_io_in),
    .io_out(RetimeWrapper_179_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_180 ( // @[package.scala 93:22:@25359.4]
    .clock(RetimeWrapper_180_clock),
    .reset(RetimeWrapper_180_reset),
    .io_flow(RetimeWrapper_180_io_flow),
    .io_in(RetimeWrapper_180_io_in),
    .io_out(RetimeWrapper_180_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_181 ( // @[package.scala 93:22:@25367.4]
    .clock(RetimeWrapper_181_clock),
    .reset(RetimeWrapper_181_reset),
    .io_flow(RetimeWrapper_181_io_flow),
    .io_in(RetimeWrapper_181_io_in),
    .io_out(RetimeWrapper_181_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_182 ( // @[package.scala 93:22:@25375.4]
    .clock(RetimeWrapper_182_clock),
    .reset(RetimeWrapper_182_reset),
    .io_flow(RetimeWrapper_182_io_flow),
    .io_in(RetimeWrapper_182_io_in),
    .io_out(RetimeWrapper_182_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_183 ( // @[package.scala 93:22:@25383.4]
    .clock(RetimeWrapper_183_clock),
    .reset(RetimeWrapper_183_reset),
    .io_flow(RetimeWrapper_183_io_flow),
    .io_in(RetimeWrapper_183_io_in),
    .io_out(RetimeWrapper_183_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_184 ( // @[package.scala 93:22:@25391.4]
    .clock(RetimeWrapper_184_clock),
    .reset(RetimeWrapper_184_reset),
    .io_flow(RetimeWrapper_184_io_flow),
    .io_in(RetimeWrapper_184_io_in),
    .io_out(RetimeWrapper_184_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_185 ( // @[package.scala 93:22:@25399.4]
    .clock(RetimeWrapper_185_clock),
    .reset(RetimeWrapper_185_reset),
    .io_flow(RetimeWrapper_185_io_flow),
    .io_in(RetimeWrapper_185_io_in),
    .io_out(RetimeWrapper_185_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_186 ( // @[package.scala 93:22:@25407.4]
    .clock(RetimeWrapper_186_clock),
    .reset(RetimeWrapper_186_reset),
    .io_flow(RetimeWrapper_186_io_flow),
    .io_in(RetimeWrapper_186_io_in),
    .io_out(RetimeWrapper_186_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_187 ( // @[package.scala 93:22:@25415.4]
    .clock(RetimeWrapper_187_clock),
    .reset(RetimeWrapper_187_reset),
    .io_flow(RetimeWrapper_187_io_flow),
    .io_in(RetimeWrapper_187_io_in),
    .io_out(RetimeWrapper_187_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_188 ( // @[package.scala 93:22:@25423.4]
    .clock(RetimeWrapper_188_clock),
    .reset(RetimeWrapper_188_reset),
    .io_flow(RetimeWrapper_188_io_flow),
    .io_in(RetimeWrapper_188_io_in),
    .io_out(RetimeWrapper_188_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_189 ( // @[package.scala 93:22:@25431.4]
    .clock(RetimeWrapper_189_clock),
    .reset(RetimeWrapper_189_reset),
    .io_flow(RetimeWrapper_189_io_flow),
    .io_in(RetimeWrapper_189_io_in),
    .io_out(RetimeWrapper_189_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_190 ( // @[package.scala 93:22:@25439.4]
    .clock(RetimeWrapper_190_clock),
    .reset(RetimeWrapper_190_reset),
    .io_flow(RetimeWrapper_190_io_flow),
    .io_in(RetimeWrapper_190_io_in),
    .io_out(RetimeWrapper_190_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_191 ( // @[package.scala 93:22:@25447.4]
    .clock(RetimeWrapper_191_clock),
    .reset(RetimeWrapper_191_reset),
    .io_flow(RetimeWrapper_191_io_flow),
    .io_in(RetimeWrapper_191_io_in),
    .io_out(RetimeWrapper_191_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_192 ( // @[package.scala 93:22:@25503.4]
    .clock(RetimeWrapper_192_clock),
    .reset(RetimeWrapper_192_reset),
    .io_flow(RetimeWrapper_192_io_flow),
    .io_in(RetimeWrapper_192_io_in),
    .io_out(RetimeWrapper_192_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_193 ( // @[package.scala 93:22:@25511.4]
    .clock(RetimeWrapper_193_clock),
    .reset(RetimeWrapper_193_reset),
    .io_flow(RetimeWrapper_193_io_flow),
    .io_in(RetimeWrapper_193_io_in),
    .io_out(RetimeWrapper_193_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_194 ( // @[package.scala 93:22:@25519.4]
    .clock(RetimeWrapper_194_clock),
    .reset(RetimeWrapper_194_reset),
    .io_flow(RetimeWrapper_194_io_flow),
    .io_in(RetimeWrapper_194_io_in),
    .io_out(RetimeWrapper_194_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_195 ( // @[package.scala 93:22:@25527.4]
    .clock(RetimeWrapper_195_clock),
    .reset(RetimeWrapper_195_reset),
    .io_flow(RetimeWrapper_195_io_flow),
    .io_in(RetimeWrapper_195_io_in),
    .io_out(RetimeWrapper_195_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_196 ( // @[package.scala 93:22:@25535.4]
    .clock(RetimeWrapper_196_clock),
    .reset(RetimeWrapper_196_reset),
    .io_flow(RetimeWrapper_196_io_flow),
    .io_in(RetimeWrapper_196_io_in),
    .io_out(RetimeWrapper_196_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_197 ( // @[package.scala 93:22:@25543.4]
    .clock(RetimeWrapper_197_clock),
    .reset(RetimeWrapper_197_reset),
    .io_flow(RetimeWrapper_197_io_flow),
    .io_in(RetimeWrapper_197_io_in),
    .io_out(RetimeWrapper_197_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_198 ( // @[package.scala 93:22:@25551.4]
    .clock(RetimeWrapper_198_clock),
    .reset(RetimeWrapper_198_reset),
    .io_flow(RetimeWrapper_198_io_flow),
    .io_in(RetimeWrapper_198_io_in),
    .io_out(RetimeWrapper_198_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_199 ( // @[package.scala 93:22:@25559.4]
    .clock(RetimeWrapper_199_clock),
    .reset(RetimeWrapper_199_reset),
    .io_flow(RetimeWrapper_199_io_flow),
    .io_in(RetimeWrapper_199_io_in),
    .io_out(RetimeWrapper_199_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_200 ( // @[package.scala 93:22:@25567.4]
    .clock(RetimeWrapper_200_clock),
    .reset(RetimeWrapper_200_reset),
    .io_flow(RetimeWrapper_200_io_flow),
    .io_in(RetimeWrapper_200_io_in),
    .io_out(RetimeWrapper_200_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_201 ( // @[package.scala 93:22:@25575.4]
    .clock(RetimeWrapper_201_clock),
    .reset(RetimeWrapper_201_reset),
    .io_flow(RetimeWrapper_201_io_flow),
    .io_in(RetimeWrapper_201_io_in),
    .io_out(RetimeWrapper_201_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_202 ( // @[package.scala 93:22:@25583.4]
    .clock(RetimeWrapper_202_clock),
    .reset(RetimeWrapper_202_reset),
    .io_flow(RetimeWrapper_202_io_flow),
    .io_in(RetimeWrapper_202_io_in),
    .io_out(RetimeWrapper_202_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_203 ( // @[package.scala 93:22:@25591.4]
    .clock(RetimeWrapper_203_clock),
    .reset(RetimeWrapper_203_reset),
    .io_flow(RetimeWrapper_203_io_flow),
    .io_in(RetimeWrapper_203_io_in),
    .io_out(RetimeWrapper_203_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_204 ( // @[package.scala 93:22:@25647.4]
    .clock(RetimeWrapper_204_clock),
    .reset(RetimeWrapper_204_reset),
    .io_flow(RetimeWrapper_204_io_flow),
    .io_in(RetimeWrapper_204_io_in),
    .io_out(RetimeWrapper_204_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_205 ( // @[package.scala 93:22:@25655.4]
    .clock(RetimeWrapper_205_clock),
    .reset(RetimeWrapper_205_reset),
    .io_flow(RetimeWrapper_205_io_flow),
    .io_in(RetimeWrapper_205_io_in),
    .io_out(RetimeWrapper_205_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_206 ( // @[package.scala 93:22:@25663.4]
    .clock(RetimeWrapper_206_clock),
    .reset(RetimeWrapper_206_reset),
    .io_flow(RetimeWrapper_206_io_flow),
    .io_in(RetimeWrapper_206_io_in),
    .io_out(RetimeWrapper_206_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_207 ( // @[package.scala 93:22:@25671.4]
    .clock(RetimeWrapper_207_clock),
    .reset(RetimeWrapper_207_reset),
    .io_flow(RetimeWrapper_207_io_flow),
    .io_in(RetimeWrapper_207_io_in),
    .io_out(RetimeWrapper_207_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_208 ( // @[package.scala 93:22:@25679.4]
    .clock(RetimeWrapper_208_clock),
    .reset(RetimeWrapper_208_reset),
    .io_flow(RetimeWrapper_208_io_flow),
    .io_in(RetimeWrapper_208_io_in),
    .io_out(RetimeWrapper_208_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_209 ( // @[package.scala 93:22:@25687.4]
    .clock(RetimeWrapper_209_clock),
    .reset(RetimeWrapper_209_reset),
    .io_flow(RetimeWrapper_209_io_flow),
    .io_in(RetimeWrapper_209_io_in),
    .io_out(RetimeWrapper_209_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_210 ( // @[package.scala 93:22:@25695.4]
    .clock(RetimeWrapper_210_clock),
    .reset(RetimeWrapper_210_reset),
    .io_flow(RetimeWrapper_210_io_flow),
    .io_in(RetimeWrapper_210_io_in),
    .io_out(RetimeWrapper_210_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_211 ( // @[package.scala 93:22:@25703.4]
    .clock(RetimeWrapper_211_clock),
    .reset(RetimeWrapper_211_reset),
    .io_flow(RetimeWrapper_211_io_flow),
    .io_in(RetimeWrapper_211_io_in),
    .io_out(RetimeWrapper_211_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_212 ( // @[package.scala 93:22:@25711.4]
    .clock(RetimeWrapper_212_clock),
    .reset(RetimeWrapper_212_reset),
    .io_flow(RetimeWrapper_212_io_flow),
    .io_in(RetimeWrapper_212_io_in),
    .io_out(RetimeWrapper_212_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_213 ( // @[package.scala 93:22:@25719.4]
    .clock(RetimeWrapper_213_clock),
    .reset(RetimeWrapper_213_reset),
    .io_flow(RetimeWrapper_213_io_flow),
    .io_in(RetimeWrapper_213_io_in),
    .io_out(RetimeWrapper_213_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_214 ( // @[package.scala 93:22:@25727.4]
    .clock(RetimeWrapper_214_clock),
    .reset(RetimeWrapper_214_reset),
    .io_flow(RetimeWrapper_214_io_flow),
    .io_in(RetimeWrapper_214_io_in),
    .io_out(RetimeWrapper_214_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_215 ( // @[package.scala 93:22:@25735.4]
    .clock(RetimeWrapper_215_clock),
    .reset(RetimeWrapper_215_reset),
    .io_flow(RetimeWrapper_215_io_flow),
    .io_in(RetimeWrapper_215_io_in),
    .io_out(RetimeWrapper_215_io_out)
  );
  assign _T_700 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@20570.4]
  assign _T_702 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@20571.4]
  assign _T_703 = _T_700 & _T_702; // @[MemPrimitives.scala 82:228:@20572.4]
  assign _T_704 = io_wPort_0_en_0 & _T_703; // @[MemPrimitives.scala 83:102:@20573.4]
  assign _T_706 = io_wPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@20574.4]
  assign _T_708 = io_wPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@20575.4]
  assign _T_709 = _T_706 & _T_708; // @[MemPrimitives.scala 82:228:@20576.4]
  assign _T_710 = io_wPort_2_en_0 & _T_709; // @[MemPrimitives.scala 83:102:@20577.4]
  assign _T_712 = {_T_704,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20579.4]
  assign _T_714 = {_T_710,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20581.4]
  assign _T_715 = _T_704 ? _T_712 : _T_714; // @[Mux.scala 31:69:@20582.4]
  assign _T_720 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@20589.4]
  assign _T_722 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@20590.4]
  assign _T_723 = _T_720 & _T_722; // @[MemPrimitives.scala 82:228:@20591.4]
  assign _T_724 = io_wPort_1_en_0 & _T_723; // @[MemPrimitives.scala 83:102:@20592.4]
  assign _T_726 = io_wPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@20593.4]
  assign _T_728 = io_wPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@20594.4]
  assign _T_729 = _T_726 & _T_728; // @[MemPrimitives.scala 82:228:@20595.4]
  assign _T_730 = io_wPort_3_en_0 & _T_729; // @[MemPrimitives.scala 83:102:@20596.4]
  assign _T_732 = {_T_724,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20598.4]
  assign _T_734 = {_T_730,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20600.4]
  assign _T_735 = _T_724 ? _T_732 : _T_734; // @[Mux.scala 31:69:@20601.4]
  assign _T_742 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@20609.4]
  assign _T_743 = _T_700 & _T_742; // @[MemPrimitives.scala 82:228:@20610.4]
  assign _T_744 = io_wPort_0_en_0 & _T_743; // @[MemPrimitives.scala 83:102:@20611.4]
  assign _T_748 = io_wPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@20613.4]
  assign _T_749 = _T_706 & _T_748; // @[MemPrimitives.scala 82:228:@20614.4]
  assign _T_750 = io_wPort_2_en_0 & _T_749; // @[MemPrimitives.scala 83:102:@20615.4]
  assign _T_752 = {_T_744,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20617.4]
  assign _T_754 = {_T_750,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20619.4]
  assign _T_755 = _T_744 ? _T_752 : _T_754; // @[Mux.scala 31:69:@20620.4]
  assign _T_762 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@20628.4]
  assign _T_763 = _T_720 & _T_762; // @[MemPrimitives.scala 82:228:@20629.4]
  assign _T_764 = io_wPort_1_en_0 & _T_763; // @[MemPrimitives.scala 83:102:@20630.4]
  assign _T_768 = io_wPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@20632.4]
  assign _T_769 = _T_726 & _T_768; // @[MemPrimitives.scala 82:228:@20633.4]
  assign _T_770 = io_wPort_3_en_0 & _T_769; // @[MemPrimitives.scala 83:102:@20634.4]
  assign _T_772 = {_T_764,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20636.4]
  assign _T_774 = {_T_770,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20638.4]
  assign _T_775 = _T_764 ? _T_772 : _T_774; // @[Mux.scala 31:69:@20639.4]
  assign _T_782 = io_wPort_0_banks_1 == 3'h4; // @[MemPrimitives.scala 82:210:@20647.4]
  assign _T_783 = _T_700 & _T_782; // @[MemPrimitives.scala 82:228:@20648.4]
  assign _T_784 = io_wPort_0_en_0 & _T_783; // @[MemPrimitives.scala 83:102:@20649.4]
  assign _T_788 = io_wPort_2_banks_1 == 3'h4; // @[MemPrimitives.scala 82:210:@20651.4]
  assign _T_789 = _T_706 & _T_788; // @[MemPrimitives.scala 82:228:@20652.4]
  assign _T_790 = io_wPort_2_en_0 & _T_789; // @[MemPrimitives.scala 83:102:@20653.4]
  assign _T_792 = {_T_784,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20655.4]
  assign _T_794 = {_T_790,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20657.4]
  assign _T_795 = _T_784 ? _T_792 : _T_794; // @[Mux.scala 31:69:@20658.4]
  assign _T_802 = io_wPort_1_banks_1 == 3'h5; // @[MemPrimitives.scala 82:210:@20666.4]
  assign _T_803 = _T_720 & _T_802; // @[MemPrimitives.scala 82:228:@20667.4]
  assign _T_804 = io_wPort_1_en_0 & _T_803; // @[MemPrimitives.scala 83:102:@20668.4]
  assign _T_808 = io_wPort_3_banks_1 == 3'h5; // @[MemPrimitives.scala 82:210:@20670.4]
  assign _T_809 = _T_726 & _T_808; // @[MemPrimitives.scala 82:228:@20671.4]
  assign _T_810 = io_wPort_3_en_0 & _T_809; // @[MemPrimitives.scala 83:102:@20672.4]
  assign _T_812 = {_T_804,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20674.4]
  assign _T_814 = {_T_810,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20676.4]
  assign _T_815 = _T_804 ? _T_812 : _T_814; // @[Mux.scala 31:69:@20677.4]
  assign _T_820 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@20684.4]
  assign _T_823 = _T_820 & _T_702; // @[MemPrimitives.scala 82:228:@20686.4]
  assign _T_824 = io_wPort_0_en_0 & _T_823; // @[MemPrimitives.scala 83:102:@20687.4]
  assign _T_826 = io_wPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@20688.4]
  assign _T_829 = _T_826 & _T_708; // @[MemPrimitives.scala 82:228:@20690.4]
  assign _T_830 = io_wPort_2_en_0 & _T_829; // @[MemPrimitives.scala 83:102:@20691.4]
  assign _T_832 = {_T_824,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20693.4]
  assign _T_834 = {_T_830,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20695.4]
  assign _T_835 = _T_824 ? _T_832 : _T_834; // @[Mux.scala 31:69:@20696.4]
  assign _T_840 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@20703.4]
  assign _T_843 = _T_840 & _T_722; // @[MemPrimitives.scala 82:228:@20705.4]
  assign _T_844 = io_wPort_1_en_0 & _T_843; // @[MemPrimitives.scala 83:102:@20706.4]
  assign _T_846 = io_wPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@20707.4]
  assign _T_849 = _T_846 & _T_728; // @[MemPrimitives.scala 82:228:@20709.4]
  assign _T_850 = io_wPort_3_en_0 & _T_849; // @[MemPrimitives.scala 83:102:@20710.4]
  assign _T_852 = {_T_844,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20712.4]
  assign _T_854 = {_T_850,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20714.4]
  assign _T_855 = _T_844 ? _T_852 : _T_854; // @[Mux.scala 31:69:@20715.4]
  assign _T_863 = _T_820 & _T_742; // @[MemPrimitives.scala 82:228:@20724.4]
  assign _T_864 = io_wPort_0_en_0 & _T_863; // @[MemPrimitives.scala 83:102:@20725.4]
  assign _T_869 = _T_826 & _T_748; // @[MemPrimitives.scala 82:228:@20728.4]
  assign _T_870 = io_wPort_2_en_0 & _T_869; // @[MemPrimitives.scala 83:102:@20729.4]
  assign _T_872 = {_T_864,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20731.4]
  assign _T_874 = {_T_870,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20733.4]
  assign _T_875 = _T_864 ? _T_872 : _T_874; // @[Mux.scala 31:69:@20734.4]
  assign _T_883 = _T_840 & _T_762; // @[MemPrimitives.scala 82:228:@20743.4]
  assign _T_884 = io_wPort_1_en_0 & _T_883; // @[MemPrimitives.scala 83:102:@20744.4]
  assign _T_889 = _T_846 & _T_768; // @[MemPrimitives.scala 82:228:@20747.4]
  assign _T_890 = io_wPort_3_en_0 & _T_889; // @[MemPrimitives.scala 83:102:@20748.4]
  assign _T_892 = {_T_884,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20750.4]
  assign _T_894 = {_T_890,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20752.4]
  assign _T_895 = _T_884 ? _T_892 : _T_894; // @[Mux.scala 31:69:@20753.4]
  assign _T_903 = _T_820 & _T_782; // @[MemPrimitives.scala 82:228:@20762.4]
  assign _T_904 = io_wPort_0_en_0 & _T_903; // @[MemPrimitives.scala 83:102:@20763.4]
  assign _T_909 = _T_826 & _T_788; // @[MemPrimitives.scala 82:228:@20766.4]
  assign _T_910 = io_wPort_2_en_0 & _T_909; // @[MemPrimitives.scala 83:102:@20767.4]
  assign _T_912 = {_T_904,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20769.4]
  assign _T_914 = {_T_910,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20771.4]
  assign _T_915 = _T_904 ? _T_912 : _T_914; // @[Mux.scala 31:69:@20772.4]
  assign _T_923 = _T_840 & _T_802; // @[MemPrimitives.scala 82:228:@20781.4]
  assign _T_924 = io_wPort_1_en_0 & _T_923; // @[MemPrimitives.scala 83:102:@20782.4]
  assign _T_929 = _T_846 & _T_808; // @[MemPrimitives.scala 82:228:@20785.4]
  assign _T_930 = io_wPort_3_en_0 & _T_929; // @[MemPrimitives.scala 83:102:@20786.4]
  assign _T_932 = {_T_924,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20788.4]
  assign _T_934 = {_T_930,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20790.4]
  assign _T_935 = _T_924 ? _T_932 : _T_934; // @[Mux.scala 31:69:@20791.4]
  assign _T_940 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20798.4]
  assign _T_943 = _T_940 & _T_702; // @[MemPrimitives.scala 82:228:@20800.4]
  assign _T_944 = io_wPort_0_en_0 & _T_943; // @[MemPrimitives.scala 83:102:@20801.4]
  assign _T_946 = io_wPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20802.4]
  assign _T_949 = _T_946 & _T_708; // @[MemPrimitives.scala 82:228:@20804.4]
  assign _T_950 = io_wPort_2_en_0 & _T_949; // @[MemPrimitives.scala 83:102:@20805.4]
  assign _T_952 = {_T_944,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20807.4]
  assign _T_954 = {_T_950,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20809.4]
  assign _T_955 = _T_944 ? _T_952 : _T_954; // @[Mux.scala 31:69:@20810.4]
  assign _T_960 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20817.4]
  assign _T_963 = _T_960 & _T_722; // @[MemPrimitives.scala 82:228:@20819.4]
  assign _T_964 = io_wPort_1_en_0 & _T_963; // @[MemPrimitives.scala 83:102:@20820.4]
  assign _T_966 = io_wPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20821.4]
  assign _T_969 = _T_966 & _T_728; // @[MemPrimitives.scala 82:228:@20823.4]
  assign _T_970 = io_wPort_3_en_0 & _T_969; // @[MemPrimitives.scala 83:102:@20824.4]
  assign _T_972 = {_T_964,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20826.4]
  assign _T_974 = {_T_970,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20828.4]
  assign _T_975 = _T_964 ? _T_972 : _T_974; // @[Mux.scala 31:69:@20829.4]
  assign _T_983 = _T_940 & _T_742; // @[MemPrimitives.scala 82:228:@20838.4]
  assign _T_984 = io_wPort_0_en_0 & _T_983; // @[MemPrimitives.scala 83:102:@20839.4]
  assign _T_989 = _T_946 & _T_748; // @[MemPrimitives.scala 82:228:@20842.4]
  assign _T_990 = io_wPort_2_en_0 & _T_989; // @[MemPrimitives.scala 83:102:@20843.4]
  assign _T_992 = {_T_984,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20845.4]
  assign _T_994 = {_T_990,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20847.4]
  assign _T_995 = _T_984 ? _T_992 : _T_994; // @[Mux.scala 31:69:@20848.4]
  assign _T_1003 = _T_960 & _T_762; // @[MemPrimitives.scala 82:228:@20857.4]
  assign _T_1004 = io_wPort_1_en_0 & _T_1003; // @[MemPrimitives.scala 83:102:@20858.4]
  assign _T_1009 = _T_966 & _T_768; // @[MemPrimitives.scala 82:228:@20861.4]
  assign _T_1010 = io_wPort_3_en_0 & _T_1009; // @[MemPrimitives.scala 83:102:@20862.4]
  assign _T_1012 = {_T_1004,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20864.4]
  assign _T_1014 = {_T_1010,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20866.4]
  assign _T_1015 = _T_1004 ? _T_1012 : _T_1014; // @[Mux.scala 31:69:@20867.4]
  assign _T_1023 = _T_940 & _T_782; // @[MemPrimitives.scala 82:228:@20876.4]
  assign _T_1024 = io_wPort_0_en_0 & _T_1023; // @[MemPrimitives.scala 83:102:@20877.4]
  assign _T_1029 = _T_946 & _T_788; // @[MemPrimitives.scala 82:228:@20880.4]
  assign _T_1030 = io_wPort_2_en_0 & _T_1029; // @[MemPrimitives.scala 83:102:@20881.4]
  assign _T_1032 = {_T_1024,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20883.4]
  assign _T_1034 = {_T_1030,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20885.4]
  assign _T_1035 = _T_1024 ? _T_1032 : _T_1034; // @[Mux.scala 31:69:@20886.4]
  assign _T_1043 = _T_960 & _T_802; // @[MemPrimitives.scala 82:228:@20895.4]
  assign _T_1044 = io_wPort_1_en_0 & _T_1043; // @[MemPrimitives.scala 83:102:@20896.4]
  assign _T_1049 = _T_966 & _T_808; // @[MemPrimitives.scala 82:228:@20899.4]
  assign _T_1050 = io_wPort_3_en_0 & _T_1049; // @[MemPrimitives.scala 83:102:@20900.4]
  assign _T_1052 = {_T_1044,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20902.4]
  assign _T_1054 = {_T_1050,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20904.4]
  assign _T_1055 = _T_1044 ? _T_1052 : _T_1054; // @[Mux.scala 31:69:@20905.4]
  assign _T_1060 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20912.4]
  assign _T_1063 = _T_1060 & _T_702; // @[MemPrimitives.scala 82:228:@20914.4]
  assign _T_1064 = io_wPort_0_en_0 & _T_1063; // @[MemPrimitives.scala 83:102:@20915.4]
  assign _T_1066 = io_wPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20916.4]
  assign _T_1069 = _T_1066 & _T_708; // @[MemPrimitives.scala 82:228:@20918.4]
  assign _T_1070 = io_wPort_2_en_0 & _T_1069; // @[MemPrimitives.scala 83:102:@20919.4]
  assign _T_1072 = {_T_1064,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20921.4]
  assign _T_1074 = {_T_1070,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20923.4]
  assign _T_1075 = _T_1064 ? _T_1072 : _T_1074; // @[Mux.scala 31:69:@20924.4]
  assign _T_1080 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20931.4]
  assign _T_1083 = _T_1080 & _T_722; // @[MemPrimitives.scala 82:228:@20933.4]
  assign _T_1084 = io_wPort_1_en_0 & _T_1083; // @[MemPrimitives.scala 83:102:@20934.4]
  assign _T_1086 = io_wPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20935.4]
  assign _T_1089 = _T_1086 & _T_728; // @[MemPrimitives.scala 82:228:@20937.4]
  assign _T_1090 = io_wPort_3_en_0 & _T_1089; // @[MemPrimitives.scala 83:102:@20938.4]
  assign _T_1092 = {_T_1084,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20940.4]
  assign _T_1094 = {_T_1090,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20942.4]
  assign _T_1095 = _T_1084 ? _T_1092 : _T_1094; // @[Mux.scala 31:69:@20943.4]
  assign _T_1103 = _T_1060 & _T_742; // @[MemPrimitives.scala 82:228:@20952.4]
  assign _T_1104 = io_wPort_0_en_0 & _T_1103; // @[MemPrimitives.scala 83:102:@20953.4]
  assign _T_1109 = _T_1066 & _T_748; // @[MemPrimitives.scala 82:228:@20956.4]
  assign _T_1110 = io_wPort_2_en_0 & _T_1109; // @[MemPrimitives.scala 83:102:@20957.4]
  assign _T_1112 = {_T_1104,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20959.4]
  assign _T_1114 = {_T_1110,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20961.4]
  assign _T_1115 = _T_1104 ? _T_1112 : _T_1114; // @[Mux.scala 31:69:@20962.4]
  assign _T_1123 = _T_1080 & _T_762; // @[MemPrimitives.scala 82:228:@20971.4]
  assign _T_1124 = io_wPort_1_en_0 & _T_1123; // @[MemPrimitives.scala 83:102:@20972.4]
  assign _T_1129 = _T_1086 & _T_768; // @[MemPrimitives.scala 82:228:@20975.4]
  assign _T_1130 = io_wPort_3_en_0 & _T_1129; // @[MemPrimitives.scala 83:102:@20976.4]
  assign _T_1132 = {_T_1124,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20978.4]
  assign _T_1134 = {_T_1130,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20980.4]
  assign _T_1135 = _T_1124 ? _T_1132 : _T_1134; // @[Mux.scala 31:69:@20981.4]
  assign _T_1143 = _T_1060 & _T_782; // @[MemPrimitives.scala 82:228:@20990.4]
  assign _T_1144 = io_wPort_0_en_0 & _T_1143; // @[MemPrimitives.scala 83:102:@20991.4]
  assign _T_1149 = _T_1066 & _T_788; // @[MemPrimitives.scala 82:228:@20994.4]
  assign _T_1150 = io_wPort_2_en_0 & _T_1149; // @[MemPrimitives.scala 83:102:@20995.4]
  assign _T_1152 = {_T_1144,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20997.4]
  assign _T_1154 = {_T_1150,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20999.4]
  assign _T_1155 = _T_1144 ? _T_1152 : _T_1154; // @[Mux.scala 31:69:@21000.4]
  assign _T_1163 = _T_1080 & _T_802; // @[MemPrimitives.scala 82:228:@21009.4]
  assign _T_1164 = io_wPort_1_en_0 & _T_1163; // @[MemPrimitives.scala 83:102:@21010.4]
  assign _T_1169 = _T_1086 & _T_808; // @[MemPrimitives.scala 82:228:@21013.4]
  assign _T_1170 = io_wPort_3_en_0 & _T_1169; // @[MemPrimitives.scala 83:102:@21014.4]
  assign _T_1172 = {_T_1164,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@21016.4]
  assign _T_1174 = {_T_1170,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@21018.4]
  assign _T_1175 = _T_1164 ? _T_1172 : _T_1174; // @[Mux.scala 31:69:@21019.4]
  assign _T_1180 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21026.4]
  assign _T_1182 = io_rPort_1_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21027.4]
  assign _T_1183 = _T_1180 & _T_1182; // @[MemPrimitives.scala 110:228:@21028.4]
  assign _T_1186 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21030.4]
  assign _T_1188 = io_rPort_3_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21031.4]
  assign _T_1189 = _T_1186 & _T_1188; // @[MemPrimitives.scala 110:228:@21032.4]
  assign _T_1192 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21034.4]
  assign _T_1194 = io_rPort_6_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21035.4]
  assign _T_1195 = _T_1192 & _T_1194; // @[MemPrimitives.scala 110:228:@21036.4]
  assign _T_1198 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21038.4]
  assign _T_1200 = io_rPort_8_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21039.4]
  assign _T_1201 = _T_1198 & _T_1200; // @[MemPrimitives.scala 110:228:@21040.4]
  assign _T_1204 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21042.4]
  assign _T_1206 = io_rPort_10_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21043.4]
  assign _T_1207 = _T_1204 & _T_1206; // @[MemPrimitives.scala 110:228:@21044.4]
  assign _T_1210 = io_rPort_12_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21046.4]
  assign _T_1212 = io_rPort_12_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21047.4]
  assign _T_1213 = _T_1210 & _T_1212; // @[MemPrimitives.scala 110:228:@21048.4]
  assign _T_1216 = io_rPort_15_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21050.4]
  assign _T_1218 = io_rPort_15_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21051.4]
  assign _T_1219 = _T_1216 & _T_1218; // @[MemPrimitives.scala 110:228:@21052.4]
  assign _T_1222 = io_rPort_16_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21054.4]
  assign _T_1224 = io_rPort_16_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21055.4]
  assign _T_1225 = _T_1222 & _T_1224; // @[MemPrimitives.scala 110:228:@21056.4]
  assign _T_1228 = io_rPort_17_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21058.4]
  assign _T_1230 = io_rPort_17_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@21059.4]
  assign _T_1231 = _T_1228 & _T_1230; // @[MemPrimitives.scala 110:228:@21060.4]
  assign _T_1233 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@21074.4]
  assign _T_1234 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@21075.4]
  assign _T_1235 = StickySelects_io_outs_2; // @[MemPrimitives.scala 126:35:@21076.4]
  assign _T_1236 = StickySelects_io_outs_3; // @[MemPrimitives.scala 126:35:@21077.4]
  assign _T_1237 = StickySelects_io_outs_4; // @[MemPrimitives.scala 126:35:@21078.4]
  assign _T_1238 = StickySelects_io_outs_5; // @[MemPrimitives.scala 126:35:@21079.4]
  assign _T_1239 = StickySelects_io_outs_6; // @[MemPrimitives.scala 126:35:@21080.4]
  assign _T_1240 = StickySelects_io_outs_7; // @[MemPrimitives.scala 126:35:@21081.4]
  assign _T_1241 = StickySelects_io_outs_8; // @[MemPrimitives.scala 126:35:@21082.4]
  assign _T_1243 = {_T_1233,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21084.4]
  assign _T_1245 = {_T_1234,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21086.4]
  assign _T_1247 = {_T_1235,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21088.4]
  assign _T_1249 = {_T_1236,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21090.4]
  assign _T_1251 = {_T_1237,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21092.4]
  assign _T_1253 = {_T_1238,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21094.4]
  assign _T_1255 = {_T_1239,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21096.4]
  assign _T_1257 = {_T_1240,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21098.4]
  assign _T_1259 = {_T_1241,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21100.4]
  assign _T_1260 = _T_1240 ? _T_1257 : _T_1259; // @[Mux.scala 31:69:@21101.4]
  assign _T_1261 = _T_1239 ? _T_1255 : _T_1260; // @[Mux.scala 31:69:@21102.4]
  assign _T_1262 = _T_1238 ? _T_1253 : _T_1261; // @[Mux.scala 31:69:@21103.4]
  assign _T_1263 = _T_1237 ? _T_1251 : _T_1262; // @[Mux.scala 31:69:@21104.4]
  assign _T_1264 = _T_1236 ? _T_1249 : _T_1263; // @[Mux.scala 31:69:@21105.4]
  assign _T_1265 = _T_1235 ? _T_1247 : _T_1264; // @[Mux.scala 31:69:@21106.4]
  assign _T_1266 = _T_1234 ? _T_1245 : _T_1265; // @[Mux.scala 31:69:@21107.4]
  assign _T_1267 = _T_1233 ? _T_1243 : _T_1266; // @[Mux.scala 31:69:@21108.4]
  assign _T_1272 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21115.4]
  assign _T_1274 = io_rPort_0_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21116.4]
  assign _T_1275 = _T_1272 & _T_1274; // @[MemPrimitives.scala 110:228:@21117.4]
  assign _T_1278 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21119.4]
  assign _T_1280 = io_rPort_2_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21120.4]
  assign _T_1281 = _T_1278 & _T_1280; // @[MemPrimitives.scala 110:228:@21121.4]
  assign _T_1284 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21123.4]
  assign _T_1286 = io_rPort_4_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21124.4]
  assign _T_1287 = _T_1284 & _T_1286; // @[MemPrimitives.scala 110:228:@21125.4]
  assign _T_1290 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21127.4]
  assign _T_1292 = io_rPort_5_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21128.4]
  assign _T_1293 = _T_1290 & _T_1292; // @[MemPrimitives.scala 110:228:@21129.4]
  assign _T_1296 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21131.4]
  assign _T_1298 = io_rPort_7_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21132.4]
  assign _T_1299 = _T_1296 & _T_1298; // @[MemPrimitives.scala 110:228:@21133.4]
  assign _T_1302 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21135.4]
  assign _T_1304 = io_rPort_9_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21136.4]
  assign _T_1305 = _T_1302 & _T_1304; // @[MemPrimitives.scala 110:228:@21137.4]
  assign _T_1308 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21139.4]
  assign _T_1310 = io_rPort_11_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21140.4]
  assign _T_1311 = _T_1308 & _T_1310; // @[MemPrimitives.scala 110:228:@21141.4]
  assign _T_1314 = io_rPort_13_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21143.4]
  assign _T_1316 = io_rPort_13_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21144.4]
  assign _T_1317 = _T_1314 & _T_1316; // @[MemPrimitives.scala 110:228:@21145.4]
  assign _T_1320 = io_rPort_14_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@21147.4]
  assign _T_1322 = io_rPort_14_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@21148.4]
  assign _T_1323 = _T_1320 & _T_1322; // @[MemPrimitives.scala 110:228:@21149.4]
  assign _T_1325 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@21163.4]
  assign _T_1326 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@21164.4]
  assign _T_1327 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@21165.4]
  assign _T_1328 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@21166.4]
  assign _T_1329 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 126:35:@21167.4]
  assign _T_1330 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 126:35:@21168.4]
  assign _T_1331 = StickySelects_1_io_outs_6; // @[MemPrimitives.scala 126:35:@21169.4]
  assign _T_1332 = StickySelects_1_io_outs_7; // @[MemPrimitives.scala 126:35:@21170.4]
  assign _T_1333 = StickySelects_1_io_outs_8; // @[MemPrimitives.scala 126:35:@21171.4]
  assign _T_1335 = {_T_1325,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21173.4]
  assign _T_1337 = {_T_1326,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21175.4]
  assign _T_1339 = {_T_1327,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21177.4]
  assign _T_1341 = {_T_1328,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21179.4]
  assign _T_1343 = {_T_1329,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21181.4]
  assign _T_1345 = {_T_1330,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21183.4]
  assign _T_1347 = {_T_1331,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21185.4]
  assign _T_1349 = {_T_1332,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21187.4]
  assign _T_1351 = {_T_1333,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21189.4]
  assign _T_1352 = _T_1332 ? _T_1349 : _T_1351; // @[Mux.scala 31:69:@21190.4]
  assign _T_1353 = _T_1331 ? _T_1347 : _T_1352; // @[Mux.scala 31:69:@21191.4]
  assign _T_1354 = _T_1330 ? _T_1345 : _T_1353; // @[Mux.scala 31:69:@21192.4]
  assign _T_1355 = _T_1329 ? _T_1343 : _T_1354; // @[Mux.scala 31:69:@21193.4]
  assign _T_1356 = _T_1328 ? _T_1341 : _T_1355; // @[Mux.scala 31:69:@21194.4]
  assign _T_1357 = _T_1327 ? _T_1339 : _T_1356; // @[Mux.scala 31:69:@21195.4]
  assign _T_1358 = _T_1326 ? _T_1337 : _T_1357; // @[Mux.scala 31:69:@21196.4]
  assign _T_1359 = _T_1325 ? _T_1335 : _T_1358; // @[Mux.scala 31:69:@21197.4]
  assign _T_1366 = io_rPort_1_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21205.4]
  assign _T_1367 = _T_1180 & _T_1366; // @[MemPrimitives.scala 110:228:@21206.4]
  assign _T_1372 = io_rPort_3_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21209.4]
  assign _T_1373 = _T_1186 & _T_1372; // @[MemPrimitives.scala 110:228:@21210.4]
  assign _T_1378 = io_rPort_6_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21213.4]
  assign _T_1379 = _T_1192 & _T_1378; // @[MemPrimitives.scala 110:228:@21214.4]
  assign _T_1384 = io_rPort_8_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21217.4]
  assign _T_1385 = _T_1198 & _T_1384; // @[MemPrimitives.scala 110:228:@21218.4]
  assign _T_1390 = io_rPort_10_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21221.4]
  assign _T_1391 = _T_1204 & _T_1390; // @[MemPrimitives.scala 110:228:@21222.4]
  assign _T_1396 = io_rPort_12_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21225.4]
  assign _T_1397 = _T_1210 & _T_1396; // @[MemPrimitives.scala 110:228:@21226.4]
  assign _T_1402 = io_rPort_15_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21229.4]
  assign _T_1403 = _T_1216 & _T_1402; // @[MemPrimitives.scala 110:228:@21230.4]
  assign _T_1408 = io_rPort_16_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21233.4]
  assign _T_1409 = _T_1222 & _T_1408; // @[MemPrimitives.scala 110:228:@21234.4]
  assign _T_1414 = io_rPort_17_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@21237.4]
  assign _T_1415 = _T_1228 & _T_1414; // @[MemPrimitives.scala 110:228:@21238.4]
  assign _T_1417 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@21252.4]
  assign _T_1418 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@21253.4]
  assign _T_1419 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 126:35:@21254.4]
  assign _T_1420 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 126:35:@21255.4]
  assign _T_1421 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 126:35:@21256.4]
  assign _T_1422 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 126:35:@21257.4]
  assign _T_1423 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 126:35:@21258.4]
  assign _T_1424 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 126:35:@21259.4]
  assign _T_1425 = StickySelects_2_io_outs_8; // @[MemPrimitives.scala 126:35:@21260.4]
  assign _T_1427 = {_T_1417,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21262.4]
  assign _T_1429 = {_T_1418,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21264.4]
  assign _T_1431 = {_T_1419,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21266.4]
  assign _T_1433 = {_T_1420,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21268.4]
  assign _T_1435 = {_T_1421,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21270.4]
  assign _T_1437 = {_T_1422,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21272.4]
  assign _T_1439 = {_T_1423,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21274.4]
  assign _T_1441 = {_T_1424,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21276.4]
  assign _T_1443 = {_T_1425,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21278.4]
  assign _T_1444 = _T_1424 ? _T_1441 : _T_1443; // @[Mux.scala 31:69:@21279.4]
  assign _T_1445 = _T_1423 ? _T_1439 : _T_1444; // @[Mux.scala 31:69:@21280.4]
  assign _T_1446 = _T_1422 ? _T_1437 : _T_1445; // @[Mux.scala 31:69:@21281.4]
  assign _T_1447 = _T_1421 ? _T_1435 : _T_1446; // @[Mux.scala 31:69:@21282.4]
  assign _T_1448 = _T_1420 ? _T_1433 : _T_1447; // @[Mux.scala 31:69:@21283.4]
  assign _T_1449 = _T_1419 ? _T_1431 : _T_1448; // @[Mux.scala 31:69:@21284.4]
  assign _T_1450 = _T_1418 ? _T_1429 : _T_1449; // @[Mux.scala 31:69:@21285.4]
  assign _T_1451 = _T_1417 ? _T_1427 : _T_1450; // @[Mux.scala 31:69:@21286.4]
  assign _T_1458 = io_rPort_0_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21294.4]
  assign _T_1459 = _T_1272 & _T_1458; // @[MemPrimitives.scala 110:228:@21295.4]
  assign _T_1464 = io_rPort_2_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21298.4]
  assign _T_1465 = _T_1278 & _T_1464; // @[MemPrimitives.scala 110:228:@21299.4]
  assign _T_1470 = io_rPort_4_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21302.4]
  assign _T_1471 = _T_1284 & _T_1470; // @[MemPrimitives.scala 110:228:@21303.4]
  assign _T_1476 = io_rPort_5_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21306.4]
  assign _T_1477 = _T_1290 & _T_1476; // @[MemPrimitives.scala 110:228:@21307.4]
  assign _T_1482 = io_rPort_7_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21310.4]
  assign _T_1483 = _T_1296 & _T_1482; // @[MemPrimitives.scala 110:228:@21311.4]
  assign _T_1488 = io_rPort_9_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21314.4]
  assign _T_1489 = _T_1302 & _T_1488; // @[MemPrimitives.scala 110:228:@21315.4]
  assign _T_1494 = io_rPort_11_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21318.4]
  assign _T_1495 = _T_1308 & _T_1494; // @[MemPrimitives.scala 110:228:@21319.4]
  assign _T_1500 = io_rPort_13_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21322.4]
  assign _T_1501 = _T_1314 & _T_1500; // @[MemPrimitives.scala 110:228:@21323.4]
  assign _T_1506 = io_rPort_14_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@21326.4]
  assign _T_1507 = _T_1320 & _T_1506; // @[MemPrimitives.scala 110:228:@21327.4]
  assign _T_1509 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@21341.4]
  assign _T_1510 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@21342.4]
  assign _T_1511 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@21343.4]
  assign _T_1512 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@21344.4]
  assign _T_1513 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 126:35:@21345.4]
  assign _T_1514 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 126:35:@21346.4]
  assign _T_1515 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 126:35:@21347.4]
  assign _T_1516 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 126:35:@21348.4]
  assign _T_1517 = StickySelects_3_io_outs_8; // @[MemPrimitives.scala 126:35:@21349.4]
  assign _T_1519 = {_T_1509,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21351.4]
  assign _T_1521 = {_T_1510,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21353.4]
  assign _T_1523 = {_T_1511,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21355.4]
  assign _T_1525 = {_T_1512,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21357.4]
  assign _T_1527 = {_T_1513,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21359.4]
  assign _T_1529 = {_T_1514,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21361.4]
  assign _T_1531 = {_T_1515,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21363.4]
  assign _T_1533 = {_T_1516,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21365.4]
  assign _T_1535 = {_T_1517,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21367.4]
  assign _T_1536 = _T_1516 ? _T_1533 : _T_1535; // @[Mux.scala 31:69:@21368.4]
  assign _T_1537 = _T_1515 ? _T_1531 : _T_1536; // @[Mux.scala 31:69:@21369.4]
  assign _T_1538 = _T_1514 ? _T_1529 : _T_1537; // @[Mux.scala 31:69:@21370.4]
  assign _T_1539 = _T_1513 ? _T_1527 : _T_1538; // @[Mux.scala 31:69:@21371.4]
  assign _T_1540 = _T_1512 ? _T_1525 : _T_1539; // @[Mux.scala 31:69:@21372.4]
  assign _T_1541 = _T_1511 ? _T_1523 : _T_1540; // @[Mux.scala 31:69:@21373.4]
  assign _T_1542 = _T_1510 ? _T_1521 : _T_1541; // @[Mux.scala 31:69:@21374.4]
  assign _T_1543 = _T_1509 ? _T_1519 : _T_1542; // @[Mux.scala 31:69:@21375.4]
  assign _T_1550 = io_rPort_1_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21383.4]
  assign _T_1551 = _T_1180 & _T_1550; // @[MemPrimitives.scala 110:228:@21384.4]
  assign _T_1556 = io_rPort_3_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21387.4]
  assign _T_1557 = _T_1186 & _T_1556; // @[MemPrimitives.scala 110:228:@21388.4]
  assign _T_1562 = io_rPort_6_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21391.4]
  assign _T_1563 = _T_1192 & _T_1562; // @[MemPrimitives.scala 110:228:@21392.4]
  assign _T_1568 = io_rPort_8_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21395.4]
  assign _T_1569 = _T_1198 & _T_1568; // @[MemPrimitives.scala 110:228:@21396.4]
  assign _T_1574 = io_rPort_10_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21399.4]
  assign _T_1575 = _T_1204 & _T_1574; // @[MemPrimitives.scala 110:228:@21400.4]
  assign _T_1580 = io_rPort_12_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21403.4]
  assign _T_1581 = _T_1210 & _T_1580; // @[MemPrimitives.scala 110:228:@21404.4]
  assign _T_1586 = io_rPort_15_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21407.4]
  assign _T_1587 = _T_1216 & _T_1586; // @[MemPrimitives.scala 110:228:@21408.4]
  assign _T_1592 = io_rPort_16_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21411.4]
  assign _T_1593 = _T_1222 & _T_1592; // @[MemPrimitives.scala 110:228:@21412.4]
  assign _T_1598 = io_rPort_17_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@21415.4]
  assign _T_1599 = _T_1228 & _T_1598; // @[MemPrimitives.scala 110:228:@21416.4]
  assign _T_1601 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@21430.4]
  assign _T_1602 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@21431.4]
  assign _T_1603 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 126:35:@21432.4]
  assign _T_1604 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 126:35:@21433.4]
  assign _T_1605 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 126:35:@21434.4]
  assign _T_1606 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 126:35:@21435.4]
  assign _T_1607 = StickySelects_4_io_outs_6; // @[MemPrimitives.scala 126:35:@21436.4]
  assign _T_1608 = StickySelects_4_io_outs_7; // @[MemPrimitives.scala 126:35:@21437.4]
  assign _T_1609 = StickySelects_4_io_outs_8; // @[MemPrimitives.scala 126:35:@21438.4]
  assign _T_1611 = {_T_1601,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21440.4]
  assign _T_1613 = {_T_1602,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21442.4]
  assign _T_1615 = {_T_1603,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21444.4]
  assign _T_1617 = {_T_1604,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21446.4]
  assign _T_1619 = {_T_1605,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21448.4]
  assign _T_1621 = {_T_1606,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21450.4]
  assign _T_1623 = {_T_1607,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21452.4]
  assign _T_1625 = {_T_1608,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21454.4]
  assign _T_1627 = {_T_1609,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21456.4]
  assign _T_1628 = _T_1608 ? _T_1625 : _T_1627; // @[Mux.scala 31:69:@21457.4]
  assign _T_1629 = _T_1607 ? _T_1623 : _T_1628; // @[Mux.scala 31:69:@21458.4]
  assign _T_1630 = _T_1606 ? _T_1621 : _T_1629; // @[Mux.scala 31:69:@21459.4]
  assign _T_1631 = _T_1605 ? _T_1619 : _T_1630; // @[Mux.scala 31:69:@21460.4]
  assign _T_1632 = _T_1604 ? _T_1617 : _T_1631; // @[Mux.scala 31:69:@21461.4]
  assign _T_1633 = _T_1603 ? _T_1615 : _T_1632; // @[Mux.scala 31:69:@21462.4]
  assign _T_1634 = _T_1602 ? _T_1613 : _T_1633; // @[Mux.scala 31:69:@21463.4]
  assign _T_1635 = _T_1601 ? _T_1611 : _T_1634; // @[Mux.scala 31:69:@21464.4]
  assign _T_1642 = io_rPort_0_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21472.4]
  assign _T_1643 = _T_1272 & _T_1642; // @[MemPrimitives.scala 110:228:@21473.4]
  assign _T_1648 = io_rPort_2_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21476.4]
  assign _T_1649 = _T_1278 & _T_1648; // @[MemPrimitives.scala 110:228:@21477.4]
  assign _T_1654 = io_rPort_4_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21480.4]
  assign _T_1655 = _T_1284 & _T_1654; // @[MemPrimitives.scala 110:228:@21481.4]
  assign _T_1660 = io_rPort_5_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21484.4]
  assign _T_1661 = _T_1290 & _T_1660; // @[MemPrimitives.scala 110:228:@21485.4]
  assign _T_1666 = io_rPort_7_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21488.4]
  assign _T_1667 = _T_1296 & _T_1666; // @[MemPrimitives.scala 110:228:@21489.4]
  assign _T_1672 = io_rPort_9_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21492.4]
  assign _T_1673 = _T_1302 & _T_1672; // @[MemPrimitives.scala 110:228:@21493.4]
  assign _T_1678 = io_rPort_11_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21496.4]
  assign _T_1679 = _T_1308 & _T_1678; // @[MemPrimitives.scala 110:228:@21497.4]
  assign _T_1684 = io_rPort_13_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21500.4]
  assign _T_1685 = _T_1314 & _T_1684; // @[MemPrimitives.scala 110:228:@21501.4]
  assign _T_1690 = io_rPort_14_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@21504.4]
  assign _T_1691 = _T_1320 & _T_1690; // @[MemPrimitives.scala 110:228:@21505.4]
  assign _T_1693 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@21519.4]
  assign _T_1694 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@21520.4]
  assign _T_1695 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@21521.4]
  assign _T_1696 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@21522.4]
  assign _T_1697 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 126:35:@21523.4]
  assign _T_1698 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 126:35:@21524.4]
  assign _T_1699 = StickySelects_5_io_outs_6; // @[MemPrimitives.scala 126:35:@21525.4]
  assign _T_1700 = StickySelects_5_io_outs_7; // @[MemPrimitives.scala 126:35:@21526.4]
  assign _T_1701 = StickySelects_5_io_outs_8; // @[MemPrimitives.scala 126:35:@21527.4]
  assign _T_1703 = {_T_1693,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21529.4]
  assign _T_1705 = {_T_1694,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21531.4]
  assign _T_1707 = {_T_1695,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21533.4]
  assign _T_1709 = {_T_1696,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21535.4]
  assign _T_1711 = {_T_1697,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21537.4]
  assign _T_1713 = {_T_1698,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21539.4]
  assign _T_1715 = {_T_1699,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21541.4]
  assign _T_1717 = {_T_1700,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21543.4]
  assign _T_1719 = {_T_1701,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21545.4]
  assign _T_1720 = _T_1700 ? _T_1717 : _T_1719; // @[Mux.scala 31:69:@21546.4]
  assign _T_1721 = _T_1699 ? _T_1715 : _T_1720; // @[Mux.scala 31:69:@21547.4]
  assign _T_1722 = _T_1698 ? _T_1713 : _T_1721; // @[Mux.scala 31:69:@21548.4]
  assign _T_1723 = _T_1697 ? _T_1711 : _T_1722; // @[Mux.scala 31:69:@21549.4]
  assign _T_1724 = _T_1696 ? _T_1709 : _T_1723; // @[Mux.scala 31:69:@21550.4]
  assign _T_1725 = _T_1695 ? _T_1707 : _T_1724; // @[Mux.scala 31:69:@21551.4]
  assign _T_1726 = _T_1694 ? _T_1705 : _T_1725; // @[Mux.scala 31:69:@21552.4]
  assign _T_1727 = _T_1693 ? _T_1703 : _T_1726; // @[Mux.scala 31:69:@21553.4]
  assign _T_1732 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21560.4]
  assign _T_1735 = _T_1732 & _T_1182; // @[MemPrimitives.scala 110:228:@21562.4]
  assign _T_1738 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21564.4]
  assign _T_1741 = _T_1738 & _T_1188; // @[MemPrimitives.scala 110:228:@21566.4]
  assign _T_1744 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21568.4]
  assign _T_1747 = _T_1744 & _T_1194; // @[MemPrimitives.scala 110:228:@21570.4]
  assign _T_1750 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21572.4]
  assign _T_1753 = _T_1750 & _T_1200; // @[MemPrimitives.scala 110:228:@21574.4]
  assign _T_1756 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21576.4]
  assign _T_1759 = _T_1756 & _T_1206; // @[MemPrimitives.scala 110:228:@21578.4]
  assign _T_1762 = io_rPort_12_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21580.4]
  assign _T_1765 = _T_1762 & _T_1212; // @[MemPrimitives.scala 110:228:@21582.4]
  assign _T_1768 = io_rPort_15_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21584.4]
  assign _T_1771 = _T_1768 & _T_1218; // @[MemPrimitives.scala 110:228:@21586.4]
  assign _T_1774 = io_rPort_16_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21588.4]
  assign _T_1777 = _T_1774 & _T_1224; // @[MemPrimitives.scala 110:228:@21590.4]
  assign _T_1780 = io_rPort_17_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21592.4]
  assign _T_1783 = _T_1780 & _T_1230; // @[MemPrimitives.scala 110:228:@21594.4]
  assign _T_1785 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@21608.4]
  assign _T_1786 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@21609.4]
  assign _T_1787 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 126:35:@21610.4]
  assign _T_1788 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 126:35:@21611.4]
  assign _T_1789 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 126:35:@21612.4]
  assign _T_1790 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 126:35:@21613.4]
  assign _T_1791 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 126:35:@21614.4]
  assign _T_1792 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 126:35:@21615.4]
  assign _T_1793 = StickySelects_6_io_outs_8; // @[MemPrimitives.scala 126:35:@21616.4]
  assign _T_1795 = {_T_1785,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21618.4]
  assign _T_1797 = {_T_1786,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21620.4]
  assign _T_1799 = {_T_1787,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21622.4]
  assign _T_1801 = {_T_1788,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21624.4]
  assign _T_1803 = {_T_1789,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21626.4]
  assign _T_1805 = {_T_1790,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21628.4]
  assign _T_1807 = {_T_1791,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21630.4]
  assign _T_1809 = {_T_1792,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21632.4]
  assign _T_1811 = {_T_1793,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21634.4]
  assign _T_1812 = _T_1792 ? _T_1809 : _T_1811; // @[Mux.scala 31:69:@21635.4]
  assign _T_1813 = _T_1791 ? _T_1807 : _T_1812; // @[Mux.scala 31:69:@21636.4]
  assign _T_1814 = _T_1790 ? _T_1805 : _T_1813; // @[Mux.scala 31:69:@21637.4]
  assign _T_1815 = _T_1789 ? _T_1803 : _T_1814; // @[Mux.scala 31:69:@21638.4]
  assign _T_1816 = _T_1788 ? _T_1801 : _T_1815; // @[Mux.scala 31:69:@21639.4]
  assign _T_1817 = _T_1787 ? _T_1799 : _T_1816; // @[Mux.scala 31:69:@21640.4]
  assign _T_1818 = _T_1786 ? _T_1797 : _T_1817; // @[Mux.scala 31:69:@21641.4]
  assign _T_1819 = _T_1785 ? _T_1795 : _T_1818; // @[Mux.scala 31:69:@21642.4]
  assign _T_1824 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21649.4]
  assign _T_1827 = _T_1824 & _T_1274; // @[MemPrimitives.scala 110:228:@21651.4]
  assign _T_1830 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21653.4]
  assign _T_1833 = _T_1830 & _T_1280; // @[MemPrimitives.scala 110:228:@21655.4]
  assign _T_1836 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21657.4]
  assign _T_1839 = _T_1836 & _T_1286; // @[MemPrimitives.scala 110:228:@21659.4]
  assign _T_1842 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21661.4]
  assign _T_1845 = _T_1842 & _T_1292; // @[MemPrimitives.scala 110:228:@21663.4]
  assign _T_1848 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21665.4]
  assign _T_1851 = _T_1848 & _T_1298; // @[MemPrimitives.scala 110:228:@21667.4]
  assign _T_1854 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21669.4]
  assign _T_1857 = _T_1854 & _T_1304; // @[MemPrimitives.scala 110:228:@21671.4]
  assign _T_1860 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21673.4]
  assign _T_1863 = _T_1860 & _T_1310; // @[MemPrimitives.scala 110:228:@21675.4]
  assign _T_1866 = io_rPort_13_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21677.4]
  assign _T_1869 = _T_1866 & _T_1316; // @[MemPrimitives.scala 110:228:@21679.4]
  assign _T_1872 = io_rPort_14_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@21681.4]
  assign _T_1875 = _T_1872 & _T_1322; // @[MemPrimitives.scala 110:228:@21683.4]
  assign _T_1877 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@21697.4]
  assign _T_1878 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@21698.4]
  assign _T_1879 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@21699.4]
  assign _T_1880 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@21700.4]
  assign _T_1881 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 126:35:@21701.4]
  assign _T_1882 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 126:35:@21702.4]
  assign _T_1883 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 126:35:@21703.4]
  assign _T_1884 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 126:35:@21704.4]
  assign _T_1885 = StickySelects_7_io_outs_8; // @[MemPrimitives.scala 126:35:@21705.4]
  assign _T_1887 = {_T_1877,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21707.4]
  assign _T_1889 = {_T_1878,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21709.4]
  assign _T_1891 = {_T_1879,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21711.4]
  assign _T_1893 = {_T_1880,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21713.4]
  assign _T_1895 = {_T_1881,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21715.4]
  assign _T_1897 = {_T_1882,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21717.4]
  assign _T_1899 = {_T_1883,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21719.4]
  assign _T_1901 = {_T_1884,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21721.4]
  assign _T_1903 = {_T_1885,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21723.4]
  assign _T_1904 = _T_1884 ? _T_1901 : _T_1903; // @[Mux.scala 31:69:@21724.4]
  assign _T_1905 = _T_1883 ? _T_1899 : _T_1904; // @[Mux.scala 31:69:@21725.4]
  assign _T_1906 = _T_1882 ? _T_1897 : _T_1905; // @[Mux.scala 31:69:@21726.4]
  assign _T_1907 = _T_1881 ? _T_1895 : _T_1906; // @[Mux.scala 31:69:@21727.4]
  assign _T_1908 = _T_1880 ? _T_1893 : _T_1907; // @[Mux.scala 31:69:@21728.4]
  assign _T_1909 = _T_1879 ? _T_1891 : _T_1908; // @[Mux.scala 31:69:@21729.4]
  assign _T_1910 = _T_1878 ? _T_1889 : _T_1909; // @[Mux.scala 31:69:@21730.4]
  assign _T_1911 = _T_1877 ? _T_1887 : _T_1910; // @[Mux.scala 31:69:@21731.4]
  assign _T_1919 = _T_1732 & _T_1366; // @[MemPrimitives.scala 110:228:@21740.4]
  assign _T_1925 = _T_1738 & _T_1372; // @[MemPrimitives.scala 110:228:@21744.4]
  assign _T_1931 = _T_1744 & _T_1378; // @[MemPrimitives.scala 110:228:@21748.4]
  assign _T_1937 = _T_1750 & _T_1384; // @[MemPrimitives.scala 110:228:@21752.4]
  assign _T_1943 = _T_1756 & _T_1390; // @[MemPrimitives.scala 110:228:@21756.4]
  assign _T_1949 = _T_1762 & _T_1396; // @[MemPrimitives.scala 110:228:@21760.4]
  assign _T_1955 = _T_1768 & _T_1402; // @[MemPrimitives.scala 110:228:@21764.4]
  assign _T_1961 = _T_1774 & _T_1408; // @[MemPrimitives.scala 110:228:@21768.4]
  assign _T_1967 = _T_1780 & _T_1414; // @[MemPrimitives.scala 110:228:@21772.4]
  assign _T_1969 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@21786.4]
  assign _T_1970 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@21787.4]
  assign _T_1971 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 126:35:@21788.4]
  assign _T_1972 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 126:35:@21789.4]
  assign _T_1973 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 126:35:@21790.4]
  assign _T_1974 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 126:35:@21791.4]
  assign _T_1975 = StickySelects_8_io_outs_6; // @[MemPrimitives.scala 126:35:@21792.4]
  assign _T_1976 = StickySelects_8_io_outs_7; // @[MemPrimitives.scala 126:35:@21793.4]
  assign _T_1977 = StickySelects_8_io_outs_8; // @[MemPrimitives.scala 126:35:@21794.4]
  assign _T_1979 = {_T_1969,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21796.4]
  assign _T_1981 = {_T_1970,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21798.4]
  assign _T_1983 = {_T_1971,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21800.4]
  assign _T_1985 = {_T_1972,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21802.4]
  assign _T_1987 = {_T_1973,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21804.4]
  assign _T_1989 = {_T_1974,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21806.4]
  assign _T_1991 = {_T_1975,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21808.4]
  assign _T_1993 = {_T_1976,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21810.4]
  assign _T_1995 = {_T_1977,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21812.4]
  assign _T_1996 = _T_1976 ? _T_1993 : _T_1995; // @[Mux.scala 31:69:@21813.4]
  assign _T_1997 = _T_1975 ? _T_1991 : _T_1996; // @[Mux.scala 31:69:@21814.4]
  assign _T_1998 = _T_1974 ? _T_1989 : _T_1997; // @[Mux.scala 31:69:@21815.4]
  assign _T_1999 = _T_1973 ? _T_1987 : _T_1998; // @[Mux.scala 31:69:@21816.4]
  assign _T_2000 = _T_1972 ? _T_1985 : _T_1999; // @[Mux.scala 31:69:@21817.4]
  assign _T_2001 = _T_1971 ? _T_1983 : _T_2000; // @[Mux.scala 31:69:@21818.4]
  assign _T_2002 = _T_1970 ? _T_1981 : _T_2001; // @[Mux.scala 31:69:@21819.4]
  assign _T_2003 = _T_1969 ? _T_1979 : _T_2002; // @[Mux.scala 31:69:@21820.4]
  assign _T_2011 = _T_1824 & _T_1458; // @[MemPrimitives.scala 110:228:@21829.4]
  assign _T_2017 = _T_1830 & _T_1464; // @[MemPrimitives.scala 110:228:@21833.4]
  assign _T_2023 = _T_1836 & _T_1470; // @[MemPrimitives.scala 110:228:@21837.4]
  assign _T_2029 = _T_1842 & _T_1476; // @[MemPrimitives.scala 110:228:@21841.4]
  assign _T_2035 = _T_1848 & _T_1482; // @[MemPrimitives.scala 110:228:@21845.4]
  assign _T_2041 = _T_1854 & _T_1488; // @[MemPrimitives.scala 110:228:@21849.4]
  assign _T_2047 = _T_1860 & _T_1494; // @[MemPrimitives.scala 110:228:@21853.4]
  assign _T_2053 = _T_1866 & _T_1500; // @[MemPrimitives.scala 110:228:@21857.4]
  assign _T_2059 = _T_1872 & _T_1506; // @[MemPrimitives.scala 110:228:@21861.4]
  assign _T_2061 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@21875.4]
  assign _T_2062 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@21876.4]
  assign _T_2063 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@21877.4]
  assign _T_2064 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@21878.4]
  assign _T_2065 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 126:35:@21879.4]
  assign _T_2066 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 126:35:@21880.4]
  assign _T_2067 = StickySelects_9_io_outs_6; // @[MemPrimitives.scala 126:35:@21881.4]
  assign _T_2068 = StickySelects_9_io_outs_7; // @[MemPrimitives.scala 126:35:@21882.4]
  assign _T_2069 = StickySelects_9_io_outs_8; // @[MemPrimitives.scala 126:35:@21883.4]
  assign _T_2071 = {_T_2061,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21885.4]
  assign _T_2073 = {_T_2062,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21887.4]
  assign _T_2075 = {_T_2063,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21889.4]
  assign _T_2077 = {_T_2064,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21891.4]
  assign _T_2079 = {_T_2065,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21893.4]
  assign _T_2081 = {_T_2066,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21895.4]
  assign _T_2083 = {_T_2067,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21897.4]
  assign _T_2085 = {_T_2068,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21899.4]
  assign _T_2087 = {_T_2069,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21901.4]
  assign _T_2088 = _T_2068 ? _T_2085 : _T_2087; // @[Mux.scala 31:69:@21902.4]
  assign _T_2089 = _T_2067 ? _T_2083 : _T_2088; // @[Mux.scala 31:69:@21903.4]
  assign _T_2090 = _T_2066 ? _T_2081 : _T_2089; // @[Mux.scala 31:69:@21904.4]
  assign _T_2091 = _T_2065 ? _T_2079 : _T_2090; // @[Mux.scala 31:69:@21905.4]
  assign _T_2092 = _T_2064 ? _T_2077 : _T_2091; // @[Mux.scala 31:69:@21906.4]
  assign _T_2093 = _T_2063 ? _T_2075 : _T_2092; // @[Mux.scala 31:69:@21907.4]
  assign _T_2094 = _T_2062 ? _T_2073 : _T_2093; // @[Mux.scala 31:69:@21908.4]
  assign _T_2095 = _T_2061 ? _T_2071 : _T_2094; // @[Mux.scala 31:69:@21909.4]
  assign _T_2103 = _T_1732 & _T_1550; // @[MemPrimitives.scala 110:228:@21918.4]
  assign _T_2109 = _T_1738 & _T_1556; // @[MemPrimitives.scala 110:228:@21922.4]
  assign _T_2115 = _T_1744 & _T_1562; // @[MemPrimitives.scala 110:228:@21926.4]
  assign _T_2121 = _T_1750 & _T_1568; // @[MemPrimitives.scala 110:228:@21930.4]
  assign _T_2127 = _T_1756 & _T_1574; // @[MemPrimitives.scala 110:228:@21934.4]
  assign _T_2133 = _T_1762 & _T_1580; // @[MemPrimitives.scala 110:228:@21938.4]
  assign _T_2139 = _T_1768 & _T_1586; // @[MemPrimitives.scala 110:228:@21942.4]
  assign _T_2145 = _T_1774 & _T_1592; // @[MemPrimitives.scala 110:228:@21946.4]
  assign _T_2151 = _T_1780 & _T_1598; // @[MemPrimitives.scala 110:228:@21950.4]
  assign _T_2153 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@21964.4]
  assign _T_2154 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@21965.4]
  assign _T_2155 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 126:35:@21966.4]
  assign _T_2156 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 126:35:@21967.4]
  assign _T_2157 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 126:35:@21968.4]
  assign _T_2158 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 126:35:@21969.4]
  assign _T_2159 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 126:35:@21970.4]
  assign _T_2160 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 126:35:@21971.4]
  assign _T_2161 = StickySelects_10_io_outs_8; // @[MemPrimitives.scala 126:35:@21972.4]
  assign _T_2163 = {_T_2153,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21974.4]
  assign _T_2165 = {_T_2154,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21976.4]
  assign _T_2167 = {_T_2155,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21978.4]
  assign _T_2169 = {_T_2156,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21980.4]
  assign _T_2171 = {_T_2157,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21982.4]
  assign _T_2173 = {_T_2158,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21984.4]
  assign _T_2175 = {_T_2159,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21986.4]
  assign _T_2177 = {_T_2160,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21988.4]
  assign _T_2179 = {_T_2161,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21990.4]
  assign _T_2180 = _T_2160 ? _T_2177 : _T_2179; // @[Mux.scala 31:69:@21991.4]
  assign _T_2181 = _T_2159 ? _T_2175 : _T_2180; // @[Mux.scala 31:69:@21992.4]
  assign _T_2182 = _T_2158 ? _T_2173 : _T_2181; // @[Mux.scala 31:69:@21993.4]
  assign _T_2183 = _T_2157 ? _T_2171 : _T_2182; // @[Mux.scala 31:69:@21994.4]
  assign _T_2184 = _T_2156 ? _T_2169 : _T_2183; // @[Mux.scala 31:69:@21995.4]
  assign _T_2185 = _T_2155 ? _T_2167 : _T_2184; // @[Mux.scala 31:69:@21996.4]
  assign _T_2186 = _T_2154 ? _T_2165 : _T_2185; // @[Mux.scala 31:69:@21997.4]
  assign _T_2187 = _T_2153 ? _T_2163 : _T_2186; // @[Mux.scala 31:69:@21998.4]
  assign _T_2195 = _T_1824 & _T_1642; // @[MemPrimitives.scala 110:228:@22007.4]
  assign _T_2201 = _T_1830 & _T_1648; // @[MemPrimitives.scala 110:228:@22011.4]
  assign _T_2207 = _T_1836 & _T_1654; // @[MemPrimitives.scala 110:228:@22015.4]
  assign _T_2213 = _T_1842 & _T_1660; // @[MemPrimitives.scala 110:228:@22019.4]
  assign _T_2219 = _T_1848 & _T_1666; // @[MemPrimitives.scala 110:228:@22023.4]
  assign _T_2225 = _T_1854 & _T_1672; // @[MemPrimitives.scala 110:228:@22027.4]
  assign _T_2231 = _T_1860 & _T_1678; // @[MemPrimitives.scala 110:228:@22031.4]
  assign _T_2237 = _T_1866 & _T_1684; // @[MemPrimitives.scala 110:228:@22035.4]
  assign _T_2243 = _T_1872 & _T_1690; // @[MemPrimitives.scala 110:228:@22039.4]
  assign _T_2245 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@22053.4]
  assign _T_2246 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@22054.4]
  assign _T_2247 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@22055.4]
  assign _T_2248 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@22056.4]
  assign _T_2249 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 126:35:@22057.4]
  assign _T_2250 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 126:35:@22058.4]
  assign _T_2251 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 126:35:@22059.4]
  assign _T_2252 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 126:35:@22060.4]
  assign _T_2253 = StickySelects_11_io_outs_8; // @[MemPrimitives.scala 126:35:@22061.4]
  assign _T_2255 = {_T_2245,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22063.4]
  assign _T_2257 = {_T_2246,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22065.4]
  assign _T_2259 = {_T_2247,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22067.4]
  assign _T_2261 = {_T_2248,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22069.4]
  assign _T_2263 = {_T_2249,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22071.4]
  assign _T_2265 = {_T_2250,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22073.4]
  assign _T_2267 = {_T_2251,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22075.4]
  assign _T_2269 = {_T_2252,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22077.4]
  assign _T_2271 = {_T_2253,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22079.4]
  assign _T_2272 = _T_2252 ? _T_2269 : _T_2271; // @[Mux.scala 31:69:@22080.4]
  assign _T_2273 = _T_2251 ? _T_2267 : _T_2272; // @[Mux.scala 31:69:@22081.4]
  assign _T_2274 = _T_2250 ? _T_2265 : _T_2273; // @[Mux.scala 31:69:@22082.4]
  assign _T_2275 = _T_2249 ? _T_2263 : _T_2274; // @[Mux.scala 31:69:@22083.4]
  assign _T_2276 = _T_2248 ? _T_2261 : _T_2275; // @[Mux.scala 31:69:@22084.4]
  assign _T_2277 = _T_2247 ? _T_2259 : _T_2276; // @[Mux.scala 31:69:@22085.4]
  assign _T_2278 = _T_2246 ? _T_2257 : _T_2277; // @[Mux.scala 31:69:@22086.4]
  assign _T_2279 = _T_2245 ? _T_2255 : _T_2278; // @[Mux.scala 31:69:@22087.4]
  assign _T_2284 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22094.4]
  assign _T_2287 = _T_2284 & _T_1182; // @[MemPrimitives.scala 110:228:@22096.4]
  assign _T_2290 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22098.4]
  assign _T_2293 = _T_2290 & _T_1188; // @[MemPrimitives.scala 110:228:@22100.4]
  assign _T_2296 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22102.4]
  assign _T_2299 = _T_2296 & _T_1194; // @[MemPrimitives.scala 110:228:@22104.4]
  assign _T_2302 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22106.4]
  assign _T_2305 = _T_2302 & _T_1200; // @[MemPrimitives.scala 110:228:@22108.4]
  assign _T_2308 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22110.4]
  assign _T_2311 = _T_2308 & _T_1206; // @[MemPrimitives.scala 110:228:@22112.4]
  assign _T_2314 = io_rPort_12_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22114.4]
  assign _T_2317 = _T_2314 & _T_1212; // @[MemPrimitives.scala 110:228:@22116.4]
  assign _T_2320 = io_rPort_15_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22118.4]
  assign _T_2323 = _T_2320 & _T_1218; // @[MemPrimitives.scala 110:228:@22120.4]
  assign _T_2326 = io_rPort_16_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22122.4]
  assign _T_2329 = _T_2326 & _T_1224; // @[MemPrimitives.scala 110:228:@22124.4]
  assign _T_2332 = io_rPort_17_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22126.4]
  assign _T_2335 = _T_2332 & _T_1230; // @[MemPrimitives.scala 110:228:@22128.4]
  assign _T_2337 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 126:35:@22142.4]
  assign _T_2338 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 126:35:@22143.4]
  assign _T_2339 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 126:35:@22144.4]
  assign _T_2340 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 126:35:@22145.4]
  assign _T_2341 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 126:35:@22146.4]
  assign _T_2342 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 126:35:@22147.4]
  assign _T_2343 = StickySelects_12_io_outs_6; // @[MemPrimitives.scala 126:35:@22148.4]
  assign _T_2344 = StickySelects_12_io_outs_7; // @[MemPrimitives.scala 126:35:@22149.4]
  assign _T_2345 = StickySelects_12_io_outs_8; // @[MemPrimitives.scala 126:35:@22150.4]
  assign _T_2347 = {_T_2337,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22152.4]
  assign _T_2349 = {_T_2338,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22154.4]
  assign _T_2351 = {_T_2339,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22156.4]
  assign _T_2353 = {_T_2340,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22158.4]
  assign _T_2355 = {_T_2341,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22160.4]
  assign _T_2357 = {_T_2342,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22162.4]
  assign _T_2359 = {_T_2343,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22164.4]
  assign _T_2361 = {_T_2344,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22166.4]
  assign _T_2363 = {_T_2345,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22168.4]
  assign _T_2364 = _T_2344 ? _T_2361 : _T_2363; // @[Mux.scala 31:69:@22169.4]
  assign _T_2365 = _T_2343 ? _T_2359 : _T_2364; // @[Mux.scala 31:69:@22170.4]
  assign _T_2366 = _T_2342 ? _T_2357 : _T_2365; // @[Mux.scala 31:69:@22171.4]
  assign _T_2367 = _T_2341 ? _T_2355 : _T_2366; // @[Mux.scala 31:69:@22172.4]
  assign _T_2368 = _T_2340 ? _T_2353 : _T_2367; // @[Mux.scala 31:69:@22173.4]
  assign _T_2369 = _T_2339 ? _T_2351 : _T_2368; // @[Mux.scala 31:69:@22174.4]
  assign _T_2370 = _T_2338 ? _T_2349 : _T_2369; // @[Mux.scala 31:69:@22175.4]
  assign _T_2371 = _T_2337 ? _T_2347 : _T_2370; // @[Mux.scala 31:69:@22176.4]
  assign _T_2376 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22183.4]
  assign _T_2379 = _T_2376 & _T_1274; // @[MemPrimitives.scala 110:228:@22185.4]
  assign _T_2382 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22187.4]
  assign _T_2385 = _T_2382 & _T_1280; // @[MemPrimitives.scala 110:228:@22189.4]
  assign _T_2388 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22191.4]
  assign _T_2391 = _T_2388 & _T_1286; // @[MemPrimitives.scala 110:228:@22193.4]
  assign _T_2394 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22195.4]
  assign _T_2397 = _T_2394 & _T_1292; // @[MemPrimitives.scala 110:228:@22197.4]
  assign _T_2400 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22199.4]
  assign _T_2403 = _T_2400 & _T_1298; // @[MemPrimitives.scala 110:228:@22201.4]
  assign _T_2406 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22203.4]
  assign _T_2409 = _T_2406 & _T_1304; // @[MemPrimitives.scala 110:228:@22205.4]
  assign _T_2412 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22207.4]
  assign _T_2415 = _T_2412 & _T_1310; // @[MemPrimitives.scala 110:228:@22209.4]
  assign _T_2418 = io_rPort_13_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22211.4]
  assign _T_2421 = _T_2418 & _T_1316; // @[MemPrimitives.scala 110:228:@22213.4]
  assign _T_2424 = io_rPort_14_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@22215.4]
  assign _T_2427 = _T_2424 & _T_1322; // @[MemPrimitives.scala 110:228:@22217.4]
  assign _T_2429 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 126:35:@22231.4]
  assign _T_2430 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 126:35:@22232.4]
  assign _T_2431 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 126:35:@22233.4]
  assign _T_2432 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 126:35:@22234.4]
  assign _T_2433 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 126:35:@22235.4]
  assign _T_2434 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 126:35:@22236.4]
  assign _T_2435 = StickySelects_13_io_outs_6; // @[MemPrimitives.scala 126:35:@22237.4]
  assign _T_2436 = StickySelects_13_io_outs_7; // @[MemPrimitives.scala 126:35:@22238.4]
  assign _T_2437 = StickySelects_13_io_outs_8; // @[MemPrimitives.scala 126:35:@22239.4]
  assign _T_2439 = {_T_2429,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22241.4]
  assign _T_2441 = {_T_2430,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22243.4]
  assign _T_2443 = {_T_2431,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22245.4]
  assign _T_2445 = {_T_2432,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22247.4]
  assign _T_2447 = {_T_2433,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22249.4]
  assign _T_2449 = {_T_2434,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22251.4]
  assign _T_2451 = {_T_2435,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22253.4]
  assign _T_2453 = {_T_2436,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22255.4]
  assign _T_2455 = {_T_2437,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22257.4]
  assign _T_2456 = _T_2436 ? _T_2453 : _T_2455; // @[Mux.scala 31:69:@22258.4]
  assign _T_2457 = _T_2435 ? _T_2451 : _T_2456; // @[Mux.scala 31:69:@22259.4]
  assign _T_2458 = _T_2434 ? _T_2449 : _T_2457; // @[Mux.scala 31:69:@22260.4]
  assign _T_2459 = _T_2433 ? _T_2447 : _T_2458; // @[Mux.scala 31:69:@22261.4]
  assign _T_2460 = _T_2432 ? _T_2445 : _T_2459; // @[Mux.scala 31:69:@22262.4]
  assign _T_2461 = _T_2431 ? _T_2443 : _T_2460; // @[Mux.scala 31:69:@22263.4]
  assign _T_2462 = _T_2430 ? _T_2441 : _T_2461; // @[Mux.scala 31:69:@22264.4]
  assign _T_2463 = _T_2429 ? _T_2439 : _T_2462; // @[Mux.scala 31:69:@22265.4]
  assign _T_2471 = _T_2284 & _T_1366; // @[MemPrimitives.scala 110:228:@22274.4]
  assign _T_2477 = _T_2290 & _T_1372; // @[MemPrimitives.scala 110:228:@22278.4]
  assign _T_2483 = _T_2296 & _T_1378; // @[MemPrimitives.scala 110:228:@22282.4]
  assign _T_2489 = _T_2302 & _T_1384; // @[MemPrimitives.scala 110:228:@22286.4]
  assign _T_2495 = _T_2308 & _T_1390; // @[MemPrimitives.scala 110:228:@22290.4]
  assign _T_2501 = _T_2314 & _T_1396; // @[MemPrimitives.scala 110:228:@22294.4]
  assign _T_2507 = _T_2320 & _T_1402; // @[MemPrimitives.scala 110:228:@22298.4]
  assign _T_2513 = _T_2326 & _T_1408; // @[MemPrimitives.scala 110:228:@22302.4]
  assign _T_2519 = _T_2332 & _T_1414; // @[MemPrimitives.scala 110:228:@22306.4]
  assign _T_2521 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 126:35:@22320.4]
  assign _T_2522 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 126:35:@22321.4]
  assign _T_2523 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 126:35:@22322.4]
  assign _T_2524 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 126:35:@22323.4]
  assign _T_2525 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 126:35:@22324.4]
  assign _T_2526 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 126:35:@22325.4]
  assign _T_2527 = StickySelects_14_io_outs_6; // @[MemPrimitives.scala 126:35:@22326.4]
  assign _T_2528 = StickySelects_14_io_outs_7; // @[MemPrimitives.scala 126:35:@22327.4]
  assign _T_2529 = StickySelects_14_io_outs_8; // @[MemPrimitives.scala 126:35:@22328.4]
  assign _T_2531 = {_T_2521,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22330.4]
  assign _T_2533 = {_T_2522,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22332.4]
  assign _T_2535 = {_T_2523,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22334.4]
  assign _T_2537 = {_T_2524,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22336.4]
  assign _T_2539 = {_T_2525,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22338.4]
  assign _T_2541 = {_T_2526,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22340.4]
  assign _T_2543 = {_T_2527,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22342.4]
  assign _T_2545 = {_T_2528,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22344.4]
  assign _T_2547 = {_T_2529,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22346.4]
  assign _T_2548 = _T_2528 ? _T_2545 : _T_2547; // @[Mux.scala 31:69:@22347.4]
  assign _T_2549 = _T_2527 ? _T_2543 : _T_2548; // @[Mux.scala 31:69:@22348.4]
  assign _T_2550 = _T_2526 ? _T_2541 : _T_2549; // @[Mux.scala 31:69:@22349.4]
  assign _T_2551 = _T_2525 ? _T_2539 : _T_2550; // @[Mux.scala 31:69:@22350.4]
  assign _T_2552 = _T_2524 ? _T_2537 : _T_2551; // @[Mux.scala 31:69:@22351.4]
  assign _T_2553 = _T_2523 ? _T_2535 : _T_2552; // @[Mux.scala 31:69:@22352.4]
  assign _T_2554 = _T_2522 ? _T_2533 : _T_2553; // @[Mux.scala 31:69:@22353.4]
  assign _T_2555 = _T_2521 ? _T_2531 : _T_2554; // @[Mux.scala 31:69:@22354.4]
  assign _T_2563 = _T_2376 & _T_1458; // @[MemPrimitives.scala 110:228:@22363.4]
  assign _T_2569 = _T_2382 & _T_1464; // @[MemPrimitives.scala 110:228:@22367.4]
  assign _T_2575 = _T_2388 & _T_1470; // @[MemPrimitives.scala 110:228:@22371.4]
  assign _T_2581 = _T_2394 & _T_1476; // @[MemPrimitives.scala 110:228:@22375.4]
  assign _T_2587 = _T_2400 & _T_1482; // @[MemPrimitives.scala 110:228:@22379.4]
  assign _T_2593 = _T_2406 & _T_1488; // @[MemPrimitives.scala 110:228:@22383.4]
  assign _T_2599 = _T_2412 & _T_1494; // @[MemPrimitives.scala 110:228:@22387.4]
  assign _T_2605 = _T_2418 & _T_1500; // @[MemPrimitives.scala 110:228:@22391.4]
  assign _T_2611 = _T_2424 & _T_1506; // @[MemPrimitives.scala 110:228:@22395.4]
  assign _T_2613 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 126:35:@22409.4]
  assign _T_2614 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 126:35:@22410.4]
  assign _T_2615 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 126:35:@22411.4]
  assign _T_2616 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 126:35:@22412.4]
  assign _T_2617 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 126:35:@22413.4]
  assign _T_2618 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 126:35:@22414.4]
  assign _T_2619 = StickySelects_15_io_outs_6; // @[MemPrimitives.scala 126:35:@22415.4]
  assign _T_2620 = StickySelects_15_io_outs_7; // @[MemPrimitives.scala 126:35:@22416.4]
  assign _T_2621 = StickySelects_15_io_outs_8; // @[MemPrimitives.scala 126:35:@22417.4]
  assign _T_2623 = {_T_2613,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22419.4]
  assign _T_2625 = {_T_2614,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22421.4]
  assign _T_2627 = {_T_2615,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22423.4]
  assign _T_2629 = {_T_2616,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22425.4]
  assign _T_2631 = {_T_2617,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22427.4]
  assign _T_2633 = {_T_2618,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22429.4]
  assign _T_2635 = {_T_2619,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22431.4]
  assign _T_2637 = {_T_2620,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22433.4]
  assign _T_2639 = {_T_2621,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22435.4]
  assign _T_2640 = _T_2620 ? _T_2637 : _T_2639; // @[Mux.scala 31:69:@22436.4]
  assign _T_2641 = _T_2619 ? _T_2635 : _T_2640; // @[Mux.scala 31:69:@22437.4]
  assign _T_2642 = _T_2618 ? _T_2633 : _T_2641; // @[Mux.scala 31:69:@22438.4]
  assign _T_2643 = _T_2617 ? _T_2631 : _T_2642; // @[Mux.scala 31:69:@22439.4]
  assign _T_2644 = _T_2616 ? _T_2629 : _T_2643; // @[Mux.scala 31:69:@22440.4]
  assign _T_2645 = _T_2615 ? _T_2627 : _T_2644; // @[Mux.scala 31:69:@22441.4]
  assign _T_2646 = _T_2614 ? _T_2625 : _T_2645; // @[Mux.scala 31:69:@22442.4]
  assign _T_2647 = _T_2613 ? _T_2623 : _T_2646; // @[Mux.scala 31:69:@22443.4]
  assign _T_2655 = _T_2284 & _T_1550; // @[MemPrimitives.scala 110:228:@22452.4]
  assign _T_2661 = _T_2290 & _T_1556; // @[MemPrimitives.scala 110:228:@22456.4]
  assign _T_2667 = _T_2296 & _T_1562; // @[MemPrimitives.scala 110:228:@22460.4]
  assign _T_2673 = _T_2302 & _T_1568; // @[MemPrimitives.scala 110:228:@22464.4]
  assign _T_2679 = _T_2308 & _T_1574; // @[MemPrimitives.scala 110:228:@22468.4]
  assign _T_2685 = _T_2314 & _T_1580; // @[MemPrimitives.scala 110:228:@22472.4]
  assign _T_2691 = _T_2320 & _T_1586; // @[MemPrimitives.scala 110:228:@22476.4]
  assign _T_2697 = _T_2326 & _T_1592; // @[MemPrimitives.scala 110:228:@22480.4]
  assign _T_2703 = _T_2332 & _T_1598; // @[MemPrimitives.scala 110:228:@22484.4]
  assign _T_2705 = StickySelects_16_io_outs_0; // @[MemPrimitives.scala 126:35:@22498.4]
  assign _T_2706 = StickySelects_16_io_outs_1; // @[MemPrimitives.scala 126:35:@22499.4]
  assign _T_2707 = StickySelects_16_io_outs_2; // @[MemPrimitives.scala 126:35:@22500.4]
  assign _T_2708 = StickySelects_16_io_outs_3; // @[MemPrimitives.scala 126:35:@22501.4]
  assign _T_2709 = StickySelects_16_io_outs_4; // @[MemPrimitives.scala 126:35:@22502.4]
  assign _T_2710 = StickySelects_16_io_outs_5; // @[MemPrimitives.scala 126:35:@22503.4]
  assign _T_2711 = StickySelects_16_io_outs_6; // @[MemPrimitives.scala 126:35:@22504.4]
  assign _T_2712 = StickySelects_16_io_outs_7; // @[MemPrimitives.scala 126:35:@22505.4]
  assign _T_2713 = StickySelects_16_io_outs_8; // @[MemPrimitives.scala 126:35:@22506.4]
  assign _T_2715 = {_T_2705,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22508.4]
  assign _T_2717 = {_T_2706,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22510.4]
  assign _T_2719 = {_T_2707,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22512.4]
  assign _T_2721 = {_T_2708,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22514.4]
  assign _T_2723 = {_T_2709,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22516.4]
  assign _T_2725 = {_T_2710,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22518.4]
  assign _T_2727 = {_T_2711,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22520.4]
  assign _T_2729 = {_T_2712,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22522.4]
  assign _T_2731 = {_T_2713,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22524.4]
  assign _T_2732 = _T_2712 ? _T_2729 : _T_2731; // @[Mux.scala 31:69:@22525.4]
  assign _T_2733 = _T_2711 ? _T_2727 : _T_2732; // @[Mux.scala 31:69:@22526.4]
  assign _T_2734 = _T_2710 ? _T_2725 : _T_2733; // @[Mux.scala 31:69:@22527.4]
  assign _T_2735 = _T_2709 ? _T_2723 : _T_2734; // @[Mux.scala 31:69:@22528.4]
  assign _T_2736 = _T_2708 ? _T_2721 : _T_2735; // @[Mux.scala 31:69:@22529.4]
  assign _T_2737 = _T_2707 ? _T_2719 : _T_2736; // @[Mux.scala 31:69:@22530.4]
  assign _T_2738 = _T_2706 ? _T_2717 : _T_2737; // @[Mux.scala 31:69:@22531.4]
  assign _T_2739 = _T_2705 ? _T_2715 : _T_2738; // @[Mux.scala 31:69:@22532.4]
  assign _T_2747 = _T_2376 & _T_1642; // @[MemPrimitives.scala 110:228:@22541.4]
  assign _T_2753 = _T_2382 & _T_1648; // @[MemPrimitives.scala 110:228:@22545.4]
  assign _T_2759 = _T_2388 & _T_1654; // @[MemPrimitives.scala 110:228:@22549.4]
  assign _T_2765 = _T_2394 & _T_1660; // @[MemPrimitives.scala 110:228:@22553.4]
  assign _T_2771 = _T_2400 & _T_1666; // @[MemPrimitives.scala 110:228:@22557.4]
  assign _T_2777 = _T_2406 & _T_1672; // @[MemPrimitives.scala 110:228:@22561.4]
  assign _T_2783 = _T_2412 & _T_1678; // @[MemPrimitives.scala 110:228:@22565.4]
  assign _T_2789 = _T_2418 & _T_1684; // @[MemPrimitives.scala 110:228:@22569.4]
  assign _T_2795 = _T_2424 & _T_1690; // @[MemPrimitives.scala 110:228:@22573.4]
  assign _T_2797 = StickySelects_17_io_outs_0; // @[MemPrimitives.scala 126:35:@22587.4]
  assign _T_2798 = StickySelects_17_io_outs_1; // @[MemPrimitives.scala 126:35:@22588.4]
  assign _T_2799 = StickySelects_17_io_outs_2; // @[MemPrimitives.scala 126:35:@22589.4]
  assign _T_2800 = StickySelects_17_io_outs_3; // @[MemPrimitives.scala 126:35:@22590.4]
  assign _T_2801 = StickySelects_17_io_outs_4; // @[MemPrimitives.scala 126:35:@22591.4]
  assign _T_2802 = StickySelects_17_io_outs_5; // @[MemPrimitives.scala 126:35:@22592.4]
  assign _T_2803 = StickySelects_17_io_outs_6; // @[MemPrimitives.scala 126:35:@22593.4]
  assign _T_2804 = StickySelects_17_io_outs_7; // @[MemPrimitives.scala 126:35:@22594.4]
  assign _T_2805 = StickySelects_17_io_outs_8; // @[MemPrimitives.scala 126:35:@22595.4]
  assign _T_2807 = {_T_2797,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22597.4]
  assign _T_2809 = {_T_2798,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22599.4]
  assign _T_2811 = {_T_2799,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22601.4]
  assign _T_2813 = {_T_2800,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22603.4]
  assign _T_2815 = {_T_2801,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22605.4]
  assign _T_2817 = {_T_2802,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22607.4]
  assign _T_2819 = {_T_2803,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22609.4]
  assign _T_2821 = {_T_2804,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22611.4]
  assign _T_2823 = {_T_2805,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22613.4]
  assign _T_2824 = _T_2804 ? _T_2821 : _T_2823; // @[Mux.scala 31:69:@22614.4]
  assign _T_2825 = _T_2803 ? _T_2819 : _T_2824; // @[Mux.scala 31:69:@22615.4]
  assign _T_2826 = _T_2802 ? _T_2817 : _T_2825; // @[Mux.scala 31:69:@22616.4]
  assign _T_2827 = _T_2801 ? _T_2815 : _T_2826; // @[Mux.scala 31:69:@22617.4]
  assign _T_2828 = _T_2800 ? _T_2813 : _T_2827; // @[Mux.scala 31:69:@22618.4]
  assign _T_2829 = _T_2799 ? _T_2811 : _T_2828; // @[Mux.scala 31:69:@22619.4]
  assign _T_2830 = _T_2798 ? _T_2809 : _T_2829; // @[Mux.scala 31:69:@22620.4]
  assign _T_2831 = _T_2797 ? _T_2807 : _T_2830; // @[Mux.scala 31:69:@22621.4]
  assign _T_2836 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22628.4]
  assign _T_2839 = _T_2836 & _T_1182; // @[MemPrimitives.scala 110:228:@22630.4]
  assign _T_2842 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22632.4]
  assign _T_2845 = _T_2842 & _T_1188; // @[MemPrimitives.scala 110:228:@22634.4]
  assign _T_2848 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22636.4]
  assign _T_2851 = _T_2848 & _T_1194; // @[MemPrimitives.scala 110:228:@22638.4]
  assign _T_2854 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22640.4]
  assign _T_2857 = _T_2854 & _T_1200; // @[MemPrimitives.scala 110:228:@22642.4]
  assign _T_2860 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22644.4]
  assign _T_2863 = _T_2860 & _T_1206; // @[MemPrimitives.scala 110:228:@22646.4]
  assign _T_2866 = io_rPort_12_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22648.4]
  assign _T_2869 = _T_2866 & _T_1212; // @[MemPrimitives.scala 110:228:@22650.4]
  assign _T_2872 = io_rPort_15_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22652.4]
  assign _T_2875 = _T_2872 & _T_1218; // @[MemPrimitives.scala 110:228:@22654.4]
  assign _T_2878 = io_rPort_16_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22656.4]
  assign _T_2881 = _T_2878 & _T_1224; // @[MemPrimitives.scala 110:228:@22658.4]
  assign _T_2884 = io_rPort_17_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22660.4]
  assign _T_2887 = _T_2884 & _T_1230; // @[MemPrimitives.scala 110:228:@22662.4]
  assign _T_2889 = StickySelects_18_io_outs_0; // @[MemPrimitives.scala 126:35:@22676.4]
  assign _T_2890 = StickySelects_18_io_outs_1; // @[MemPrimitives.scala 126:35:@22677.4]
  assign _T_2891 = StickySelects_18_io_outs_2; // @[MemPrimitives.scala 126:35:@22678.4]
  assign _T_2892 = StickySelects_18_io_outs_3; // @[MemPrimitives.scala 126:35:@22679.4]
  assign _T_2893 = StickySelects_18_io_outs_4; // @[MemPrimitives.scala 126:35:@22680.4]
  assign _T_2894 = StickySelects_18_io_outs_5; // @[MemPrimitives.scala 126:35:@22681.4]
  assign _T_2895 = StickySelects_18_io_outs_6; // @[MemPrimitives.scala 126:35:@22682.4]
  assign _T_2896 = StickySelects_18_io_outs_7; // @[MemPrimitives.scala 126:35:@22683.4]
  assign _T_2897 = StickySelects_18_io_outs_8; // @[MemPrimitives.scala 126:35:@22684.4]
  assign _T_2899 = {_T_2889,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22686.4]
  assign _T_2901 = {_T_2890,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22688.4]
  assign _T_2903 = {_T_2891,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22690.4]
  assign _T_2905 = {_T_2892,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22692.4]
  assign _T_2907 = {_T_2893,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22694.4]
  assign _T_2909 = {_T_2894,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22696.4]
  assign _T_2911 = {_T_2895,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22698.4]
  assign _T_2913 = {_T_2896,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22700.4]
  assign _T_2915 = {_T_2897,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22702.4]
  assign _T_2916 = _T_2896 ? _T_2913 : _T_2915; // @[Mux.scala 31:69:@22703.4]
  assign _T_2917 = _T_2895 ? _T_2911 : _T_2916; // @[Mux.scala 31:69:@22704.4]
  assign _T_2918 = _T_2894 ? _T_2909 : _T_2917; // @[Mux.scala 31:69:@22705.4]
  assign _T_2919 = _T_2893 ? _T_2907 : _T_2918; // @[Mux.scala 31:69:@22706.4]
  assign _T_2920 = _T_2892 ? _T_2905 : _T_2919; // @[Mux.scala 31:69:@22707.4]
  assign _T_2921 = _T_2891 ? _T_2903 : _T_2920; // @[Mux.scala 31:69:@22708.4]
  assign _T_2922 = _T_2890 ? _T_2901 : _T_2921; // @[Mux.scala 31:69:@22709.4]
  assign _T_2923 = _T_2889 ? _T_2899 : _T_2922; // @[Mux.scala 31:69:@22710.4]
  assign _T_2928 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22717.4]
  assign _T_2931 = _T_2928 & _T_1274; // @[MemPrimitives.scala 110:228:@22719.4]
  assign _T_2934 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22721.4]
  assign _T_2937 = _T_2934 & _T_1280; // @[MemPrimitives.scala 110:228:@22723.4]
  assign _T_2940 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22725.4]
  assign _T_2943 = _T_2940 & _T_1286; // @[MemPrimitives.scala 110:228:@22727.4]
  assign _T_2946 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22729.4]
  assign _T_2949 = _T_2946 & _T_1292; // @[MemPrimitives.scala 110:228:@22731.4]
  assign _T_2952 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22733.4]
  assign _T_2955 = _T_2952 & _T_1298; // @[MemPrimitives.scala 110:228:@22735.4]
  assign _T_2958 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22737.4]
  assign _T_2961 = _T_2958 & _T_1304; // @[MemPrimitives.scala 110:228:@22739.4]
  assign _T_2964 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22741.4]
  assign _T_2967 = _T_2964 & _T_1310; // @[MemPrimitives.scala 110:228:@22743.4]
  assign _T_2970 = io_rPort_13_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22745.4]
  assign _T_2973 = _T_2970 & _T_1316; // @[MemPrimitives.scala 110:228:@22747.4]
  assign _T_2976 = io_rPort_14_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@22749.4]
  assign _T_2979 = _T_2976 & _T_1322; // @[MemPrimitives.scala 110:228:@22751.4]
  assign _T_2981 = StickySelects_19_io_outs_0; // @[MemPrimitives.scala 126:35:@22765.4]
  assign _T_2982 = StickySelects_19_io_outs_1; // @[MemPrimitives.scala 126:35:@22766.4]
  assign _T_2983 = StickySelects_19_io_outs_2; // @[MemPrimitives.scala 126:35:@22767.4]
  assign _T_2984 = StickySelects_19_io_outs_3; // @[MemPrimitives.scala 126:35:@22768.4]
  assign _T_2985 = StickySelects_19_io_outs_4; // @[MemPrimitives.scala 126:35:@22769.4]
  assign _T_2986 = StickySelects_19_io_outs_5; // @[MemPrimitives.scala 126:35:@22770.4]
  assign _T_2987 = StickySelects_19_io_outs_6; // @[MemPrimitives.scala 126:35:@22771.4]
  assign _T_2988 = StickySelects_19_io_outs_7; // @[MemPrimitives.scala 126:35:@22772.4]
  assign _T_2989 = StickySelects_19_io_outs_8; // @[MemPrimitives.scala 126:35:@22773.4]
  assign _T_2991 = {_T_2981,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22775.4]
  assign _T_2993 = {_T_2982,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22777.4]
  assign _T_2995 = {_T_2983,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22779.4]
  assign _T_2997 = {_T_2984,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22781.4]
  assign _T_2999 = {_T_2985,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22783.4]
  assign _T_3001 = {_T_2986,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22785.4]
  assign _T_3003 = {_T_2987,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22787.4]
  assign _T_3005 = {_T_2988,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22789.4]
  assign _T_3007 = {_T_2989,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22791.4]
  assign _T_3008 = _T_2988 ? _T_3005 : _T_3007; // @[Mux.scala 31:69:@22792.4]
  assign _T_3009 = _T_2987 ? _T_3003 : _T_3008; // @[Mux.scala 31:69:@22793.4]
  assign _T_3010 = _T_2986 ? _T_3001 : _T_3009; // @[Mux.scala 31:69:@22794.4]
  assign _T_3011 = _T_2985 ? _T_2999 : _T_3010; // @[Mux.scala 31:69:@22795.4]
  assign _T_3012 = _T_2984 ? _T_2997 : _T_3011; // @[Mux.scala 31:69:@22796.4]
  assign _T_3013 = _T_2983 ? _T_2995 : _T_3012; // @[Mux.scala 31:69:@22797.4]
  assign _T_3014 = _T_2982 ? _T_2993 : _T_3013; // @[Mux.scala 31:69:@22798.4]
  assign _T_3015 = _T_2981 ? _T_2991 : _T_3014; // @[Mux.scala 31:69:@22799.4]
  assign _T_3023 = _T_2836 & _T_1366; // @[MemPrimitives.scala 110:228:@22808.4]
  assign _T_3029 = _T_2842 & _T_1372; // @[MemPrimitives.scala 110:228:@22812.4]
  assign _T_3035 = _T_2848 & _T_1378; // @[MemPrimitives.scala 110:228:@22816.4]
  assign _T_3041 = _T_2854 & _T_1384; // @[MemPrimitives.scala 110:228:@22820.4]
  assign _T_3047 = _T_2860 & _T_1390; // @[MemPrimitives.scala 110:228:@22824.4]
  assign _T_3053 = _T_2866 & _T_1396; // @[MemPrimitives.scala 110:228:@22828.4]
  assign _T_3059 = _T_2872 & _T_1402; // @[MemPrimitives.scala 110:228:@22832.4]
  assign _T_3065 = _T_2878 & _T_1408; // @[MemPrimitives.scala 110:228:@22836.4]
  assign _T_3071 = _T_2884 & _T_1414; // @[MemPrimitives.scala 110:228:@22840.4]
  assign _T_3073 = StickySelects_20_io_outs_0; // @[MemPrimitives.scala 126:35:@22854.4]
  assign _T_3074 = StickySelects_20_io_outs_1; // @[MemPrimitives.scala 126:35:@22855.4]
  assign _T_3075 = StickySelects_20_io_outs_2; // @[MemPrimitives.scala 126:35:@22856.4]
  assign _T_3076 = StickySelects_20_io_outs_3; // @[MemPrimitives.scala 126:35:@22857.4]
  assign _T_3077 = StickySelects_20_io_outs_4; // @[MemPrimitives.scala 126:35:@22858.4]
  assign _T_3078 = StickySelects_20_io_outs_5; // @[MemPrimitives.scala 126:35:@22859.4]
  assign _T_3079 = StickySelects_20_io_outs_6; // @[MemPrimitives.scala 126:35:@22860.4]
  assign _T_3080 = StickySelects_20_io_outs_7; // @[MemPrimitives.scala 126:35:@22861.4]
  assign _T_3081 = StickySelects_20_io_outs_8; // @[MemPrimitives.scala 126:35:@22862.4]
  assign _T_3083 = {_T_3073,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22864.4]
  assign _T_3085 = {_T_3074,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22866.4]
  assign _T_3087 = {_T_3075,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22868.4]
  assign _T_3089 = {_T_3076,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22870.4]
  assign _T_3091 = {_T_3077,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22872.4]
  assign _T_3093 = {_T_3078,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22874.4]
  assign _T_3095 = {_T_3079,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22876.4]
  assign _T_3097 = {_T_3080,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22878.4]
  assign _T_3099 = {_T_3081,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22880.4]
  assign _T_3100 = _T_3080 ? _T_3097 : _T_3099; // @[Mux.scala 31:69:@22881.4]
  assign _T_3101 = _T_3079 ? _T_3095 : _T_3100; // @[Mux.scala 31:69:@22882.4]
  assign _T_3102 = _T_3078 ? _T_3093 : _T_3101; // @[Mux.scala 31:69:@22883.4]
  assign _T_3103 = _T_3077 ? _T_3091 : _T_3102; // @[Mux.scala 31:69:@22884.4]
  assign _T_3104 = _T_3076 ? _T_3089 : _T_3103; // @[Mux.scala 31:69:@22885.4]
  assign _T_3105 = _T_3075 ? _T_3087 : _T_3104; // @[Mux.scala 31:69:@22886.4]
  assign _T_3106 = _T_3074 ? _T_3085 : _T_3105; // @[Mux.scala 31:69:@22887.4]
  assign _T_3107 = _T_3073 ? _T_3083 : _T_3106; // @[Mux.scala 31:69:@22888.4]
  assign _T_3115 = _T_2928 & _T_1458; // @[MemPrimitives.scala 110:228:@22897.4]
  assign _T_3121 = _T_2934 & _T_1464; // @[MemPrimitives.scala 110:228:@22901.4]
  assign _T_3127 = _T_2940 & _T_1470; // @[MemPrimitives.scala 110:228:@22905.4]
  assign _T_3133 = _T_2946 & _T_1476; // @[MemPrimitives.scala 110:228:@22909.4]
  assign _T_3139 = _T_2952 & _T_1482; // @[MemPrimitives.scala 110:228:@22913.4]
  assign _T_3145 = _T_2958 & _T_1488; // @[MemPrimitives.scala 110:228:@22917.4]
  assign _T_3151 = _T_2964 & _T_1494; // @[MemPrimitives.scala 110:228:@22921.4]
  assign _T_3157 = _T_2970 & _T_1500; // @[MemPrimitives.scala 110:228:@22925.4]
  assign _T_3163 = _T_2976 & _T_1506; // @[MemPrimitives.scala 110:228:@22929.4]
  assign _T_3165 = StickySelects_21_io_outs_0; // @[MemPrimitives.scala 126:35:@22943.4]
  assign _T_3166 = StickySelects_21_io_outs_1; // @[MemPrimitives.scala 126:35:@22944.4]
  assign _T_3167 = StickySelects_21_io_outs_2; // @[MemPrimitives.scala 126:35:@22945.4]
  assign _T_3168 = StickySelects_21_io_outs_3; // @[MemPrimitives.scala 126:35:@22946.4]
  assign _T_3169 = StickySelects_21_io_outs_4; // @[MemPrimitives.scala 126:35:@22947.4]
  assign _T_3170 = StickySelects_21_io_outs_5; // @[MemPrimitives.scala 126:35:@22948.4]
  assign _T_3171 = StickySelects_21_io_outs_6; // @[MemPrimitives.scala 126:35:@22949.4]
  assign _T_3172 = StickySelects_21_io_outs_7; // @[MemPrimitives.scala 126:35:@22950.4]
  assign _T_3173 = StickySelects_21_io_outs_8; // @[MemPrimitives.scala 126:35:@22951.4]
  assign _T_3175 = {_T_3165,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22953.4]
  assign _T_3177 = {_T_3166,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22955.4]
  assign _T_3179 = {_T_3167,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22957.4]
  assign _T_3181 = {_T_3168,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22959.4]
  assign _T_3183 = {_T_3169,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22961.4]
  assign _T_3185 = {_T_3170,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22963.4]
  assign _T_3187 = {_T_3171,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22965.4]
  assign _T_3189 = {_T_3172,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22967.4]
  assign _T_3191 = {_T_3173,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22969.4]
  assign _T_3192 = _T_3172 ? _T_3189 : _T_3191; // @[Mux.scala 31:69:@22970.4]
  assign _T_3193 = _T_3171 ? _T_3187 : _T_3192; // @[Mux.scala 31:69:@22971.4]
  assign _T_3194 = _T_3170 ? _T_3185 : _T_3193; // @[Mux.scala 31:69:@22972.4]
  assign _T_3195 = _T_3169 ? _T_3183 : _T_3194; // @[Mux.scala 31:69:@22973.4]
  assign _T_3196 = _T_3168 ? _T_3181 : _T_3195; // @[Mux.scala 31:69:@22974.4]
  assign _T_3197 = _T_3167 ? _T_3179 : _T_3196; // @[Mux.scala 31:69:@22975.4]
  assign _T_3198 = _T_3166 ? _T_3177 : _T_3197; // @[Mux.scala 31:69:@22976.4]
  assign _T_3199 = _T_3165 ? _T_3175 : _T_3198; // @[Mux.scala 31:69:@22977.4]
  assign _T_3207 = _T_2836 & _T_1550; // @[MemPrimitives.scala 110:228:@22986.4]
  assign _T_3213 = _T_2842 & _T_1556; // @[MemPrimitives.scala 110:228:@22990.4]
  assign _T_3219 = _T_2848 & _T_1562; // @[MemPrimitives.scala 110:228:@22994.4]
  assign _T_3225 = _T_2854 & _T_1568; // @[MemPrimitives.scala 110:228:@22998.4]
  assign _T_3231 = _T_2860 & _T_1574; // @[MemPrimitives.scala 110:228:@23002.4]
  assign _T_3237 = _T_2866 & _T_1580; // @[MemPrimitives.scala 110:228:@23006.4]
  assign _T_3243 = _T_2872 & _T_1586; // @[MemPrimitives.scala 110:228:@23010.4]
  assign _T_3249 = _T_2878 & _T_1592; // @[MemPrimitives.scala 110:228:@23014.4]
  assign _T_3255 = _T_2884 & _T_1598; // @[MemPrimitives.scala 110:228:@23018.4]
  assign _T_3257 = StickySelects_22_io_outs_0; // @[MemPrimitives.scala 126:35:@23032.4]
  assign _T_3258 = StickySelects_22_io_outs_1; // @[MemPrimitives.scala 126:35:@23033.4]
  assign _T_3259 = StickySelects_22_io_outs_2; // @[MemPrimitives.scala 126:35:@23034.4]
  assign _T_3260 = StickySelects_22_io_outs_3; // @[MemPrimitives.scala 126:35:@23035.4]
  assign _T_3261 = StickySelects_22_io_outs_4; // @[MemPrimitives.scala 126:35:@23036.4]
  assign _T_3262 = StickySelects_22_io_outs_5; // @[MemPrimitives.scala 126:35:@23037.4]
  assign _T_3263 = StickySelects_22_io_outs_6; // @[MemPrimitives.scala 126:35:@23038.4]
  assign _T_3264 = StickySelects_22_io_outs_7; // @[MemPrimitives.scala 126:35:@23039.4]
  assign _T_3265 = StickySelects_22_io_outs_8; // @[MemPrimitives.scala 126:35:@23040.4]
  assign _T_3267 = {_T_3257,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@23042.4]
  assign _T_3269 = {_T_3258,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@23044.4]
  assign _T_3271 = {_T_3259,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@23046.4]
  assign _T_3273 = {_T_3260,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@23048.4]
  assign _T_3275 = {_T_3261,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@23050.4]
  assign _T_3277 = {_T_3262,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@23052.4]
  assign _T_3279 = {_T_3263,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@23054.4]
  assign _T_3281 = {_T_3264,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@23056.4]
  assign _T_3283 = {_T_3265,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@23058.4]
  assign _T_3284 = _T_3264 ? _T_3281 : _T_3283; // @[Mux.scala 31:69:@23059.4]
  assign _T_3285 = _T_3263 ? _T_3279 : _T_3284; // @[Mux.scala 31:69:@23060.4]
  assign _T_3286 = _T_3262 ? _T_3277 : _T_3285; // @[Mux.scala 31:69:@23061.4]
  assign _T_3287 = _T_3261 ? _T_3275 : _T_3286; // @[Mux.scala 31:69:@23062.4]
  assign _T_3288 = _T_3260 ? _T_3273 : _T_3287; // @[Mux.scala 31:69:@23063.4]
  assign _T_3289 = _T_3259 ? _T_3271 : _T_3288; // @[Mux.scala 31:69:@23064.4]
  assign _T_3290 = _T_3258 ? _T_3269 : _T_3289; // @[Mux.scala 31:69:@23065.4]
  assign _T_3291 = _T_3257 ? _T_3267 : _T_3290; // @[Mux.scala 31:69:@23066.4]
  assign _T_3299 = _T_2928 & _T_1642; // @[MemPrimitives.scala 110:228:@23075.4]
  assign _T_3305 = _T_2934 & _T_1648; // @[MemPrimitives.scala 110:228:@23079.4]
  assign _T_3311 = _T_2940 & _T_1654; // @[MemPrimitives.scala 110:228:@23083.4]
  assign _T_3317 = _T_2946 & _T_1660; // @[MemPrimitives.scala 110:228:@23087.4]
  assign _T_3323 = _T_2952 & _T_1666; // @[MemPrimitives.scala 110:228:@23091.4]
  assign _T_3329 = _T_2958 & _T_1672; // @[MemPrimitives.scala 110:228:@23095.4]
  assign _T_3335 = _T_2964 & _T_1678; // @[MemPrimitives.scala 110:228:@23099.4]
  assign _T_3341 = _T_2970 & _T_1684; // @[MemPrimitives.scala 110:228:@23103.4]
  assign _T_3347 = _T_2976 & _T_1690; // @[MemPrimitives.scala 110:228:@23107.4]
  assign _T_3349 = StickySelects_23_io_outs_0; // @[MemPrimitives.scala 126:35:@23121.4]
  assign _T_3350 = StickySelects_23_io_outs_1; // @[MemPrimitives.scala 126:35:@23122.4]
  assign _T_3351 = StickySelects_23_io_outs_2; // @[MemPrimitives.scala 126:35:@23123.4]
  assign _T_3352 = StickySelects_23_io_outs_3; // @[MemPrimitives.scala 126:35:@23124.4]
  assign _T_3353 = StickySelects_23_io_outs_4; // @[MemPrimitives.scala 126:35:@23125.4]
  assign _T_3354 = StickySelects_23_io_outs_5; // @[MemPrimitives.scala 126:35:@23126.4]
  assign _T_3355 = StickySelects_23_io_outs_6; // @[MemPrimitives.scala 126:35:@23127.4]
  assign _T_3356 = StickySelects_23_io_outs_7; // @[MemPrimitives.scala 126:35:@23128.4]
  assign _T_3357 = StickySelects_23_io_outs_8; // @[MemPrimitives.scala 126:35:@23129.4]
  assign _T_3359 = {_T_3349,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@23131.4]
  assign _T_3361 = {_T_3350,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@23133.4]
  assign _T_3363 = {_T_3351,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@23135.4]
  assign _T_3365 = {_T_3352,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@23137.4]
  assign _T_3367 = {_T_3353,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@23139.4]
  assign _T_3369 = {_T_3354,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@23141.4]
  assign _T_3371 = {_T_3355,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@23143.4]
  assign _T_3373 = {_T_3356,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@23145.4]
  assign _T_3375 = {_T_3357,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@23147.4]
  assign _T_3376 = _T_3356 ? _T_3373 : _T_3375; // @[Mux.scala 31:69:@23148.4]
  assign _T_3377 = _T_3355 ? _T_3371 : _T_3376; // @[Mux.scala 31:69:@23149.4]
  assign _T_3378 = _T_3354 ? _T_3369 : _T_3377; // @[Mux.scala 31:69:@23150.4]
  assign _T_3379 = _T_3353 ? _T_3367 : _T_3378; // @[Mux.scala 31:69:@23151.4]
  assign _T_3380 = _T_3352 ? _T_3365 : _T_3379; // @[Mux.scala 31:69:@23152.4]
  assign _T_3381 = _T_3351 ? _T_3363 : _T_3380; // @[Mux.scala 31:69:@23153.4]
  assign _T_3382 = _T_3350 ? _T_3361 : _T_3381; // @[Mux.scala 31:69:@23154.4]
  assign _T_3383 = _T_3349 ? _T_3359 : _T_3382; // @[Mux.scala 31:69:@23155.4]
  assign _T_3479 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@23284.4 package.scala 96:25:@23285.4]
  assign _T_3483 = _T_3479 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@23294.4]
  assign _T_3476 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@23276.4 package.scala 96:25:@23277.4]
  assign _T_3484 = _T_3476 ? Mem1D_19_io_output : _T_3483; // @[Mux.scala 31:69:@23295.4]
  assign _T_3473 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@23268.4 package.scala 96:25:@23269.4]
  assign _T_3485 = _T_3473 ? Mem1D_17_io_output : _T_3484; // @[Mux.scala 31:69:@23296.4]
  assign _T_3470 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@23260.4 package.scala 96:25:@23261.4]
  assign _T_3486 = _T_3470 ? Mem1D_15_io_output : _T_3485; // @[Mux.scala 31:69:@23297.4]
  assign _T_3467 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@23252.4 package.scala 96:25:@23253.4]
  assign _T_3487 = _T_3467 ? Mem1D_13_io_output : _T_3486; // @[Mux.scala 31:69:@23298.4]
  assign _T_3464 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@23244.4 package.scala 96:25:@23245.4]
  assign _T_3488 = _T_3464 ? Mem1D_11_io_output : _T_3487; // @[Mux.scala 31:69:@23299.4]
  assign _T_3461 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@23236.4 package.scala 96:25:@23237.4]
  assign _T_3489 = _T_3461 ? Mem1D_9_io_output : _T_3488; // @[Mux.scala 31:69:@23300.4]
  assign _T_3458 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@23228.4 package.scala 96:25:@23229.4]
  assign _T_3490 = _T_3458 ? Mem1D_7_io_output : _T_3489; // @[Mux.scala 31:69:@23301.4]
  assign _T_3455 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@23220.4 package.scala 96:25:@23221.4]
  assign _T_3491 = _T_3455 ? Mem1D_5_io_output : _T_3490; // @[Mux.scala 31:69:@23302.4]
  assign _T_3452 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@23212.4 package.scala 96:25:@23213.4]
  assign _T_3492 = _T_3452 ? Mem1D_3_io_output : _T_3491; // @[Mux.scala 31:69:@23303.4]
  assign _T_3449 = RetimeWrapper_io_out; // @[package.scala 96:25:@23204.4 package.scala 96:25:@23205.4]
  assign _T_3586 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@23428.4 package.scala 96:25:@23429.4]
  assign _T_3590 = _T_3586 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@23438.4]
  assign _T_3583 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@23420.4 package.scala 96:25:@23421.4]
  assign _T_3591 = _T_3583 ? Mem1D_18_io_output : _T_3590; // @[Mux.scala 31:69:@23439.4]
  assign _T_3580 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@23412.4 package.scala 96:25:@23413.4]
  assign _T_3592 = _T_3580 ? Mem1D_16_io_output : _T_3591; // @[Mux.scala 31:69:@23440.4]
  assign _T_3577 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@23404.4 package.scala 96:25:@23405.4]
  assign _T_3593 = _T_3577 ? Mem1D_14_io_output : _T_3592; // @[Mux.scala 31:69:@23441.4]
  assign _T_3574 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@23396.4 package.scala 96:25:@23397.4]
  assign _T_3594 = _T_3574 ? Mem1D_12_io_output : _T_3593; // @[Mux.scala 31:69:@23442.4]
  assign _T_3571 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@23388.4 package.scala 96:25:@23389.4]
  assign _T_3595 = _T_3571 ? Mem1D_10_io_output : _T_3594; // @[Mux.scala 31:69:@23443.4]
  assign _T_3568 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@23380.4 package.scala 96:25:@23381.4]
  assign _T_3596 = _T_3568 ? Mem1D_8_io_output : _T_3595; // @[Mux.scala 31:69:@23444.4]
  assign _T_3565 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@23372.4 package.scala 96:25:@23373.4]
  assign _T_3597 = _T_3565 ? Mem1D_6_io_output : _T_3596; // @[Mux.scala 31:69:@23445.4]
  assign _T_3562 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@23364.4 package.scala 96:25:@23365.4]
  assign _T_3598 = _T_3562 ? Mem1D_4_io_output : _T_3597; // @[Mux.scala 31:69:@23446.4]
  assign _T_3559 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@23356.4 package.scala 96:25:@23357.4]
  assign _T_3599 = _T_3559 ? Mem1D_2_io_output : _T_3598; // @[Mux.scala 31:69:@23447.4]
  assign _T_3556 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@23348.4 package.scala 96:25:@23349.4]
  assign _T_3693 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@23572.4 package.scala 96:25:@23573.4]
  assign _T_3697 = _T_3693 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@23582.4]
  assign _T_3690 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@23564.4 package.scala 96:25:@23565.4]
  assign _T_3698 = _T_3690 ? Mem1D_19_io_output : _T_3697; // @[Mux.scala 31:69:@23583.4]
  assign _T_3687 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@23556.4 package.scala 96:25:@23557.4]
  assign _T_3699 = _T_3687 ? Mem1D_17_io_output : _T_3698; // @[Mux.scala 31:69:@23584.4]
  assign _T_3684 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@23548.4 package.scala 96:25:@23549.4]
  assign _T_3700 = _T_3684 ? Mem1D_15_io_output : _T_3699; // @[Mux.scala 31:69:@23585.4]
  assign _T_3681 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@23540.4 package.scala 96:25:@23541.4]
  assign _T_3701 = _T_3681 ? Mem1D_13_io_output : _T_3700; // @[Mux.scala 31:69:@23586.4]
  assign _T_3678 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@23532.4 package.scala 96:25:@23533.4]
  assign _T_3702 = _T_3678 ? Mem1D_11_io_output : _T_3701; // @[Mux.scala 31:69:@23587.4]
  assign _T_3675 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@23524.4 package.scala 96:25:@23525.4]
  assign _T_3703 = _T_3675 ? Mem1D_9_io_output : _T_3702; // @[Mux.scala 31:69:@23588.4]
  assign _T_3672 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@23516.4 package.scala 96:25:@23517.4]
  assign _T_3704 = _T_3672 ? Mem1D_7_io_output : _T_3703; // @[Mux.scala 31:69:@23589.4]
  assign _T_3669 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@23508.4 package.scala 96:25:@23509.4]
  assign _T_3705 = _T_3669 ? Mem1D_5_io_output : _T_3704; // @[Mux.scala 31:69:@23590.4]
  assign _T_3666 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@23500.4 package.scala 96:25:@23501.4]
  assign _T_3706 = _T_3666 ? Mem1D_3_io_output : _T_3705; // @[Mux.scala 31:69:@23591.4]
  assign _T_3663 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@23492.4 package.scala 96:25:@23493.4]
  assign _T_3800 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@23716.4 package.scala 96:25:@23717.4]
  assign _T_3804 = _T_3800 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@23726.4]
  assign _T_3797 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@23708.4 package.scala 96:25:@23709.4]
  assign _T_3805 = _T_3797 ? Mem1D_18_io_output : _T_3804; // @[Mux.scala 31:69:@23727.4]
  assign _T_3794 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@23700.4 package.scala 96:25:@23701.4]
  assign _T_3806 = _T_3794 ? Mem1D_16_io_output : _T_3805; // @[Mux.scala 31:69:@23728.4]
  assign _T_3791 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@23692.4 package.scala 96:25:@23693.4]
  assign _T_3807 = _T_3791 ? Mem1D_14_io_output : _T_3806; // @[Mux.scala 31:69:@23729.4]
  assign _T_3788 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@23684.4 package.scala 96:25:@23685.4]
  assign _T_3808 = _T_3788 ? Mem1D_12_io_output : _T_3807; // @[Mux.scala 31:69:@23730.4]
  assign _T_3785 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@23676.4 package.scala 96:25:@23677.4]
  assign _T_3809 = _T_3785 ? Mem1D_10_io_output : _T_3808; // @[Mux.scala 31:69:@23731.4]
  assign _T_3782 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@23668.4 package.scala 96:25:@23669.4]
  assign _T_3810 = _T_3782 ? Mem1D_8_io_output : _T_3809; // @[Mux.scala 31:69:@23732.4]
  assign _T_3779 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@23660.4 package.scala 96:25:@23661.4]
  assign _T_3811 = _T_3779 ? Mem1D_6_io_output : _T_3810; // @[Mux.scala 31:69:@23733.4]
  assign _T_3776 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@23652.4 package.scala 96:25:@23653.4]
  assign _T_3812 = _T_3776 ? Mem1D_4_io_output : _T_3811; // @[Mux.scala 31:69:@23734.4]
  assign _T_3773 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@23644.4 package.scala 96:25:@23645.4]
  assign _T_3813 = _T_3773 ? Mem1D_2_io_output : _T_3812; // @[Mux.scala 31:69:@23735.4]
  assign _T_3770 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@23636.4 package.scala 96:25:@23637.4]
  assign _T_3907 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@23860.4 package.scala 96:25:@23861.4]
  assign _T_3911 = _T_3907 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@23870.4]
  assign _T_3904 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@23852.4 package.scala 96:25:@23853.4]
  assign _T_3912 = _T_3904 ? Mem1D_19_io_output : _T_3911; // @[Mux.scala 31:69:@23871.4]
  assign _T_3901 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@23844.4 package.scala 96:25:@23845.4]
  assign _T_3913 = _T_3901 ? Mem1D_17_io_output : _T_3912; // @[Mux.scala 31:69:@23872.4]
  assign _T_3898 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@23836.4 package.scala 96:25:@23837.4]
  assign _T_3914 = _T_3898 ? Mem1D_15_io_output : _T_3913; // @[Mux.scala 31:69:@23873.4]
  assign _T_3895 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@23828.4 package.scala 96:25:@23829.4]
  assign _T_3915 = _T_3895 ? Mem1D_13_io_output : _T_3914; // @[Mux.scala 31:69:@23874.4]
  assign _T_3892 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@23820.4 package.scala 96:25:@23821.4]
  assign _T_3916 = _T_3892 ? Mem1D_11_io_output : _T_3915; // @[Mux.scala 31:69:@23875.4]
  assign _T_3889 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@23812.4 package.scala 96:25:@23813.4]
  assign _T_3917 = _T_3889 ? Mem1D_9_io_output : _T_3916; // @[Mux.scala 31:69:@23876.4]
  assign _T_3886 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@23804.4 package.scala 96:25:@23805.4]
  assign _T_3918 = _T_3886 ? Mem1D_7_io_output : _T_3917; // @[Mux.scala 31:69:@23877.4]
  assign _T_3883 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@23796.4 package.scala 96:25:@23797.4]
  assign _T_3919 = _T_3883 ? Mem1D_5_io_output : _T_3918; // @[Mux.scala 31:69:@23878.4]
  assign _T_3880 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@23788.4 package.scala 96:25:@23789.4]
  assign _T_3920 = _T_3880 ? Mem1D_3_io_output : _T_3919; // @[Mux.scala 31:69:@23879.4]
  assign _T_3877 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@23780.4 package.scala 96:25:@23781.4]
  assign _T_4014 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@24004.4 package.scala 96:25:@24005.4]
  assign _T_4018 = _T_4014 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@24014.4]
  assign _T_4011 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@23996.4 package.scala 96:25:@23997.4]
  assign _T_4019 = _T_4011 ? Mem1D_19_io_output : _T_4018; // @[Mux.scala 31:69:@24015.4]
  assign _T_4008 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@23988.4 package.scala 96:25:@23989.4]
  assign _T_4020 = _T_4008 ? Mem1D_17_io_output : _T_4019; // @[Mux.scala 31:69:@24016.4]
  assign _T_4005 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@23980.4 package.scala 96:25:@23981.4]
  assign _T_4021 = _T_4005 ? Mem1D_15_io_output : _T_4020; // @[Mux.scala 31:69:@24017.4]
  assign _T_4002 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@23972.4 package.scala 96:25:@23973.4]
  assign _T_4022 = _T_4002 ? Mem1D_13_io_output : _T_4021; // @[Mux.scala 31:69:@24018.4]
  assign _T_3999 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@23964.4 package.scala 96:25:@23965.4]
  assign _T_4023 = _T_3999 ? Mem1D_11_io_output : _T_4022; // @[Mux.scala 31:69:@24019.4]
  assign _T_3996 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@23956.4 package.scala 96:25:@23957.4]
  assign _T_4024 = _T_3996 ? Mem1D_9_io_output : _T_4023; // @[Mux.scala 31:69:@24020.4]
  assign _T_3993 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@23948.4 package.scala 96:25:@23949.4]
  assign _T_4025 = _T_3993 ? Mem1D_7_io_output : _T_4024; // @[Mux.scala 31:69:@24021.4]
  assign _T_3990 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@23940.4 package.scala 96:25:@23941.4]
  assign _T_4026 = _T_3990 ? Mem1D_5_io_output : _T_4025; // @[Mux.scala 31:69:@24022.4]
  assign _T_3987 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@23932.4 package.scala 96:25:@23933.4]
  assign _T_4027 = _T_3987 ? Mem1D_3_io_output : _T_4026; // @[Mux.scala 31:69:@24023.4]
  assign _T_3984 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@23924.4 package.scala 96:25:@23925.4]
  assign _T_4121 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@24148.4 package.scala 96:25:@24149.4]
  assign _T_4125 = _T_4121 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@24158.4]
  assign _T_4118 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@24140.4 package.scala 96:25:@24141.4]
  assign _T_4126 = _T_4118 ? Mem1D_18_io_output : _T_4125; // @[Mux.scala 31:69:@24159.4]
  assign _T_4115 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@24132.4 package.scala 96:25:@24133.4]
  assign _T_4127 = _T_4115 ? Mem1D_16_io_output : _T_4126; // @[Mux.scala 31:69:@24160.4]
  assign _T_4112 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@24124.4 package.scala 96:25:@24125.4]
  assign _T_4128 = _T_4112 ? Mem1D_14_io_output : _T_4127; // @[Mux.scala 31:69:@24161.4]
  assign _T_4109 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@24116.4 package.scala 96:25:@24117.4]
  assign _T_4129 = _T_4109 ? Mem1D_12_io_output : _T_4128; // @[Mux.scala 31:69:@24162.4]
  assign _T_4106 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@24108.4 package.scala 96:25:@24109.4]
  assign _T_4130 = _T_4106 ? Mem1D_10_io_output : _T_4129; // @[Mux.scala 31:69:@24163.4]
  assign _T_4103 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@24100.4 package.scala 96:25:@24101.4]
  assign _T_4131 = _T_4103 ? Mem1D_8_io_output : _T_4130; // @[Mux.scala 31:69:@24164.4]
  assign _T_4100 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@24092.4 package.scala 96:25:@24093.4]
  assign _T_4132 = _T_4100 ? Mem1D_6_io_output : _T_4131; // @[Mux.scala 31:69:@24165.4]
  assign _T_4097 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@24084.4 package.scala 96:25:@24085.4]
  assign _T_4133 = _T_4097 ? Mem1D_4_io_output : _T_4132; // @[Mux.scala 31:69:@24166.4]
  assign _T_4094 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@24076.4 package.scala 96:25:@24077.4]
  assign _T_4134 = _T_4094 ? Mem1D_2_io_output : _T_4133; // @[Mux.scala 31:69:@24167.4]
  assign _T_4091 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@24068.4 package.scala 96:25:@24069.4]
  assign _T_4228 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@24292.4 package.scala 96:25:@24293.4]
  assign _T_4232 = _T_4228 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@24302.4]
  assign _T_4225 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@24284.4 package.scala 96:25:@24285.4]
  assign _T_4233 = _T_4225 ? Mem1D_19_io_output : _T_4232; // @[Mux.scala 31:69:@24303.4]
  assign _T_4222 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@24276.4 package.scala 96:25:@24277.4]
  assign _T_4234 = _T_4222 ? Mem1D_17_io_output : _T_4233; // @[Mux.scala 31:69:@24304.4]
  assign _T_4219 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@24268.4 package.scala 96:25:@24269.4]
  assign _T_4235 = _T_4219 ? Mem1D_15_io_output : _T_4234; // @[Mux.scala 31:69:@24305.4]
  assign _T_4216 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@24260.4 package.scala 96:25:@24261.4]
  assign _T_4236 = _T_4216 ? Mem1D_13_io_output : _T_4235; // @[Mux.scala 31:69:@24306.4]
  assign _T_4213 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@24252.4 package.scala 96:25:@24253.4]
  assign _T_4237 = _T_4213 ? Mem1D_11_io_output : _T_4236; // @[Mux.scala 31:69:@24307.4]
  assign _T_4210 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@24244.4 package.scala 96:25:@24245.4]
  assign _T_4238 = _T_4210 ? Mem1D_9_io_output : _T_4237; // @[Mux.scala 31:69:@24308.4]
  assign _T_4207 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@24236.4 package.scala 96:25:@24237.4]
  assign _T_4239 = _T_4207 ? Mem1D_7_io_output : _T_4238; // @[Mux.scala 31:69:@24309.4]
  assign _T_4204 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@24228.4 package.scala 96:25:@24229.4]
  assign _T_4240 = _T_4204 ? Mem1D_5_io_output : _T_4239; // @[Mux.scala 31:69:@24310.4]
  assign _T_4201 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@24220.4 package.scala 96:25:@24221.4]
  assign _T_4241 = _T_4201 ? Mem1D_3_io_output : _T_4240; // @[Mux.scala 31:69:@24311.4]
  assign _T_4198 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@24212.4 package.scala 96:25:@24213.4]
  assign _T_4335 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@24436.4 package.scala 96:25:@24437.4]
  assign _T_4339 = _T_4335 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@24446.4]
  assign _T_4332 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@24428.4 package.scala 96:25:@24429.4]
  assign _T_4340 = _T_4332 ? Mem1D_18_io_output : _T_4339; // @[Mux.scala 31:69:@24447.4]
  assign _T_4329 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@24420.4 package.scala 96:25:@24421.4]
  assign _T_4341 = _T_4329 ? Mem1D_16_io_output : _T_4340; // @[Mux.scala 31:69:@24448.4]
  assign _T_4326 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@24412.4 package.scala 96:25:@24413.4]
  assign _T_4342 = _T_4326 ? Mem1D_14_io_output : _T_4341; // @[Mux.scala 31:69:@24449.4]
  assign _T_4323 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@24404.4 package.scala 96:25:@24405.4]
  assign _T_4343 = _T_4323 ? Mem1D_12_io_output : _T_4342; // @[Mux.scala 31:69:@24450.4]
  assign _T_4320 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@24396.4 package.scala 96:25:@24397.4]
  assign _T_4344 = _T_4320 ? Mem1D_10_io_output : _T_4343; // @[Mux.scala 31:69:@24451.4]
  assign _T_4317 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@24388.4 package.scala 96:25:@24389.4]
  assign _T_4345 = _T_4317 ? Mem1D_8_io_output : _T_4344; // @[Mux.scala 31:69:@24452.4]
  assign _T_4314 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@24380.4 package.scala 96:25:@24381.4]
  assign _T_4346 = _T_4314 ? Mem1D_6_io_output : _T_4345; // @[Mux.scala 31:69:@24453.4]
  assign _T_4311 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@24372.4 package.scala 96:25:@24373.4]
  assign _T_4347 = _T_4311 ? Mem1D_4_io_output : _T_4346; // @[Mux.scala 31:69:@24454.4]
  assign _T_4308 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@24364.4 package.scala 96:25:@24365.4]
  assign _T_4348 = _T_4308 ? Mem1D_2_io_output : _T_4347; // @[Mux.scala 31:69:@24455.4]
  assign _T_4305 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@24356.4 package.scala 96:25:@24357.4]
  assign _T_4442 = RetimeWrapper_118_io_out; // @[package.scala 96:25:@24580.4 package.scala 96:25:@24581.4]
  assign _T_4446 = _T_4442 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@24590.4]
  assign _T_4439 = RetimeWrapper_117_io_out; // @[package.scala 96:25:@24572.4 package.scala 96:25:@24573.4]
  assign _T_4447 = _T_4439 ? Mem1D_19_io_output : _T_4446; // @[Mux.scala 31:69:@24591.4]
  assign _T_4436 = RetimeWrapper_116_io_out; // @[package.scala 96:25:@24564.4 package.scala 96:25:@24565.4]
  assign _T_4448 = _T_4436 ? Mem1D_17_io_output : _T_4447; // @[Mux.scala 31:69:@24592.4]
  assign _T_4433 = RetimeWrapper_115_io_out; // @[package.scala 96:25:@24556.4 package.scala 96:25:@24557.4]
  assign _T_4449 = _T_4433 ? Mem1D_15_io_output : _T_4448; // @[Mux.scala 31:69:@24593.4]
  assign _T_4430 = RetimeWrapper_114_io_out; // @[package.scala 96:25:@24548.4 package.scala 96:25:@24549.4]
  assign _T_4450 = _T_4430 ? Mem1D_13_io_output : _T_4449; // @[Mux.scala 31:69:@24594.4]
  assign _T_4427 = RetimeWrapper_113_io_out; // @[package.scala 96:25:@24540.4 package.scala 96:25:@24541.4]
  assign _T_4451 = _T_4427 ? Mem1D_11_io_output : _T_4450; // @[Mux.scala 31:69:@24595.4]
  assign _T_4424 = RetimeWrapper_112_io_out; // @[package.scala 96:25:@24532.4 package.scala 96:25:@24533.4]
  assign _T_4452 = _T_4424 ? Mem1D_9_io_output : _T_4451; // @[Mux.scala 31:69:@24596.4]
  assign _T_4421 = RetimeWrapper_111_io_out; // @[package.scala 96:25:@24524.4 package.scala 96:25:@24525.4]
  assign _T_4453 = _T_4421 ? Mem1D_7_io_output : _T_4452; // @[Mux.scala 31:69:@24597.4]
  assign _T_4418 = RetimeWrapper_110_io_out; // @[package.scala 96:25:@24516.4 package.scala 96:25:@24517.4]
  assign _T_4454 = _T_4418 ? Mem1D_5_io_output : _T_4453; // @[Mux.scala 31:69:@24598.4]
  assign _T_4415 = RetimeWrapper_109_io_out; // @[package.scala 96:25:@24508.4 package.scala 96:25:@24509.4]
  assign _T_4455 = _T_4415 ? Mem1D_3_io_output : _T_4454; // @[Mux.scala 31:69:@24599.4]
  assign _T_4412 = RetimeWrapper_108_io_out; // @[package.scala 96:25:@24500.4 package.scala 96:25:@24501.4]
  assign _T_4549 = RetimeWrapper_130_io_out; // @[package.scala 96:25:@24724.4 package.scala 96:25:@24725.4]
  assign _T_4553 = _T_4549 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@24734.4]
  assign _T_4546 = RetimeWrapper_129_io_out; // @[package.scala 96:25:@24716.4 package.scala 96:25:@24717.4]
  assign _T_4554 = _T_4546 ? Mem1D_18_io_output : _T_4553; // @[Mux.scala 31:69:@24735.4]
  assign _T_4543 = RetimeWrapper_128_io_out; // @[package.scala 96:25:@24708.4 package.scala 96:25:@24709.4]
  assign _T_4555 = _T_4543 ? Mem1D_16_io_output : _T_4554; // @[Mux.scala 31:69:@24736.4]
  assign _T_4540 = RetimeWrapper_127_io_out; // @[package.scala 96:25:@24700.4 package.scala 96:25:@24701.4]
  assign _T_4556 = _T_4540 ? Mem1D_14_io_output : _T_4555; // @[Mux.scala 31:69:@24737.4]
  assign _T_4537 = RetimeWrapper_126_io_out; // @[package.scala 96:25:@24692.4 package.scala 96:25:@24693.4]
  assign _T_4557 = _T_4537 ? Mem1D_12_io_output : _T_4556; // @[Mux.scala 31:69:@24738.4]
  assign _T_4534 = RetimeWrapper_125_io_out; // @[package.scala 96:25:@24684.4 package.scala 96:25:@24685.4]
  assign _T_4558 = _T_4534 ? Mem1D_10_io_output : _T_4557; // @[Mux.scala 31:69:@24739.4]
  assign _T_4531 = RetimeWrapper_124_io_out; // @[package.scala 96:25:@24676.4 package.scala 96:25:@24677.4]
  assign _T_4559 = _T_4531 ? Mem1D_8_io_output : _T_4558; // @[Mux.scala 31:69:@24740.4]
  assign _T_4528 = RetimeWrapper_123_io_out; // @[package.scala 96:25:@24668.4 package.scala 96:25:@24669.4]
  assign _T_4560 = _T_4528 ? Mem1D_6_io_output : _T_4559; // @[Mux.scala 31:69:@24741.4]
  assign _T_4525 = RetimeWrapper_122_io_out; // @[package.scala 96:25:@24660.4 package.scala 96:25:@24661.4]
  assign _T_4561 = _T_4525 ? Mem1D_4_io_output : _T_4560; // @[Mux.scala 31:69:@24742.4]
  assign _T_4522 = RetimeWrapper_121_io_out; // @[package.scala 96:25:@24652.4 package.scala 96:25:@24653.4]
  assign _T_4562 = _T_4522 ? Mem1D_2_io_output : _T_4561; // @[Mux.scala 31:69:@24743.4]
  assign _T_4519 = RetimeWrapper_120_io_out; // @[package.scala 96:25:@24644.4 package.scala 96:25:@24645.4]
  assign _T_4656 = RetimeWrapper_142_io_out; // @[package.scala 96:25:@24868.4 package.scala 96:25:@24869.4]
  assign _T_4660 = _T_4656 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@24878.4]
  assign _T_4653 = RetimeWrapper_141_io_out; // @[package.scala 96:25:@24860.4 package.scala 96:25:@24861.4]
  assign _T_4661 = _T_4653 ? Mem1D_19_io_output : _T_4660; // @[Mux.scala 31:69:@24879.4]
  assign _T_4650 = RetimeWrapper_140_io_out; // @[package.scala 96:25:@24852.4 package.scala 96:25:@24853.4]
  assign _T_4662 = _T_4650 ? Mem1D_17_io_output : _T_4661; // @[Mux.scala 31:69:@24880.4]
  assign _T_4647 = RetimeWrapper_139_io_out; // @[package.scala 96:25:@24844.4 package.scala 96:25:@24845.4]
  assign _T_4663 = _T_4647 ? Mem1D_15_io_output : _T_4662; // @[Mux.scala 31:69:@24881.4]
  assign _T_4644 = RetimeWrapper_138_io_out; // @[package.scala 96:25:@24836.4 package.scala 96:25:@24837.4]
  assign _T_4664 = _T_4644 ? Mem1D_13_io_output : _T_4663; // @[Mux.scala 31:69:@24882.4]
  assign _T_4641 = RetimeWrapper_137_io_out; // @[package.scala 96:25:@24828.4 package.scala 96:25:@24829.4]
  assign _T_4665 = _T_4641 ? Mem1D_11_io_output : _T_4664; // @[Mux.scala 31:69:@24883.4]
  assign _T_4638 = RetimeWrapper_136_io_out; // @[package.scala 96:25:@24820.4 package.scala 96:25:@24821.4]
  assign _T_4666 = _T_4638 ? Mem1D_9_io_output : _T_4665; // @[Mux.scala 31:69:@24884.4]
  assign _T_4635 = RetimeWrapper_135_io_out; // @[package.scala 96:25:@24812.4 package.scala 96:25:@24813.4]
  assign _T_4667 = _T_4635 ? Mem1D_7_io_output : _T_4666; // @[Mux.scala 31:69:@24885.4]
  assign _T_4632 = RetimeWrapper_134_io_out; // @[package.scala 96:25:@24804.4 package.scala 96:25:@24805.4]
  assign _T_4668 = _T_4632 ? Mem1D_5_io_output : _T_4667; // @[Mux.scala 31:69:@24886.4]
  assign _T_4629 = RetimeWrapper_133_io_out; // @[package.scala 96:25:@24796.4 package.scala 96:25:@24797.4]
  assign _T_4669 = _T_4629 ? Mem1D_3_io_output : _T_4668; // @[Mux.scala 31:69:@24887.4]
  assign _T_4626 = RetimeWrapper_132_io_out; // @[package.scala 96:25:@24788.4 package.scala 96:25:@24789.4]
  assign _T_4763 = RetimeWrapper_154_io_out; // @[package.scala 96:25:@25012.4 package.scala 96:25:@25013.4]
  assign _T_4767 = _T_4763 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@25022.4]
  assign _T_4760 = RetimeWrapper_153_io_out; // @[package.scala 96:25:@25004.4 package.scala 96:25:@25005.4]
  assign _T_4768 = _T_4760 ? Mem1D_18_io_output : _T_4767; // @[Mux.scala 31:69:@25023.4]
  assign _T_4757 = RetimeWrapper_152_io_out; // @[package.scala 96:25:@24996.4 package.scala 96:25:@24997.4]
  assign _T_4769 = _T_4757 ? Mem1D_16_io_output : _T_4768; // @[Mux.scala 31:69:@25024.4]
  assign _T_4754 = RetimeWrapper_151_io_out; // @[package.scala 96:25:@24988.4 package.scala 96:25:@24989.4]
  assign _T_4770 = _T_4754 ? Mem1D_14_io_output : _T_4769; // @[Mux.scala 31:69:@25025.4]
  assign _T_4751 = RetimeWrapper_150_io_out; // @[package.scala 96:25:@24980.4 package.scala 96:25:@24981.4]
  assign _T_4771 = _T_4751 ? Mem1D_12_io_output : _T_4770; // @[Mux.scala 31:69:@25026.4]
  assign _T_4748 = RetimeWrapper_149_io_out; // @[package.scala 96:25:@24972.4 package.scala 96:25:@24973.4]
  assign _T_4772 = _T_4748 ? Mem1D_10_io_output : _T_4771; // @[Mux.scala 31:69:@25027.4]
  assign _T_4745 = RetimeWrapper_148_io_out; // @[package.scala 96:25:@24964.4 package.scala 96:25:@24965.4]
  assign _T_4773 = _T_4745 ? Mem1D_8_io_output : _T_4772; // @[Mux.scala 31:69:@25028.4]
  assign _T_4742 = RetimeWrapper_147_io_out; // @[package.scala 96:25:@24956.4 package.scala 96:25:@24957.4]
  assign _T_4774 = _T_4742 ? Mem1D_6_io_output : _T_4773; // @[Mux.scala 31:69:@25029.4]
  assign _T_4739 = RetimeWrapper_146_io_out; // @[package.scala 96:25:@24948.4 package.scala 96:25:@24949.4]
  assign _T_4775 = _T_4739 ? Mem1D_4_io_output : _T_4774; // @[Mux.scala 31:69:@25030.4]
  assign _T_4736 = RetimeWrapper_145_io_out; // @[package.scala 96:25:@24940.4 package.scala 96:25:@24941.4]
  assign _T_4776 = _T_4736 ? Mem1D_2_io_output : _T_4775; // @[Mux.scala 31:69:@25031.4]
  assign _T_4733 = RetimeWrapper_144_io_out; // @[package.scala 96:25:@24932.4 package.scala 96:25:@24933.4]
  assign _T_4870 = RetimeWrapper_166_io_out; // @[package.scala 96:25:@25156.4 package.scala 96:25:@25157.4]
  assign _T_4874 = _T_4870 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@25166.4]
  assign _T_4867 = RetimeWrapper_165_io_out; // @[package.scala 96:25:@25148.4 package.scala 96:25:@25149.4]
  assign _T_4875 = _T_4867 ? Mem1D_19_io_output : _T_4874; // @[Mux.scala 31:69:@25167.4]
  assign _T_4864 = RetimeWrapper_164_io_out; // @[package.scala 96:25:@25140.4 package.scala 96:25:@25141.4]
  assign _T_4876 = _T_4864 ? Mem1D_17_io_output : _T_4875; // @[Mux.scala 31:69:@25168.4]
  assign _T_4861 = RetimeWrapper_163_io_out; // @[package.scala 96:25:@25132.4 package.scala 96:25:@25133.4]
  assign _T_4877 = _T_4861 ? Mem1D_15_io_output : _T_4876; // @[Mux.scala 31:69:@25169.4]
  assign _T_4858 = RetimeWrapper_162_io_out; // @[package.scala 96:25:@25124.4 package.scala 96:25:@25125.4]
  assign _T_4878 = _T_4858 ? Mem1D_13_io_output : _T_4877; // @[Mux.scala 31:69:@25170.4]
  assign _T_4855 = RetimeWrapper_161_io_out; // @[package.scala 96:25:@25116.4 package.scala 96:25:@25117.4]
  assign _T_4879 = _T_4855 ? Mem1D_11_io_output : _T_4878; // @[Mux.scala 31:69:@25171.4]
  assign _T_4852 = RetimeWrapper_160_io_out; // @[package.scala 96:25:@25108.4 package.scala 96:25:@25109.4]
  assign _T_4880 = _T_4852 ? Mem1D_9_io_output : _T_4879; // @[Mux.scala 31:69:@25172.4]
  assign _T_4849 = RetimeWrapper_159_io_out; // @[package.scala 96:25:@25100.4 package.scala 96:25:@25101.4]
  assign _T_4881 = _T_4849 ? Mem1D_7_io_output : _T_4880; // @[Mux.scala 31:69:@25173.4]
  assign _T_4846 = RetimeWrapper_158_io_out; // @[package.scala 96:25:@25092.4 package.scala 96:25:@25093.4]
  assign _T_4882 = _T_4846 ? Mem1D_5_io_output : _T_4881; // @[Mux.scala 31:69:@25174.4]
  assign _T_4843 = RetimeWrapper_157_io_out; // @[package.scala 96:25:@25084.4 package.scala 96:25:@25085.4]
  assign _T_4883 = _T_4843 ? Mem1D_3_io_output : _T_4882; // @[Mux.scala 31:69:@25175.4]
  assign _T_4840 = RetimeWrapper_156_io_out; // @[package.scala 96:25:@25076.4 package.scala 96:25:@25077.4]
  assign _T_4977 = RetimeWrapper_178_io_out; // @[package.scala 96:25:@25300.4 package.scala 96:25:@25301.4]
  assign _T_4981 = _T_4977 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@25310.4]
  assign _T_4974 = RetimeWrapper_177_io_out; // @[package.scala 96:25:@25292.4 package.scala 96:25:@25293.4]
  assign _T_4982 = _T_4974 ? Mem1D_19_io_output : _T_4981; // @[Mux.scala 31:69:@25311.4]
  assign _T_4971 = RetimeWrapper_176_io_out; // @[package.scala 96:25:@25284.4 package.scala 96:25:@25285.4]
  assign _T_4983 = _T_4971 ? Mem1D_17_io_output : _T_4982; // @[Mux.scala 31:69:@25312.4]
  assign _T_4968 = RetimeWrapper_175_io_out; // @[package.scala 96:25:@25276.4 package.scala 96:25:@25277.4]
  assign _T_4984 = _T_4968 ? Mem1D_15_io_output : _T_4983; // @[Mux.scala 31:69:@25313.4]
  assign _T_4965 = RetimeWrapper_174_io_out; // @[package.scala 96:25:@25268.4 package.scala 96:25:@25269.4]
  assign _T_4985 = _T_4965 ? Mem1D_13_io_output : _T_4984; // @[Mux.scala 31:69:@25314.4]
  assign _T_4962 = RetimeWrapper_173_io_out; // @[package.scala 96:25:@25260.4 package.scala 96:25:@25261.4]
  assign _T_4986 = _T_4962 ? Mem1D_11_io_output : _T_4985; // @[Mux.scala 31:69:@25315.4]
  assign _T_4959 = RetimeWrapper_172_io_out; // @[package.scala 96:25:@25252.4 package.scala 96:25:@25253.4]
  assign _T_4987 = _T_4959 ? Mem1D_9_io_output : _T_4986; // @[Mux.scala 31:69:@25316.4]
  assign _T_4956 = RetimeWrapper_171_io_out; // @[package.scala 96:25:@25244.4 package.scala 96:25:@25245.4]
  assign _T_4988 = _T_4956 ? Mem1D_7_io_output : _T_4987; // @[Mux.scala 31:69:@25317.4]
  assign _T_4953 = RetimeWrapper_170_io_out; // @[package.scala 96:25:@25236.4 package.scala 96:25:@25237.4]
  assign _T_4989 = _T_4953 ? Mem1D_5_io_output : _T_4988; // @[Mux.scala 31:69:@25318.4]
  assign _T_4950 = RetimeWrapper_169_io_out; // @[package.scala 96:25:@25228.4 package.scala 96:25:@25229.4]
  assign _T_4990 = _T_4950 ? Mem1D_3_io_output : _T_4989; // @[Mux.scala 31:69:@25319.4]
  assign _T_4947 = RetimeWrapper_168_io_out; // @[package.scala 96:25:@25220.4 package.scala 96:25:@25221.4]
  assign _T_5084 = RetimeWrapper_190_io_out; // @[package.scala 96:25:@25444.4 package.scala 96:25:@25445.4]
  assign _T_5088 = _T_5084 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@25454.4]
  assign _T_5081 = RetimeWrapper_189_io_out; // @[package.scala 96:25:@25436.4 package.scala 96:25:@25437.4]
  assign _T_5089 = _T_5081 ? Mem1D_18_io_output : _T_5088; // @[Mux.scala 31:69:@25455.4]
  assign _T_5078 = RetimeWrapper_188_io_out; // @[package.scala 96:25:@25428.4 package.scala 96:25:@25429.4]
  assign _T_5090 = _T_5078 ? Mem1D_16_io_output : _T_5089; // @[Mux.scala 31:69:@25456.4]
  assign _T_5075 = RetimeWrapper_187_io_out; // @[package.scala 96:25:@25420.4 package.scala 96:25:@25421.4]
  assign _T_5091 = _T_5075 ? Mem1D_14_io_output : _T_5090; // @[Mux.scala 31:69:@25457.4]
  assign _T_5072 = RetimeWrapper_186_io_out; // @[package.scala 96:25:@25412.4 package.scala 96:25:@25413.4]
  assign _T_5092 = _T_5072 ? Mem1D_12_io_output : _T_5091; // @[Mux.scala 31:69:@25458.4]
  assign _T_5069 = RetimeWrapper_185_io_out; // @[package.scala 96:25:@25404.4 package.scala 96:25:@25405.4]
  assign _T_5093 = _T_5069 ? Mem1D_10_io_output : _T_5092; // @[Mux.scala 31:69:@25459.4]
  assign _T_5066 = RetimeWrapper_184_io_out; // @[package.scala 96:25:@25396.4 package.scala 96:25:@25397.4]
  assign _T_5094 = _T_5066 ? Mem1D_8_io_output : _T_5093; // @[Mux.scala 31:69:@25460.4]
  assign _T_5063 = RetimeWrapper_183_io_out; // @[package.scala 96:25:@25388.4 package.scala 96:25:@25389.4]
  assign _T_5095 = _T_5063 ? Mem1D_6_io_output : _T_5094; // @[Mux.scala 31:69:@25461.4]
  assign _T_5060 = RetimeWrapper_182_io_out; // @[package.scala 96:25:@25380.4 package.scala 96:25:@25381.4]
  assign _T_5096 = _T_5060 ? Mem1D_4_io_output : _T_5095; // @[Mux.scala 31:69:@25462.4]
  assign _T_5057 = RetimeWrapper_181_io_out; // @[package.scala 96:25:@25372.4 package.scala 96:25:@25373.4]
  assign _T_5097 = _T_5057 ? Mem1D_2_io_output : _T_5096; // @[Mux.scala 31:69:@25463.4]
  assign _T_5054 = RetimeWrapper_180_io_out; // @[package.scala 96:25:@25364.4 package.scala 96:25:@25365.4]
  assign _T_5191 = RetimeWrapper_202_io_out; // @[package.scala 96:25:@25588.4 package.scala 96:25:@25589.4]
  assign _T_5195 = _T_5191 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@25598.4]
  assign _T_5188 = RetimeWrapper_201_io_out; // @[package.scala 96:25:@25580.4 package.scala 96:25:@25581.4]
  assign _T_5196 = _T_5188 ? Mem1D_18_io_output : _T_5195; // @[Mux.scala 31:69:@25599.4]
  assign _T_5185 = RetimeWrapper_200_io_out; // @[package.scala 96:25:@25572.4 package.scala 96:25:@25573.4]
  assign _T_5197 = _T_5185 ? Mem1D_16_io_output : _T_5196; // @[Mux.scala 31:69:@25600.4]
  assign _T_5182 = RetimeWrapper_199_io_out; // @[package.scala 96:25:@25564.4 package.scala 96:25:@25565.4]
  assign _T_5198 = _T_5182 ? Mem1D_14_io_output : _T_5197; // @[Mux.scala 31:69:@25601.4]
  assign _T_5179 = RetimeWrapper_198_io_out; // @[package.scala 96:25:@25556.4 package.scala 96:25:@25557.4]
  assign _T_5199 = _T_5179 ? Mem1D_12_io_output : _T_5198; // @[Mux.scala 31:69:@25602.4]
  assign _T_5176 = RetimeWrapper_197_io_out; // @[package.scala 96:25:@25548.4 package.scala 96:25:@25549.4]
  assign _T_5200 = _T_5176 ? Mem1D_10_io_output : _T_5199; // @[Mux.scala 31:69:@25603.4]
  assign _T_5173 = RetimeWrapper_196_io_out; // @[package.scala 96:25:@25540.4 package.scala 96:25:@25541.4]
  assign _T_5201 = _T_5173 ? Mem1D_8_io_output : _T_5200; // @[Mux.scala 31:69:@25604.4]
  assign _T_5170 = RetimeWrapper_195_io_out; // @[package.scala 96:25:@25532.4 package.scala 96:25:@25533.4]
  assign _T_5202 = _T_5170 ? Mem1D_6_io_output : _T_5201; // @[Mux.scala 31:69:@25605.4]
  assign _T_5167 = RetimeWrapper_194_io_out; // @[package.scala 96:25:@25524.4 package.scala 96:25:@25525.4]
  assign _T_5203 = _T_5167 ? Mem1D_4_io_output : _T_5202; // @[Mux.scala 31:69:@25606.4]
  assign _T_5164 = RetimeWrapper_193_io_out; // @[package.scala 96:25:@25516.4 package.scala 96:25:@25517.4]
  assign _T_5204 = _T_5164 ? Mem1D_2_io_output : _T_5203; // @[Mux.scala 31:69:@25607.4]
  assign _T_5161 = RetimeWrapper_192_io_out; // @[package.scala 96:25:@25508.4 package.scala 96:25:@25509.4]
  assign _T_5298 = RetimeWrapper_214_io_out; // @[package.scala 96:25:@25732.4 package.scala 96:25:@25733.4]
  assign _T_5302 = _T_5298 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@25742.4]
  assign _T_5295 = RetimeWrapper_213_io_out; // @[package.scala 96:25:@25724.4 package.scala 96:25:@25725.4]
  assign _T_5303 = _T_5295 ? Mem1D_18_io_output : _T_5302; // @[Mux.scala 31:69:@25743.4]
  assign _T_5292 = RetimeWrapper_212_io_out; // @[package.scala 96:25:@25716.4 package.scala 96:25:@25717.4]
  assign _T_5304 = _T_5292 ? Mem1D_16_io_output : _T_5303; // @[Mux.scala 31:69:@25744.4]
  assign _T_5289 = RetimeWrapper_211_io_out; // @[package.scala 96:25:@25708.4 package.scala 96:25:@25709.4]
  assign _T_5305 = _T_5289 ? Mem1D_14_io_output : _T_5304; // @[Mux.scala 31:69:@25745.4]
  assign _T_5286 = RetimeWrapper_210_io_out; // @[package.scala 96:25:@25700.4 package.scala 96:25:@25701.4]
  assign _T_5306 = _T_5286 ? Mem1D_12_io_output : _T_5305; // @[Mux.scala 31:69:@25746.4]
  assign _T_5283 = RetimeWrapper_209_io_out; // @[package.scala 96:25:@25692.4 package.scala 96:25:@25693.4]
  assign _T_5307 = _T_5283 ? Mem1D_10_io_output : _T_5306; // @[Mux.scala 31:69:@25747.4]
  assign _T_5280 = RetimeWrapper_208_io_out; // @[package.scala 96:25:@25684.4 package.scala 96:25:@25685.4]
  assign _T_5308 = _T_5280 ? Mem1D_8_io_output : _T_5307; // @[Mux.scala 31:69:@25748.4]
  assign _T_5277 = RetimeWrapper_207_io_out; // @[package.scala 96:25:@25676.4 package.scala 96:25:@25677.4]
  assign _T_5309 = _T_5277 ? Mem1D_6_io_output : _T_5308; // @[Mux.scala 31:69:@25749.4]
  assign _T_5274 = RetimeWrapper_206_io_out; // @[package.scala 96:25:@25668.4 package.scala 96:25:@25669.4]
  assign _T_5310 = _T_5274 ? Mem1D_4_io_output : _T_5309; // @[Mux.scala 31:69:@25750.4]
  assign _T_5271 = RetimeWrapper_205_io_out; // @[package.scala 96:25:@25660.4 package.scala 96:25:@25661.4]
  assign _T_5311 = _T_5271 ? Mem1D_2_io_output : _T_5310; // @[Mux.scala 31:69:@25751.4]
  assign _T_5268 = RetimeWrapper_204_io_out; // @[package.scala 96:25:@25652.4 package.scala 96:25:@25653.4]
  assign io_rPort_17_output_0 = _T_5268 ? Mem1D_io_output : _T_5311; // @[MemPrimitives.scala 152:13:@25753.4]
  assign io_rPort_16_output_0 = _T_5161 ? Mem1D_io_output : _T_5204; // @[MemPrimitives.scala 152:13:@25609.4]
  assign io_rPort_15_output_0 = _T_5054 ? Mem1D_io_output : _T_5097; // @[MemPrimitives.scala 152:13:@25465.4]
  assign io_rPort_14_output_0 = _T_4947 ? Mem1D_1_io_output : _T_4990; // @[MemPrimitives.scala 152:13:@25321.4]
  assign io_rPort_13_output_0 = _T_4840 ? Mem1D_1_io_output : _T_4883; // @[MemPrimitives.scala 152:13:@25177.4]
  assign io_rPort_12_output_0 = _T_4733 ? Mem1D_io_output : _T_4776; // @[MemPrimitives.scala 152:13:@25033.4]
  assign io_rPort_11_output_0 = _T_4626 ? Mem1D_1_io_output : _T_4669; // @[MemPrimitives.scala 152:13:@24889.4]
  assign io_rPort_10_output_0 = _T_4519 ? Mem1D_io_output : _T_4562; // @[MemPrimitives.scala 152:13:@24745.4]
  assign io_rPort_9_output_0 = _T_4412 ? Mem1D_1_io_output : _T_4455; // @[MemPrimitives.scala 152:13:@24601.4]
  assign io_rPort_8_output_0 = _T_4305 ? Mem1D_io_output : _T_4348; // @[MemPrimitives.scala 152:13:@24457.4]
  assign io_rPort_7_output_0 = _T_4198 ? Mem1D_1_io_output : _T_4241; // @[MemPrimitives.scala 152:13:@24313.4]
  assign io_rPort_6_output_0 = _T_4091 ? Mem1D_io_output : _T_4134; // @[MemPrimitives.scala 152:13:@24169.4]
  assign io_rPort_5_output_0 = _T_3984 ? Mem1D_1_io_output : _T_4027; // @[MemPrimitives.scala 152:13:@24025.4]
  assign io_rPort_4_output_0 = _T_3877 ? Mem1D_1_io_output : _T_3920; // @[MemPrimitives.scala 152:13:@23881.4]
  assign io_rPort_3_output_0 = _T_3770 ? Mem1D_io_output : _T_3813; // @[MemPrimitives.scala 152:13:@23737.4]
  assign io_rPort_2_output_0 = _T_3663 ? Mem1D_1_io_output : _T_3706; // @[MemPrimitives.scala 152:13:@23593.4]
  assign io_rPort_1_output_0 = _T_3556 ? Mem1D_io_output : _T_3599; // @[MemPrimitives.scala 152:13:@23449.4]
  assign io_rPort_0_output_0 = _T_3449 ? Mem1D_1_io_output : _T_3492; // @[MemPrimitives.scala 152:13:@23305.4]
  assign Mem1D_clock = clock; // @[:@20187.4]
  assign Mem1D_reset = reset; // @[:@20188.4]
  assign Mem1D_io_r_ofs_0 = _T_1267[8:0]; // @[MemPrimitives.scala 131:28:@21112.4]
  assign Mem1D_io_r_backpressure = _T_1267[9]; // @[MemPrimitives.scala 132:32:@21113.4]
  assign Mem1D_io_w_ofs_0 = _T_715[8:0]; // @[MemPrimitives.scala 94:28:@20586.4]
  assign Mem1D_io_w_data_0 = _T_715[40:9]; // @[MemPrimitives.scala 95:29:@20587.4]
  assign Mem1D_io_w_en_0 = _T_715[41]; // @[MemPrimitives.scala 96:27:@20588.4]
  assign Mem1D_1_clock = clock; // @[:@20203.4]
  assign Mem1D_1_reset = reset; // @[:@20204.4]
  assign Mem1D_1_io_r_ofs_0 = _T_1359[8:0]; // @[MemPrimitives.scala 131:28:@21201.4]
  assign Mem1D_1_io_r_backpressure = _T_1359[9]; // @[MemPrimitives.scala 132:32:@21202.4]
  assign Mem1D_1_io_w_ofs_0 = _T_735[8:0]; // @[MemPrimitives.scala 94:28:@20605.4]
  assign Mem1D_1_io_w_data_0 = _T_735[40:9]; // @[MemPrimitives.scala 95:29:@20606.4]
  assign Mem1D_1_io_w_en_0 = _T_735[41]; // @[MemPrimitives.scala 96:27:@20607.4]
  assign Mem1D_2_clock = clock; // @[:@20219.4]
  assign Mem1D_2_reset = reset; // @[:@20220.4]
  assign Mem1D_2_io_r_ofs_0 = _T_1451[8:0]; // @[MemPrimitives.scala 131:28:@21290.4]
  assign Mem1D_2_io_r_backpressure = _T_1451[9]; // @[MemPrimitives.scala 132:32:@21291.4]
  assign Mem1D_2_io_w_ofs_0 = _T_755[8:0]; // @[MemPrimitives.scala 94:28:@20624.4]
  assign Mem1D_2_io_w_data_0 = _T_755[40:9]; // @[MemPrimitives.scala 95:29:@20625.4]
  assign Mem1D_2_io_w_en_0 = _T_755[41]; // @[MemPrimitives.scala 96:27:@20626.4]
  assign Mem1D_3_clock = clock; // @[:@20235.4]
  assign Mem1D_3_reset = reset; // @[:@20236.4]
  assign Mem1D_3_io_r_ofs_0 = _T_1543[8:0]; // @[MemPrimitives.scala 131:28:@21379.4]
  assign Mem1D_3_io_r_backpressure = _T_1543[9]; // @[MemPrimitives.scala 132:32:@21380.4]
  assign Mem1D_3_io_w_ofs_0 = _T_775[8:0]; // @[MemPrimitives.scala 94:28:@20643.4]
  assign Mem1D_3_io_w_data_0 = _T_775[40:9]; // @[MemPrimitives.scala 95:29:@20644.4]
  assign Mem1D_3_io_w_en_0 = _T_775[41]; // @[MemPrimitives.scala 96:27:@20645.4]
  assign Mem1D_4_clock = clock; // @[:@20251.4]
  assign Mem1D_4_reset = reset; // @[:@20252.4]
  assign Mem1D_4_io_r_ofs_0 = _T_1635[8:0]; // @[MemPrimitives.scala 131:28:@21468.4]
  assign Mem1D_4_io_r_backpressure = _T_1635[9]; // @[MemPrimitives.scala 132:32:@21469.4]
  assign Mem1D_4_io_w_ofs_0 = _T_795[8:0]; // @[MemPrimitives.scala 94:28:@20662.4]
  assign Mem1D_4_io_w_data_0 = _T_795[40:9]; // @[MemPrimitives.scala 95:29:@20663.4]
  assign Mem1D_4_io_w_en_0 = _T_795[41]; // @[MemPrimitives.scala 96:27:@20664.4]
  assign Mem1D_5_clock = clock; // @[:@20267.4]
  assign Mem1D_5_reset = reset; // @[:@20268.4]
  assign Mem1D_5_io_r_ofs_0 = _T_1727[8:0]; // @[MemPrimitives.scala 131:28:@21557.4]
  assign Mem1D_5_io_r_backpressure = _T_1727[9]; // @[MemPrimitives.scala 132:32:@21558.4]
  assign Mem1D_5_io_w_ofs_0 = _T_815[8:0]; // @[MemPrimitives.scala 94:28:@20681.4]
  assign Mem1D_5_io_w_data_0 = _T_815[40:9]; // @[MemPrimitives.scala 95:29:@20682.4]
  assign Mem1D_5_io_w_en_0 = _T_815[41]; // @[MemPrimitives.scala 96:27:@20683.4]
  assign Mem1D_6_clock = clock; // @[:@20283.4]
  assign Mem1D_6_reset = reset; // @[:@20284.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1819[8:0]; // @[MemPrimitives.scala 131:28:@21646.4]
  assign Mem1D_6_io_r_backpressure = _T_1819[9]; // @[MemPrimitives.scala 132:32:@21647.4]
  assign Mem1D_6_io_w_ofs_0 = _T_835[8:0]; // @[MemPrimitives.scala 94:28:@20700.4]
  assign Mem1D_6_io_w_data_0 = _T_835[40:9]; // @[MemPrimitives.scala 95:29:@20701.4]
  assign Mem1D_6_io_w_en_0 = _T_835[41]; // @[MemPrimitives.scala 96:27:@20702.4]
  assign Mem1D_7_clock = clock; // @[:@20299.4]
  assign Mem1D_7_reset = reset; // @[:@20300.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1911[8:0]; // @[MemPrimitives.scala 131:28:@21735.4]
  assign Mem1D_7_io_r_backpressure = _T_1911[9]; // @[MemPrimitives.scala 132:32:@21736.4]
  assign Mem1D_7_io_w_ofs_0 = _T_855[8:0]; // @[MemPrimitives.scala 94:28:@20719.4]
  assign Mem1D_7_io_w_data_0 = _T_855[40:9]; // @[MemPrimitives.scala 95:29:@20720.4]
  assign Mem1D_7_io_w_en_0 = _T_855[41]; // @[MemPrimitives.scala 96:27:@20721.4]
  assign Mem1D_8_clock = clock; // @[:@20315.4]
  assign Mem1D_8_reset = reset; // @[:@20316.4]
  assign Mem1D_8_io_r_ofs_0 = _T_2003[8:0]; // @[MemPrimitives.scala 131:28:@21824.4]
  assign Mem1D_8_io_r_backpressure = _T_2003[9]; // @[MemPrimitives.scala 132:32:@21825.4]
  assign Mem1D_8_io_w_ofs_0 = _T_875[8:0]; // @[MemPrimitives.scala 94:28:@20738.4]
  assign Mem1D_8_io_w_data_0 = _T_875[40:9]; // @[MemPrimitives.scala 95:29:@20739.4]
  assign Mem1D_8_io_w_en_0 = _T_875[41]; // @[MemPrimitives.scala 96:27:@20740.4]
  assign Mem1D_9_clock = clock; // @[:@20331.4]
  assign Mem1D_9_reset = reset; // @[:@20332.4]
  assign Mem1D_9_io_r_ofs_0 = _T_2095[8:0]; // @[MemPrimitives.scala 131:28:@21913.4]
  assign Mem1D_9_io_r_backpressure = _T_2095[9]; // @[MemPrimitives.scala 132:32:@21914.4]
  assign Mem1D_9_io_w_ofs_0 = _T_895[8:0]; // @[MemPrimitives.scala 94:28:@20757.4]
  assign Mem1D_9_io_w_data_0 = _T_895[40:9]; // @[MemPrimitives.scala 95:29:@20758.4]
  assign Mem1D_9_io_w_en_0 = _T_895[41]; // @[MemPrimitives.scala 96:27:@20759.4]
  assign Mem1D_10_clock = clock; // @[:@20347.4]
  assign Mem1D_10_reset = reset; // @[:@20348.4]
  assign Mem1D_10_io_r_ofs_0 = _T_2187[8:0]; // @[MemPrimitives.scala 131:28:@22002.4]
  assign Mem1D_10_io_r_backpressure = _T_2187[9]; // @[MemPrimitives.scala 132:32:@22003.4]
  assign Mem1D_10_io_w_ofs_0 = _T_915[8:0]; // @[MemPrimitives.scala 94:28:@20776.4]
  assign Mem1D_10_io_w_data_0 = _T_915[40:9]; // @[MemPrimitives.scala 95:29:@20777.4]
  assign Mem1D_10_io_w_en_0 = _T_915[41]; // @[MemPrimitives.scala 96:27:@20778.4]
  assign Mem1D_11_clock = clock; // @[:@20363.4]
  assign Mem1D_11_reset = reset; // @[:@20364.4]
  assign Mem1D_11_io_r_ofs_0 = _T_2279[8:0]; // @[MemPrimitives.scala 131:28:@22091.4]
  assign Mem1D_11_io_r_backpressure = _T_2279[9]; // @[MemPrimitives.scala 132:32:@22092.4]
  assign Mem1D_11_io_w_ofs_0 = _T_935[8:0]; // @[MemPrimitives.scala 94:28:@20795.4]
  assign Mem1D_11_io_w_data_0 = _T_935[40:9]; // @[MemPrimitives.scala 95:29:@20796.4]
  assign Mem1D_11_io_w_en_0 = _T_935[41]; // @[MemPrimitives.scala 96:27:@20797.4]
  assign Mem1D_12_clock = clock; // @[:@20379.4]
  assign Mem1D_12_reset = reset; // @[:@20380.4]
  assign Mem1D_12_io_r_ofs_0 = _T_2371[8:0]; // @[MemPrimitives.scala 131:28:@22180.4]
  assign Mem1D_12_io_r_backpressure = _T_2371[9]; // @[MemPrimitives.scala 132:32:@22181.4]
  assign Mem1D_12_io_w_ofs_0 = _T_955[8:0]; // @[MemPrimitives.scala 94:28:@20814.4]
  assign Mem1D_12_io_w_data_0 = _T_955[40:9]; // @[MemPrimitives.scala 95:29:@20815.4]
  assign Mem1D_12_io_w_en_0 = _T_955[41]; // @[MemPrimitives.scala 96:27:@20816.4]
  assign Mem1D_13_clock = clock; // @[:@20395.4]
  assign Mem1D_13_reset = reset; // @[:@20396.4]
  assign Mem1D_13_io_r_ofs_0 = _T_2463[8:0]; // @[MemPrimitives.scala 131:28:@22269.4]
  assign Mem1D_13_io_r_backpressure = _T_2463[9]; // @[MemPrimitives.scala 132:32:@22270.4]
  assign Mem1D_13_io_w_ofs_0 = _T_975[8:0]; // @[MemPrimitives.scala 94:28:@20833.4]
  assign Mem1D_13_io_w_data_0 = _T_975[40:9]; // @[MemPrimitives.scala 95:29:@20834.4]
  assign Mem1D_13_io_w_en_0 = _T_975[41]; // @[MemPrimitives.scala 96:27:@20835.4]
  assign Mem1D_14_clock = clock; // @[:@20411.4]
  assign Mem1D_14_reset = reset; // @[:@20412.4]
  assign Mem1D_14_io_r_ofs_0 = _T_2555[8:0]; // @[MemPrimitives.scala 131:28:@22358.4]
  assign Mem1D_14_io_r_backpressure = _T_2555[9]; // @[MemPrimitives.scala 132:32:@22359.4]
  assign Mem1D_14_io_w_ofs_0 = _T_995[8:0]; // @[MemPrimitives.scala 94:28:@20852.4]
  assign Mem1D_14_io_w_data_0 = _T_995[40:9]; // @[MemPrimitives.scala 95:29:@20853.4]
  assign Mem1D_14_io_w_en_0 = _T_995[41]; // @[MemPrimitives.scala 96:27:@20854.4]
  assign Mem1D_15_clock = clock; // @[:@20427.4]
  assign Mem1D_15_reset = reset; // @[:@20428.4]
  assign Mem1D_15_io_r_ofs_0 = _T_2647[8:0]; // @[MemPrimitives.scala 131:28:@22447.4]
  assign Mem1D_15_io_r_backpressure = _T_2647[9]; // @[MemPrimitives.scala 132:32:@22448.4]
  assign Mem1D_15_io_w_ofs_0 = _T_1015[8:0]; // @[MemPrimitives.scala 94:28:@20871.4]
  assign Mem1D_15_io_w_data_0 = _T_1015[40:9]; // @[MemPrimitives.scala 95:29:@20872.4]
  assign Mem1D_15_io_w_en_0 = _T_1015[41]; // @[MemPrimitives.scala 96:27:@20873.4]
  assign Mem1D_16_clock = clock; // @[:@20443.4]
  assign Mem1D_16_reset = reset; // @[:@20444.4]
  assign Mem1D_16_io_r_ofs_0 = _T_2739[8:0]; // @[MemPrimitives.scala 131:28:@22536.4]
  assign Mem1D_16_io_r_backpressure = _T_2739[9]; // @[MemPrimitives.scala 132:32:@22537.4]
  assign Mem1D_16_io_w_ofs_0 = _T_1035[8:0]; // @[MemPrimitives.scala 94:28:@20890.4]
  assign Mem1D_16_io_w_data_0 = _T_1035[40:9]; // @[MemPrimitives.scala 95:29:@20891.4]
  assign Mem1D_16_io_w_en_0 = _T_1035[41]; // @[MemPrimitives.scala 96:27:@20892.4]
  assign Mem1D_17_clock = clock; // @[:@20459.4]
  assign Mem1D_17_reset = reset; // @[:@20460.4]
  assign Mem1D_17_io_r_ofs_0 = _T_2831[8:0]; // @[MemPrimitives.scala 131:28:@22625.4]
  assign Mem1D_17_io_r_backpressure = _T_2831[9]; // @[MemPrimitives.scala 132:32:@22626.4]
  assign Mem1D_17_io_w_ofs_0 = _T_1055[8:0]; // @[MemPrimitives.scala 94:28:@20909.4]
  assign Mem1D_17_io_w_data_0 = _T_1055[40:9]; // @[MemPrimitives.scala 95:29:@20910.4]
  assign Mem1D_17_io_w_en_0 = _T_1055[41]; // @[MemPrimitives.scala 96:27:@20911.4]
  assign Mem1D_18_clock = clock; // @[:@20475.4]
  assign Mem1D_18_reset = reset; // @[:@20476.4]
  assign Mem1D_18_io_r_ofs_0 = _T_2923[8:0]; // @[MemPrimitives.scala 131:28:@22714.4]
  assign Mem1D_18_io_r_backpressure = _T_2923[9]; // @[MemPrimitives.scala 132:32:@22715.4]
  assign Mem1D_18_io_w_ofs_0 = _T_1075[8:0]; // @[MemPrimitives.scala 94:28:@20928.4]
  assign Mem1D_18_io_w_data_0 = _T_1075[40:9]; // @[MemPrimitives.scala 95:29:@20929.4]
  assign Mem1D_18_io_w_en_0 = _T_1075[41]; // @[MemPrimitives.scala 96:27:@20930.4]
  assign Mem1D_19_clock = clock; // @[:@20491.4]
  assign Mem1D_19_reset = reset; // @[:@20492.4]
  assign Mem1D_19_io_r_ofs_0 = _T_3015[8:0]; // @[MemPrimitives.scala 131:28:@22803.4]
  assign Mem1D_19_io_r_backpressure = _T_3015[9]; // @[MemPrimitives.scala 132:32:@22804.4]
  assign Mem1D_19_io_w_ofs_0 = _T_1095[8:0]; // @[MemPrimitives.scala 94:28:@20947.4]
  assign Mem1D_19_io_w_data_0 = _T_1095[40:9]; // @[MemPrimitives.scala 95:29:@20948.4]
  assign Mem1D_19_io_w_en_0 = _T_1095[41]; // @[MemPrimitives.scala 96:27:@20949.4]
  assign Mem1D_20_clock = clock; // @[:@20507.4]
  assign Mem1D_20_reset = reset; // @[:@20508.4]
  assign Mem1D_20_io_r_ofs_0 = _T_3107[8:0]; // @[MemPrimitives.scala 131:28:@22892.4]
  assign Mem1D_20_io_r_backpressure = _T_3107[9]; // @[MemPrimitives.scala 132:32:@22893.4]
  assign Mem1D_20_io_w_ofs_0 = _T_1115[8:0]; // @[MemPrimitives.scala 94:28:@20966.4]
  assign Mem1D_20_io_w_data_0 = _T_1115[40:9]; // @[MemPrimitives.scala 95:29:@20967.4]
  assign Mem1D_20_io_w_en_0 = _T_1115[41]; // @[MemPrimitives.scala 96:27:@20968.4]
  assign Mem1D_21_clock = clock; // @[:@20523.4]
  assign Mem1D_21_reset = reset; // @[:@20524.4]
  assign Mem1D_21_io_r_ofs_0 = _T_3199[8:0]; // @[MemPrimitives.scala 131:28:@22981.4]
  assign Mem1D_21_io_r_backpressure = _T_3199[9]; // @[MemPrimitives.scala 132:32:@22982.4]
  assign Mem1D_21_io_w_ofs_0 = _T_1135[8:0]; // @[MemPrimitives.scala 94:28:@20985.4]
  assign Mem1D_21_io_w_data_0 = _T_1135[40:9]; // @[MemPrimitives.scala 95:29:@20986.4]
  assign Mem1D_21_io_w_en_0 = _T_1135[41]; // @[MemPrimitives.scala 96:27:@20987.4]
  assign Mem1D_22_clock = clock; // @[:@20539.4]
  assign Mem1D_22_reset = reset; // @[:@20540.4]
  assign Mem1D_22_io_r_ofs_0 = _T_3291[8:0]; // @[MemPrimitives.scala 131:28:@23070.4]
  assign Mem1D_22_io_r_backpressure = _T_3291[9]; // @[MemPrimitives.scala 132:32:@23071.4]
  assign Mem1D_22_io_w_ofs_0 = _T_1155[8:0]; // @[MemPrimitives.scala 94:28:@21004.4]
  assign Mem1D_22_io_w_data_0 = _T_1155[40:9]; // @[MemPrimitives.scala 95:29:@21005.4]
  assign Mem1D_22_io_w_en_0 = _T_1155[41]; // @[MemPrimitives.scala 96:27:@21006.4]
  assign Mem1D_23_clock = clock; // @[:@20555.4]
  assign Mem1D_23_reset = reset; // @[:@20556.4]
  assign Mem1D_23_io_r_ofs_0 = _T_3383[8:0]; // @[MemPrimitives.scala 131:28:@23159.4]
  assign Mem1D_23_io_r_backpressure = _T_3383[9]; // @[MemPrimitives.scala 132:32:@23160.4]
  assign Mem1D_23_io_w_ofs_0 = _T_1175[8:0]; // @[MemPrimitives.scala 94:28:@21023.4]
  assign Mem1D_23_io_w_data_0 = _T_1175[40:9]; // @[MemPrimitives.scala 95:29:@21024.4]
  assign Mem1D_23_io_w_en_0 = _T_1175[41]; // @[MemPrimitives.scala 96:27:@21025.4]
  assign StickySelects_clock = clock; // @[:@21063.4]
  assign StickySelects_reset = reset; // @[:@21064.4]
  assign StickySelects_io_ins_0 = io_rPort_1_en_0 & _T_1183; // @[MemPrimitives.scala 125:64:@21065.4]
  assign StickySelects_io_ins_1 = io_rPort_3_en_0 & _T_1189; // @[MemPrimitives.scala 125:64:@21066.4]
  assign StickySelects_io_ins_2 = io_rPort_6_en_0 & _T_1195; // @[MemPrimitives.scala 125:64:@21067.4]
  assign StickySelects_io_ins_3 = io_rPort_8_en_0 & _T_1201; // @[MemPrimitives.scala 125:64:@21068.4]
  assign StickySelects_io_ins_4 = io_rPort_10_en_0 & _T_1207; // @[MemPrimitives.scala 125:64:@21069.4]
  assign StickySelects_io_ins_5 = io_rPort_12_en_0 & _T_1213; // @[MemPrimitives.scala 125:64:@21070.4]
  assign StickySelects_io_ins_6 = io_rPort_15_en_0 & _T_1219; // @[MemPrimitives.scala 125:64:@21071.4]
  assign StickySelects_io_ins_7 = io_rPort_16_en_0 & _T_1225; // @[MemPrimitives.scala 125:64:@21072.4]
  assign StickySelects_io_ins_8 = io_rPort_17_en_0 & _T_1231; // @[MemPrimitives.scala 125:64:@21073.4]
  assign StickySelects_1_clock = clock; // @[:@21152.4]
  assign StickySelects_1_reset = reset; // @[:@21153.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_1275; // @[MemPrimitives.scala 125:64:@21154.4]
  assign StickySelects_1_io_ins_1 = io_rPort_2_en_0 & _T_1281; // @[MemPrimitives.scala 125:64:@21155.4]
  assign StickySelects_1_io_ins_2 = io_rPort_4_en_0 & _T_1287; // @[MemPrimitives.scala 125:64:@21156.4]
  assign StickySelects_1_io_ins_3 = io_rPort_5_en_0 & _T_1293; // @[MemPrimitives.scala 125:64:@21157.4]
  assign StickySelects_1_io_ins_4 = io_rPort_7_en_0 & _T_1299; // @[MemPrimitives.scala 125:64:@21158.4]
  assign StickySelects_1_io_ins_5 = io_rPort_9_en_0 & _T_1305; // @[MemPrimitives.scala 125:64:@21159.4]
  assign StickySelects_1_io_ins_6 = io_rPort_11_en_0 & _T_1311; // @[MemPrimitives.scala 125:64:@21160.4]
  assign StickySelects_1_io_ins_7 = io_rPort_13_en_0 & _T_1317; // @[MemPrimitives.scala 125:64:@21161.4]
  assign StickySelects_1_io_ins_8 = io_rPort_14_en_0 & _T_1323; // @[MemPrimitives.scala 125:64:@21162.4]
  assign StickySelects_2_clock = clock; // @[:@21241.4]
  assign StickySelects_2_reset = reset; // @[:@21242.4]
  assign StickySelects_2_io_ins_0 = io_rPort_1_en_0 & _T_1367; // @[MemPrimitives.scala 125:64:@21243.4]
  assign StickySelects_2_io_ins_1 = io_rPort_3_en_0 & _T_1373; // @[MemPrimitives.scala 125:64:@21244.4]
  assign StickySelects_2_io_ins_2 = io_rPort_6_en_0 & _T_1379; // @[MemPrimitives.scala 125:64:@21245.4]
  assign StickySelects_2_io_ins_3 = io_rPort_8_en_0 & _T_1385; // @[MemPrimitives.scala 125:64:@21246.4]
  assign StickySelects_2_io_ins_4 = io_rPort_10_en_0 & _T_1391; // @[MemPrimitives.scala 125:64:@21247.4]
  assign StickySelects_2_io_ins_5 = io_rPort_12_en_0 & _T_1397; // @[MemPrimitives.scala 125:64:@21248.4]
  assign StickySelects_2_io_ins_6 = io_rPort_15_en_0 & _T_1403; // @[MemPrimitives.scala 125:64:@21249.4]
  assign StickySelects_2_io_ins_7 = io_rPort_16_en_0 & _T_1409; // @[MemPrimitives.scala 125:64:@21250.4]
  assign StickySelects_2_io_ins_8 = io_rPort_17_en_0 & _T_1415; // @[MemPrimitives.scala 125:64:@21251.4]
  assign StickySelects_3_clock = clock; // @[:@21330.4]
  assign StickySelects_3_reset = reset; // @[:@21331.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_1459; // @[MemPrimitives.scala 125:64:@21332.4]
  assign StickySelects_3_io_ins_1 = io_rPort_2_en_0 & _T_1465; // @[MemPrimitives.scala 125:64:@21333.4]
  assign StickySelects_3_io_ins_2 = io_rPort_4_en_0 & _T_1471; // @[MemPrimitives.scala 125:64:@21334.4]
  assign StickySelects_3_io_ins_3 = io_rPort_5_en_0 & _T_1477; // @[MemPrimitives.scala 125:64:@21335.4]
  assign StickySelects_3_io_ins_4 = io_rPort_7_en_0 & _T_1483; // @[MemPrimitives.scala 125:64:@21336.4]
  assign StickySelects_3_io_ins_5 = io_rPort_9_en_0 & _T_1489; // @[MemPrimitives.scala 125:64:@21337.4]
  assign StickySelects_3_io_ins_6 = io_rPort_11_en_0 & _T_1495; // @[MemPrimitives.scala 125:64:@21338.4]
  assign StickySelects_3_io_ins_7 = io_rPort_13_en_0 & _T_1501; // @[MemPrimitives.scala 125:64:@21339.4]
  assign StickySelects_3_io_ins_8 = io_rPort_14_en_0 & _T_1507; // @[MemPrimitives.scala 125:64:@21340.4]
  assign StickySelects_4_clock = clock; // @[:@21419.4]
  assign StickySelects_4_reset = reset; // @[:@21420.4]
  assign StickySelects_4_io_ins_0 = io_rPort_1_en_0 & _T_1551; // @[MemPrimitives.scala 125:64:@21421.4]
  assign StickySelects_4_io_ins_1 = io_rPort_3_en_0 & _T_1557; // @[MemPrimitives.scala 125:64:@21422.4]
  assign StickySelects_4_io_ins_2 = io_rPort_6_en_0 & _T_1563; // @[MemPrimitives.scala 125:64:@21423.4]
  assign StickySelects_4_io_ins_3 = io_rPort_8_en_0 & _T_1569; // @[MemPrimitives.scala 125:64:@21424.4]
  assign StickySelects_4_io_ins_4 = io_rPort_10_en_0 & _T_1575; // @[MemPrimitives.scala 125:64:@21425.4]
  assign StickySelects_4_io_ins_5 = io_rPort_12_en_0 & _T_1581; // @[MemPrimitives.scala 125:64:@21426.4]
  assign StickySelects_4_io_ins_6 = io_rPort_15_en_0 & _T_1587; // @[MemPrimitives.scala 125:64:@21427.4]
  assign StickySelects_4_io_ins_7 = io_rPort_16_en_0 & _T_1593; // @[MemPrimitives.scala 125:64:@21428.4]
  assign StickySelects_4_io_ins_8 = io_rPort_17_en_0 & _T_1599; // @[MemPrimitives.scala 125:64:@21429.4]
  assign StickySelects_5_clock = clock; // @[:@21508.4]
  assign StickySelects_5_reset = reset; // @[:@21509.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_1643; // @[MemPrimitives.scala 125:64:@21510.4]
  assign StickySelects_5_io_ins_1 = io_rPort_2_en_0 & _T_1649; // @[MemPrimitives.scala 125:64:@21511.4]
  assign StickySelects_5_io_ins_2 = io_rPort_4_en_0 & _T_1655; // @[MemPrimitives.scala 125:64:@21512.4]
  assign StickySelects_5_io_ins_3 = io_rPort_5_en_0 & _T_1661; // @[MemPrimitives.scala 125:64:@21513.4]
  assign StickySelects_5_io_ins_4 = io_rPort_7_en_0 & _T_1667; // @[MemPrimitives.scala 125:64:@21514.4]
  assign StickySelects_5_io_ins_5 = io_rPort_9_en_0 & _T_1673; // @[MemPrimitives.scala 125:64:@21515.4]
  assign StickySelects_5_io_ins_6 = io_rPort_11_en_0 & _T_1679; // @[MemPrimitives.scala 125:64:@21516.4]
  assign StickySelects_5_io_ins_7 = io_rPort_13_en_0 & _T_1685; // @[MemPrimitives.scala 125:64:@21517.4]
  assign StickySelects_5_io_ins_8 = io_rPort_14_en_0 & _T_1691; // @[MemPrimitives.scala 125:64:@21518.4]
  assign StickySelects_6_clock = clock; // @[:@21597.4]
  assign StickySelects_6_reset = reset; // @[:@21598.4]
  assign StickySelects_6_io_ins_0 = io_rPort_1_en_0 & _T_1735; // @[MemPrimitives.scala 125:64:@21599.4]
  assign StickySelects_6_io_ins_1 = io_rPort_3_en_0 & _T_1741; // @[MemPrimitives.scala 125:64:@21600.4]
  assign StickySelects_6_io_ins_2 = io_rPort_6_en_0 & _T_1747; // @[MemPrimitives.scala 125:64:@21601.4]
  assign StickySelects_6_io_ins_3 = io_rPort_8_en_0 & _T_1753; // @[MemPrimitives.scala 125:64:@21602.4]
  assign StickySelects_6_io_ins_4 = io_rPort_10_en_0 & _T_1759; // @[MemPrimitives.scala 125:64:@21603.4]
  assign StickySelects_6_io_ins_5 = io_rPort_12_en_0 & _T_1765; // @[MemPrimitives.scala 125:64:@21604.4]
  assign StickySelects_6_io_ins_6 = io_rPort_15_en_0 & _T_1771; // @[MemPrimitives.scala 125:64:@21605.4]
  assign StickySelects_6_io_ins_7 = io_rPort_16_en_0 & _T_1777; // @[MemPrimitives.scala 125:64:@21606.4]
  assign StickySelects_6_io_ins_8 = io_rPort_17_en_0 & _T_1783; // @[MemPrimitives.scala 125:64:@21607.4]
  assign StickySelects_7_clock = clock; // @[:@21686.4]
  assign StickySelects_7_reset = reset; // @[:@21687.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1827; // @[MemPrimitives.scala 125:64:@21688.4]
  assign StickySelects_7_io_ins_1 = io_rPort_2_en_0 & _T_1833; // @[MemPrimitives.scala 125:64:@21689.4]
  assign StickySelects_7_io_ins_2 = io_rPort_4_en_0 & _T_1839; // @[MemPrimitives.scala 125:64:@21690.4]
  assign StickySelects_7_io_ins_3 = io_rPort_5_en_0 & _T_1845; // @[MemPrimitives.scala 125:64:@21691.4]
  assign StickySelects_7_io_ins_4 = io_rPort_7_en_0 & _T_1851; // @[MemPrimitives.scala 125:64:@21692.4]
  assign StickySelects_7_io_ins_5 = io_rPort_9_en_0 & _T_1857; // @[MemPrimitives.scala 125:64:@21693.4]
  assign StickySelects_7_io_ins_6 = io_rPort_11_en_0 & _T_1863; // @[MemPrimitives.scala 125:64:@21694.4]
  assign StickySelects_7_io_ins_7 = io_rPort_13_en_0 & _T_1869; // @[MemPrimitives.scala 125:64:@21695.4]
  assign StickySelects_7_io_ins_8 = io_rPort_14_en_0 & _T_1875; // @[MemPrimitives.scala 125:64:@21696.4]
  assign StickySelects_8_clock = clock; // @[:@21775.4]
  assign StickySelects_8_reset = reset; // @[:@21776.4]
  assign StickySelects_8_io_ins_0 = io_rPort_1_en_0 & _T_1919; // @[MemPrimitives.scala 125:64:@21777.4]
  assign StickySelects_8_io_ins_1 = io_rPort_3_en_0 & _T_1925; // @[MemPrimitives.scala 125:64:@21778.4]
  assign StickySelects_8_io_ins_2 = io_rPort_6_en_0 & _T_1931; // @[MemPrimitives.scala 125:64:@21779.4]
  assign StickySelects_8_io_ins_3 = io_rPort_8_en_0 & _T_1937; // @[MemPrimitives.scala 125:64:@21780.4]
  assign StickySelects_8_io_ins_4 = io_rPort_10_en_0 & _T_1943; // @[MemPrimitives.scala 125:64:@21781.4]
  assign StickySelects_8_io_ins_5 = io_rPort_12_en_0 & _T_1949; // @[MemPrimitives.scala 125:64:@21782.4]
  assign StickySelects_8_io_ins_6 = io_rPort_15_en_0 & _T_1955; // @[MemPrimitives.scala 125:64:@21783.4]
  assign StickySelects_8_io_ins_7 = io_rPort_16_en_0 & _T_1961; // @[MemPrimitives.scala 125:64:@21784.4]
  assign StickySelects_8_io_ins_8 = io_rPort_17_en_0 & _T_1967; // @[MemPrimitives.scala 125:64:@21785.4]
  assign StickySelects_9_clock = clock; // @[:@21864.4]
  assign StickySelects_9_reset = reset; // @[:@21865.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_2011; // @[MemPrimitives.scala 125:64:@21866.4]
  assign StickySelects_9_io_ins_1 = io_rPort_2_en_0 & _T_2017; // @[MemPrimitives.scala 125:64:@21867.4]
  assign StickySelects_9_io_ins_2 = io_rPort_4_en_0 & _T_2023; // @[MemPrimitives.scala 125:64:@21868.4]
  assign StickySelects_9_io_ins_3 = io_rPort_5_en_0 & _T_2029; // @[MemPrimitives.scala 125:64:@21869.4]
  assign StickySelects_9_io_ins_4 = io_rPort_7_en_0 & _T_2035; // @[MemPrimitives.scala 125:64:@21870.4]
  assign StickySelects_9_io_ins_5 = io_rPort_9_en_0 & _T_2041; // @[MemPrimitives.scala 125:64:@21871.4]
  assign StickySelects_9_io_ins_6 = io_rPort_11_en_0 & _T_2047; // @[MemPrimitives.scala 125:64:@21872.4]
  assign StickySelects_9_io_ins_7 = io_rPort_13_en_0 & _T_2053; // @[MemPrimitives.scala 125:64:@21873.4]
  assign StickySelects_9_io_ins_8 = io_rPort_14_en_0 & _T_2059; // @[MemPrimitives.scala 125:64:@21874.4]
  assign StickySelects_10_clock = clock; // @[:@21953.4]
  assign StickySelects_10_reset = reset; // @[:@21954.4]
  assign StickySelects_10_io_ins_0 = io_rPort_1_en_0 & _T_2103; // @[MemPrimitives.scala 125:64:@21955.4]
  assign StickySelects_10_io_ins_1 = io_rPort_3_en_0 & _T_2109; // @[MemPrimitives.scala 125:64:@21956.4]
  assign StickySelects_10_io_ins_2 = io_rPort_6_en_0 & _T_2115; // @[MemPrimitives.scala 125:64:@21957.4]
  assign StickySelects_10_io_ins_3 = io_rPort_8_en_0 & _T_2121; // @[MemPrimitives.scala 125:64:@21958.4]
  assign StickySelects_10_io_ins_4 = io_rPort_10_en_0 & _T_2127; // @[MemPrimitives.scala 125:64:@21959.4]
  assign StickySelects_10_io_ins_5 = io_rPort_12_en_0 & _T_2133; // @[MemPrimitives.scala 125:64:@21960.4]
  assign StickySelects_10_io_ins_6 = io_rPort_15_en_0 & _T_2139; // @[MemPrimitives.scala 125:64:@21961.4]
  assign StickySelects_10_io_ins_7 = io_rPort_16_en_0 & _T_2145; // @[MemPrimitives.scala 125:64:@21962.4]
  assign StickySelects_10_io_ins_8 = io_rPort_17_en_0 & _T_2151; // @[MemPrimitives.scala 125:64:@21963.4]
  assign StickySelects_11_clock = clock; // @[:@22042.4]
  assign StickySelects_11_reset = reset; // @[:@22043.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_2195; // @[MemPrimitives.scala 125:64:@22044.4]
  assign StickySelects_11_io_ins_1 = io_rPort_2_en_0 & _T_2201; // @[MemPrimitives.scala 125:64:@22045.4]
  assign StickySelects_11_io_ins_2 = io_rPort_4_en_0 & _T_2207; // @[MemPrimitives.scala 125:64:@22046.4]
  assign StickySelects_11_io_ins_3 = io_rPort_5_en_0 & _T_2213; // @[MemPrimitives.scala 125:64:@22047.4]
  assign StickySelects_11_io_ins_4 = io_rPort_7_en_0 & _T_2219; // @[MemPrimitives.scala 125:64:@22048.4]
  assign StickySelects_11_io_ins_5 = io_rPort_9_en_0 & _T_2225; // @[MemPrimitives.scala 125:64:@22049.4]
  assign StickySelects_11_io_ins_6 = io_rPort_11_en_0 & _T_2231; // @[MemPrimitives.scala 125:64:@22050.4]
  assign StickySelects_11_io_ins_7 = io_rPort_13_en_0 & _T_2237; // @[MemPrimitives.scala 125:64:@22051.4]
  assign StickySelects_11_io_ins_8 = io_rPort_14_en_0 & _T_2243; // @[MemPrimitives.scala 125:64:@22052.4]
  assign StickySelects_12_clock = clock; // @[:@22131.4]
  assign StickySelects_12_reset = reset; // @[:@22132.4]
  assign StickySelects_12_io_ins_0 = io_rPort_1_en_0 & _T_2287; // @[MemPrimitives.scala 125:64:@22133.4]
  assign StickySelects_12_io_ins_1 = io_rPort_3_en_0 & _T_2293; // @[MemPrimitives.scala 125:64:@22134.4]
  assign StickySelects_12_io_ins_2 = io_rPort_6_en_0 & _T_2299; // @[MemPrimitives.scala 125:64:@22135.4]
  assign StickySelects_12_io_ins_3 = io_rPort_8_en_0 & _T_2305; // @[MemPrimitives.scala 125:64:@22136.4]
  assign StickySelects_12_io_ins_4 = io_rPort_10_en_0 & _T_2311; // @[MemPrimitives.scala 125:64:@22137.4]
  assign StickySelects_12_io_ins_5 = io_rPort_12_en_0 & _T_2317; // @[MemPrimitives.scala 125:64:@22138.4]
  assign StickySelects_12_io_ins_6 = io_rPort_15_en_0 & _T_2323; // @[MemPrimitives.scala 125:64:@22139.4]
  assign StickySelects_12_io_ins_7 = io_rPort_16_en_0 & _T_2329; // @[MemPrimitives.scala 125:64:@22140.4]
  assign StickySelects_12_io_ins_8 = io_rPort_17_en_0 & _T_2335; // @[MemPrimitives.scala 125:64:@22141.4]
  assign StickySelects_13_clock = clock; // @[:@22220.4]
  assign StickySelects_13_reset = reset; // @[:@22221.4]
  assign StickySelects_13_io_ins_0 = io_rPort_0_en_0 & _T_2379; // @[MemPrimitives.scala 125:64:@22222.4]
  assign StickySelects_13_io_ins_1 = io_rPort_2_en_0 & _T_2385; // @[MemPrimitives.scala 125:64:@22223.4]
  assign StickySelects_13_io_ins_2 = io_rPort_4_en_0 & _T_2391; // @[MemPrimitives.scala 125:64:@22224.4]
  assign StickySelects_13_io_ins_3 = io_rPort_5_en_0 & _T_2397; // @[MemPrimitives.scala 125:64:@22225.4]
  assign StickySelects_13_io_ins_4 = io_rPort_7_en_0 & _T_2403; // @[MemPrimitives.scala 125:64:@22226.4]
  assign StickySelects_13_io_ins_5 = io_rPort_9_en_0 & _T_2409; // @[MemPrimitives.scala 125:64:@22227.4]
  assign StickySelects_13_io_ins_6 = io_rPort_11_en_0 & _T_2415; // @[MemPrimitives.scala 125:64:@22228.4]
  assign StickySelects_13_io_ins_7 = io_rPort_13_en_0 & _T_2421; // @[MemPrimitives.scala 125:64:@22229.4]
  assign StickySelects_13_io_ins_8 = io_rPort_14_en_0 & _T_2427; // @[MemPrimitives.scala 125:64:@22230.4]
  assign StickySelects_14_clock = clock; // @[:@22309.4]
  assign StickySelects_14_reset = reset; // @[:@22310.4]
  assign StickySelects_14_io_ins_0 = io_rPort_1_en_0 & _T_2471; // @[MemPrimitives.scala 125:64:@22311.4]
  assign StickySelects_14_io_ins_1 = io_rPort_3_en_0 & _T_2477; // @[MemPrimitives.scala 125:64:@22312.4]
  assign StickySelects_14_io_ins_2 = io_rPort_6_en_0 & _T_2483; // @[MemPrimitives.scala 125:64:@22313.4]
  assign StickySelects_14_io_ins_3 = io_rPort_8_en_0 & _T_2489; // @[MemPrimitives.scala 125:64:@22314.4]
  assign StickySelects_14_io_ins_4 = io_rPort_10_en_0 & _T_2495; // @[MemPrimitives.scala 125:64:@22315.4]
  assign StickySelects_14_io_ins_5 = io_rPort_12_en_0 & _T_2501; // @[MemPrimitives.scala 125:64:@22316.4]
  assign StickySelects_14_io_ins_6 = io_rPort_15_en_0 & _T_2507; // @[MemPrimitives.scala 125:64:@22317.4]
  assign StickySelects_14_io_ins_7 = io_rPort_16_en_0 & _T_2513; // @[MemPrimitives.scala 125:64:@22318.4]
  assign StickySelects_14_io_ins_8 = io_rPort_17_en_0 & _T_2519; // @[MemPrimitives.scala 125:64:@22319.4]
  assign StickySelects_15_clock = clock; // @[:@22398.4]
  assign StickySelects_15_reset = reset; // @[:@22399.4]
  assign StickySelects_15_io_ins_0 = io_rPort_0_en_0 & _T_2563; // @[MemPrimitives.scala 125:64:@22400.4]
  assign StickySelects_15_io_ins_1 = io_rPort_2_en_0 & _T_2569; // @[MemPrimitives.scala 125:64:@22401.4]
  assign StickySelects_15_io_ins_2 = io_rPort_4_en_0 & _T_2575; // @[MemPrimitives.scala 125:64:@22402.4]
  assign StickySelects_15_io_ins_3 = io_rPort_5_en_0 & _T_2581; // @[MemPrimitives.scala 125:64:@22403.4]
  assign StickySelects_15_io_ins_4 = io_rPort_7_en_0 & _T_2587; // @[MemPrimitives.scala 125:64:@22404.4]
  assign StickySelects_15_io_ins_5 = io_rPort_9_en_0 & _T_2593; // @[MemPrimitives.scala 125:64:@22405.4]
  assign StickySelects_15_io_ins_6 = io_rPort_11_en_0 & _T_2599; // @[MemPrimitives.scala 125:64:@22406.4]
  assign StickySelects_15_io_ins_7 = io_rPort_13_en_0 & _T_2605; // @[MemPrimitives.scala 125:64:@22407.4]
  assign StickySelects_15_io_ins_8 = io_rPort_14_en_0 & _T_2611; // @[MemPrimitives.scala 125:64:@22408.4]
  assign StickySelects_16_clock = clock; // @[:@22487.4]
  assign StickySelects_16_reset = reset; // @[:@22488.4]
  assign StickySelects_16_io_ins_0 = io_rPort_1_en_0 & _T_2655; // @[MemPrimitives.scala 125:64:@22489.4]
  assign StickySelects_16_io_ins_1 = io_rPort_3_en_0 & _T_2661; // @[MemPrimitives.scala 125:64:@22490.4]
  assign StickySelects_16_io_ins_2 = io_rPort_6_en_0 & _T_2667; // @[MemPrimitives.scala 125:64:@22491.4]
  assign StickySelects_16_io_ins_3 = io_rPort_8_en_0 & _T_2673; // @[MemPrimitives.scala 125:64:@22492.4]
  assign StickySelects_16_io_ins_4 = io_rPort_10_en_0 & _T_2679; // @[MemPrimitives.scala 125:64:@22493.4]
  assign StickySelects_16_io_ins_5 = io_rPort_12_en_0 & _T_2685; // @[MemPrimitives.scala 125:64:@22494.4]
  assign StickySelects_16_io_ins_6 = io_rPort_15_en_0 & _T_2691; // @[MemPrimitives.scala 125:64:@22495.4]
  assign StickySelects_16_io_ins_7 = io_rPort_16_en_0 & _T_2697; // @[MemPrimitives.scala 125:64:@22496.4]
  assign StickySelects_16_io_ins_8 = io_rPort_17_en_0 & _T_2703; // @[MemPrimitives.scala 125:64:@22497.4]
  assign StickySelects_17_clock = clock; // @[:@22576.4]
  assign StickySelects_17_reset = reset; // @[:@22577.4]
  assign StickySelects_17_io_ins_0 = io_rPort_0_en_0 & _T_2747; // @[MemPrimitives.scala 125:64:@22578.4]
  assign StickySelects_17_io_ins_1 = io_rPort_2_en_0 & _T_2753; // @[MemPrimitives.scala 125:64:@22579.4]
  assign StickySelects_17_io_ins_2 = io_rPort_4_en_0 & _T_2759; // @[MemPrimitives.scala 125:64:@22580.4]
  assign StickySelects_17_io_ins_3 = io_rPort_5_en_0 & _T_2765; // @[MemPrimitives.scala 125:64:@22581.4]
  assign StickySelects_17_io_ins_4 = io_rPort_7_en_0 & _T_2771; // @[MemPrimitives.scala 125:64:@22582.4]
  assign StickySelects_17_io_ins_5 = io_rPort_9_en_0 & _T_2777; // @[MemPrimitives.scala 125:64:@22583.4]
  assign StickySelects_17_io_ins_6 = io_rPort_11_en_0 & _T_2783; // @[MemPrimitives.scala 125:64:@22584.4]
  assign StickySelects_17_io_ins_7 = io_rPort_13_en_0 & _T_2789; // @[MemPrimitives.scala 125:64:@22585.4]
  assign StickySelects_17_io_ins_8 = io_rPort_14_en_0 & _T_2795; // @[MemPrimitives.scala 125:64:@22586.4]
  assign StickySelects_18_clock = clock; // @[:@22665.4]
  assign StickySelects_18_reset = reset; // @[:@22666.4]
  assign StickySelects_18_io_ins_0 = io_rPort_1_en_0 & _T_2839; // @[MemPrimitives.scala 125:64:@22667.4]
  assign StickySelects_18_io_ins_1 = io_rPort_3_en_0 & _T_2845; // @[MemPrimitives.scala 125:64:@22668.4]
  assign StickySelects_18_io_ins_2 = io_rPort_6_en_0 & _T_2851; // @[MemPrimitives.scala 125:64:@22669.4]
  assign StickySelects_18_io_ins_3 = io_rPort_8_en_0 & _T_2857; // @[MemPrimitives.scala 125:64:@22670.4]
  assign StickySelects_18_io_ins_4 = io_rPort_10_en_0 & _T_2863; // @[MemPrimitives.scala 125:64:@22671.4]
  assign StickySelects_18_io_ins_5 = io_rPort_12_en_0 & _T_2869; // @[MemPrimitives.scala 125:64:@22672.4]
  assign StickySelects_18_io_ins_6 = io_rPort_15_en_0 & _T_2875; // @[MemPrimitives.scala 125:64:@22673.4]
  assign StickySelects_18_io_ins_7 = io_rPort_16_en_0 & _T_2881; // @[MemPrimitives.scala 125:64:@22674.4]
  assign StickySelects_18_io_ins_8 = io_rPort_17_en_0 & _T_2887; // @[MemPrimitives.scala 125:64:@22675.4]
  assign StickySelects_19_clock = clock; // @[:@22754.4]
  assign StickySelects_19_reset = reset; // @[:@22755.4]
  assign StickySelects_19_io_ins_0 = io_rPort_0_en_0 & _T_2931; // @[MemPrimitives.scala 125:64:@22756.4]
  assign StickySelects_19_io_ins_1 = io_rPort_2_en_0 & _T_2937; // @[MemPrimitives.scala 125:64:@22757.4]
  assign StickySelects_19_io_ins_2 = io_rPort_4_en_0 & _T_2943; // @[MemPrimitives.scala 125:64:@22758.4]
  assign StickySelects_19_io_ins_3 = io_rPort_5_en_0 & _T_2949; // @[MemPrimitives.scala 125:64:@22759.4]
  assign StickySelects_19_io_ins_4 = io_rPort_7_en_0 & _T_2955; // @[MemPrimitives.scala 125:64:@22760.4]
  assign StickySelects_19_io_ins_5 = io_rPort_9_en_0 & _T_2961; // @[MemPrimitives.scala 125:64:@22761.4]
  assign StickySelects_19_io_ins_6 = io_rPort_11_en_0 & _T_2967; // @[MemPrimitives.scala 125:64:@22762.4]
  assign StickySelects_19_io_ins_7 = io_rPort_13_en_0 & _T_2973; // @[MemPrimitives.scala 125:64:@22763.4]
  assign StickySelects_19_io_ins_8 = io_rPort_14_en_0 & _T_2979; // @[MemPrimitives.scala 125:64:@22764.4]
  assign StickySelects_20_clock = clock; // @[:@22843.4]
  assign StickySelects_20_reset = reset; // @[:@22844.4]
  assign StickySelects_20_io_ins_0 = io_rPort_1_en_0 & _T_3023; // @[MemPrimitives.scala 125:64:@22845.4]
  assign StickySelects_20_io_ins_1 = io_rPort_3_en_0 & _T_3029; // @[MemPrimitives.scala 125:64:@22846.4]
  assign StickySelects_20_io_ins_2 = io_rPort_6_en_0 & _T_3035; // @[MemPrimitives.scala 125:64:@22847.4]
  assign StickySelects_20_io_ins_3 = io_rPort_8_en_0 & _T_3041; // @[MemPrimitives.scala 125:64:@22848.4]
  assign StickySelects_20_io_ins_4 = io_rPort_10_en_0 & _T_3047; // @[MemPrimitives.scala 125:64:@22849.4]
  assign StickySelects_20_io_ins_5 = io_rPort_12_en_0 & _T_3053; // @[MemPrimitives.scala 125:64:@22850.4]
  assign StickySelects_20_io_ins_6 = io_rPort_15_en_0 & _T_3059; // @[MemPrimitives.scala 125:64:@22851.4]
  assign StickySelects_20_io_ins_7 = io_rPort_16_en_0 & _T_3065; // @[MemPrimitives.scala 125:64:@22852.4]
  assign StickySelects_20_io_ins_8 = io_rPort_17_en_0 & _T_3071; // @[MemPrimitives.scala 125:64:@22853.4]
  assign StickySelects_21_clock = clock; // @[:@22932.4]
  assign StickySelects_21_reset = reset; // @[:@22933.4]
  assign StickySelects_21_io_ins_0 = io_rPort_0_en_0 & _T_3115; // @[MemPrimitives.scala 125:64:@22934.4]
  assign StickySelects_21_io_ins_1 = io_rPort_2_en_0 & _T_3121; // @[MemPrimitives.scala 125:64:@22935.4]
  assign StickySelects_21_io_ins_2 = io_rPort_4_en_0 & _T_3127; // @[MemPrimitives.scala 125:64:@22936.4]
  assign StickySelects_21_io_ins_3 = io_rPort_5_en_0 & _T_3133; // @[MemPrimitives.scala 125:64:@22937.4]
  assign StickySelects_21_io_ins_4 = io_rPort_7_en_0 & _T_3139; // @[MemPrimitives.scala 125:64:@22938.4]
  assign StickySelects_21_io_ins_5 = io_rPort_9_en_0 & _T_3145; // @[MemPrimitives.scala 125:64:@22939.4]
  assign StickySelects_21_io_ins_6 = io_rPort_11_en_0 & _T_3151; // @[MemPrimitives.scala 125:64:@22940.4]
  assign StickySelects_21_io_ins_7 = io_rPort_13_en_0 & _T_3157; // @[MemPrimitives.scala 125:64:@22941.4]
  assign StickySelects_21_io_ins_8 = io_rPort_14_en_0 & _T_3163; // @[MemPrimitives.scala 125:64:@22942.4]
  assign StickySelects_22_clock = clock; // @[:@23021.4]
  assign StickySelects_22_reset = reset; // @[:@23022.4]
  assign StickySelects_22_io_ins_0 = io_rPort_1_en_0 & _T_3207; // @[MemPrimitives.scala 125:64:@23023.4]
  assign StickySelects_22_io_ins_1 = io_rPort_3_en_0 & _T_3213; // @[MemPrimitives.scala 125:64:@23024.4]
  assign StickySelects_22_io_ins_2 = io_rPort_6_en_0 & _T_3219; // @[MemPrimitives.scala 125:64:@23025.4]
  assign StickySelects_22_io_ins_3 = io_rPort_8_en_0 & _T_3225; // @[MemPrimitives.scala 125:64:@23026.4]
  assign StickySelects_22_io_ins_4 = io_rPort_10_en_0 & _T_3231; // @[MemPrimitives.scala 125:64:@23027.4]
  assign StickySelects_22_io_ins_5 = io_rPort_12_en_0 & _T_3237; // @[MemPrimitives.scala 125:64:@23028.4]
  assign StickySelects_22_io_ins_6 = io_rPort_15_en_0 & _T_3243; // @[MemPrimitives.scala 125:64:@23029.4]
  assign StickySelects_22_io_ins_7 = io_rPort_16_en_0 & _T_3249; // @[MemPrimitives.scala 125:64:@23030.4]
  assign StickySelects_22_io_ins_8 = io_rPort_17_en_0 & _T_3255; // @[MemPrimitives.scala 125:64:@23031.4]
  assign StickySelects_23_clock = clock; // @[:@23110.4]
  assign StickySelects_23_reset = reset; // @[:@23111.4]
  assign StickySelects_23_io_ins_0 = io_rPort_0_en_0 & _T_3299; // @[MemPrimitives.scala 125:64:@23112.4]
  assign StickySelects_23_io_ins_1 = io_rPort_2_en_0 & _T_3305; // @[MemPrimitives.scala 125:64:@23113.4]
  assign StickySelects_23_io_ins_2 = io_rPort_4_en_0 & _T_3311; // @[MemPrimitives.scala 125:64:@23114.4]
  assign StickySelects_23_io_ins_3 = io_rPort_5_en_0 & _T_3317; // @[MemPrimitives.scala 125:64:@23115.4]
  assign StickySelects_23_io_ins_4 = io_rPort_7_en_0 & _T_3323; // @[MemPrimitives.scala 125:64:@23116.4]
  assign StickySelects_23_io_ins_5 = io_rPort_9_en_0 & _T_3329; // @[MemPrimitives.scala 125:64:@23117.4]
  assign StickySelects_23_io_ins_6 = io_rPort_11_en_0 & _T_3335; // @[MemPrimitives.scala 125:64:@23118.4]
  assign StickySelects_23_io_ins_7 = io_rPort_13_en_0 & _T_3341; // @[MemPrimitives.scala 125:64:@23119.4]
  assign StickySelects_23_io_ins_8 = io_rPort_14_en_0 & _T_3347; // @[MemPrimitives.scala 125:64:@23120.4]
  assign RetimeWrapper_clock = clock; // @[:@23200.4]
  assign RetimeWrapper_reset = reset; // @[:@23201.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23203.4]
  assign RetimeWrapper_io_in = _T_1275 & io_rPort_0_en_0; // @[package.scala 94:16:@23202.4]
  assign RetimeWrapper_1_clock = clock; // @[:@23208.4]
  assign RetimeWrapper_1_reset = reset; // @[:@23209.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23211.4]
  assign RetimeWrapper_1_io_in = _T_1459 & io_rPort_0_en_0; // @[package.scala 94:16:@23210.4]
  assign RetimeWrapper_2_clock = clock; // @[:@23216.4]
  assign RetimeWrapper_2_reset = reset; // @[:@23217.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23219.4]
  assign RetimeWrapper_2_io_in = _T_1643 & io_rPort_0_en_0; // @[package.scala 94:16:@23218.4]
  assign RetimeWrapper_3_clock = clock; // @[:@23224.4]
  assign RetimeWrapper_3_reset = reset; // @[:@23225.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23227.4]
  assign RetimeWrapper_3_io_in = _T_1827 & io_rPort_0_en_0; // @[package.scala 94:16:@23226.4]
  assign RetimeWrapper_4_clock = clock; // @[:@23232.4]
  assign RetimeWrapper_4_reset = reset; // @[:@23233.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23235.4]
  assign RetimeWrapper_4_io_in = _T_2011 & io_rPort_0_en_0; // @[package.scala 94:16:@23234.4]
  assign RetimeWrapper_5_clock = clock; // @[:@23240.4]
  assign RetimeWrapper_5_reset = reset; // @[:@23241.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23243.4]
  assign RetimeWrapper_5_io_in = _T_2195 & io_rPort_0_en_0; // @[package.scala 94:16:@23242.4]
  assign RetimeWrapper_6_clock = clock; // @[:@23248.4]
  assign RetimeWrapper_6_reset = reset; // @[:@23249.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23251.4]
  assign RetimeWrapper_6_io_in = _T_2379 & io_rPort_0_en_0; // @[package.scala 94:16:@23250.4]
  assign RetimeWrapper_7_clock = clock; // @[:@23256.4]
  assign RetimeWrapper_7_reset = reset; // @[:@23257.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23259.4]
  assign RetimeWrapper_7_io_in = _T_2563 & io_rPort_0_en_0; // @[package.scala 94:16:@23258.4]
  assign RetimeWrapper_8_clock = clock; // @[:@23264.4]
  assign RetimeWrapper_8_reset = reset; // @[:@23265.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23267.4]
  assign RetimeWrapper_8_io_in = _T_2747 & io_rPort_0_en_0; // @[package.scala 94:16:@23266.4]
  assign RetimeWrapper_9_clock = clock; // @[:@23272.4]
  assign RetimeWrapper_9_reset = reset; // @[:@23273.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23275.4]
  assign RetimeWrapper_9_io_in = _T_2931 & io_rPort_0_en_0; // @[package.scala 94:16:@23274.4]
  assign RetimeWrapper_10_clock = clock; // @[:@23280.4]
  assign RetimeWrapper_10_reset = reset; // @[:@23281.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23283.4]
  assign RetimeWrapper_10_io_in = _T_3115 & io_rPort_0_en_0; // @[package.scala 94:16:@23282.4]
  assign RetimeWrapper_11_clock = clock; // @[:@23288.4]
  assign RetimeWrapper_11_reset = reset; // @[:@23289.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@23291.4]
  assign RetimeWrapper_11_io_in = _T_3299 & io_rPort_0_en_0; // @[package.scala 94:16:@23290.4]
  assign RetimeWrapper_12_clock = clock; // @[:@23344.4]
  assign RetimeWrapper_12_reset = reset; // @[:@23345.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23347.4]
  assign RetimeWrapper_12_io_in = _T_1183 & io_rPort_1_en_0; // @[package.scala 94:16:@23346.4]
  assign RetimeWrapper_13_clock = clock; // @[:@23352.4]
  assign RetimeWrapper_13_reset = reset; // @[:@23353.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23355.4]
  assign RetimeWrapper_13_io_in = _T_1367 & io_rPort_1_en_0; // @[package.scala 94:16:@23354.4]
  assign RetimeWrapper_14_clock = clock; // @[:@23360.4]
  assign RetimeWrapper_14_reset = reset; // @[:@23361.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23363.4]
  assign RetimeWrapper_14_io_in = _T_1551 & io_rPort_1_en_0; // @[package.scala 94:16:@23362.4]
  assign RetimeWrapper_15_clock = clock; // @[:@23368.4]
  assign RetimeWrapper_15_reset = reset; // @[:@23369.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23371.4]
  assign RetimeWrapper_15_io_in = _T_1735 & io_rPort_1_en_0; // @[package.scala 94:16:@23370.4]
  assign RetimeWrapper_16_clock = clock; // @[:@23376.4]
  assign RetimeWrapper_16_reset = reset; // @[:@23377.4]
  assign RetimeWrapper_16_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23379.4]
  assign RetimeWrapper_16_io_in = _T_1919 & io_rPort_1_en_0; // @[package.scala 94:16:@23378.4]
  assign RetimeWrapper_17_clock = clock; // @[:@23384.4]
  assign RetimeWrapper_17_reset = reset; // @[:@23385.4]
  assign RetimeWrapper_17_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23387.4]
  assign RetimeWrapper_17_io_in = _T_2103 & io_rPort_1_en_0; // @[package.scala 94:16:@23386.4]
  assign RetimeWrapper_18_clock = clock; // @[:@23392.4]
  assign RetimeWrapper_18_reset = reset; // @[:@23393.4]
  assign RetimeWrapper_18_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23395.4]
  assign RetimeWrapper_18_io_in = _T_2287 & io_rPort_1_en_0; // @[package.scala 94:16:@23394.4]
  assign RetimeWrapper_19_clock = clock; // @[:@23400.4]
  assign RetimeWrapper_19_reset = reset; // @[:@23401.4]
  assign RetimeWrapper_19_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23403.4]
  assign RetimeWrapper_19_io_in = _T_2471 & io_rPort_1_en_0; // @[package.scala 94:16:@23402.4]
  assign RetimeWrapper_20_clock = clock; // @[:@23408.4]
  assign RetimeWrapper_20_reset = reset; // @[:@23409.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23411.4]
  assign RetimeWrapper_20_io_in = _T_2655 & io_rPort_1_en_0; // @[package.scala 94:16:@23410.4]
  assign RetimeWrapper_21_clock = clock; // @[:@23416.4]
  assign RetimeWrapper_21_reset = reset; // @[:@23417.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23419.4]
  assign RetimeWrapper_21_io_in = _T_2839 & io_rPort_1_en_0; // @[package.scala 94:16:@23418.4]
  assign RetimeWrapper_22_clock = clock; // @[:@23424.4]
  assign RetimeWrapper_22_reset = reset; // @[:@23425.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23427.4]
  assign RetimeWrapper_22_io_in = _T_3023 & io_rPort_1_en_0; // @[package.scala 94:16:@23426.4]
  assign RetimeWrapper_23_clock = clock; // @[:@23432.4]
  assign RetimeWrapper_23_reset = reset; // @[:@23433.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@23435.4]
  assign RetimeWrapper_23_io_in = _T_3207 & io_rPort_1_en_0; // @[package.scala 94:16:@23434.4]
  assign RetimeWrapper_24_clock = clock; // @[:@23488.4]
  assign RetimeWrapper_24_reset = reset; // @[:@23489.4]
  assign RetimeWrapper_24_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23491.4]
  assign RetimeWrapper_24_io_in = _T_1281 & io_rPort_2_en_0; // @[package.scala 94:16:@23490.4]
  assign RetimeWrapper_25_clock = clock; // @[:@23496.4]
  assign RetimeWrapper_25_reset = reset; // @[:@23497.4]
  assign RetimeWrapper_25_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23499.4]
  assign RetimeWrapper_25_io_in = _T_1465 & io_rPort_2_en_0; // @[package.scala 94:16:@23498.4]
  assign RetimeWrapper_26_clock = clock; // @[:@23504.4]
  assign RetimeWrapper_26_reset = reset; // @[:@23505.4]
  assign RetimeWrapper_26_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23507.4]
  assign RetimeWrapper_26_io_in = _T_1649 & io_rPort_2_en_0; // @[package.scala 94:16:@23506.4]
  assign RetimeWrapper_27_clock = clock; // @[:@23512.4]
  assign RetimeWrapper_27_reset = reset; // @[:@23513.4]
  assign RetimeWrapper_27_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23515.4]
  assign RetimeWrapper_27_io_in = _T_1833 & io_rPort_2_en_0; // @[package.scala 94:16:@23514.4]
  assign RetimeWrapper_28_clock = clock; // @[:@23520.4]
  assign RetimeWrapper_28_reset = reset; // @[:@23521.4]
  assign RetimeWrapper_28_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23523.4]
  assign RetimeWrapper_28_io_in = _T_2017 & io_rPort_2_en_0; // @[package.scala 94:16:@23522.4]
  assign RetimeWrapper_29_clock = clock; // @[:@23528.4]
  assign RetimeWrapper_29_reset = reset; // @[:@23529.4]
  assign RetimeWrapper_29_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23531.4]
  assign RetimeWrapper_29_io_in = _T_2201 & io_rPort_2_en_0; // @[package.scala 94:16:@23530.4]
  assign RetimeWrapper_30_clock = clock; // @[:@23536.4]
  assign RetimeWrapper_30_reset = reset; // @[:@23537.4]
  assign RetimeWrapper_30_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23539.4]
  assign RetimeWrapper_30_io_in = _T_2385 & io_rPort_2_en_0; // @[package.scala 94:16:@23538.4]
  assign RetimeWrapper_31_clock = clock; // @[:@23544.4]
  assign RetimeWrapper_31_reset = reset; // @[:@23545.4]
  assign RetimeWrapper_31_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23547.4]
  assign RetimeWrapper_31_io_in = _T_2569 & io_rPort_2_en_0; // @[package.scala 94:16:@23546.4]
  assign RetimeWrapper_32_clock = clock; // @[:@23552.4]
  assign RetimeWrapper_32_reset = reset; // @[:@23553.4]
  assign RetimeWrapper_32_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23555.4]
  assign RetimeWrapper_32_io_in = _T_2753 & io_rPort_2_en_0; // @[package.scala 94:16:@23554.4]
  assign RetimeWrapper_33_clock = clock; // @[:@23560.4]
  assign RetimeWrapper_33_reset = reset; // @[:@23561.4]
  assign RetimeWrapper_33_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23563.4]
  assign RetimeWrapper_33_io_in = _T_2937 & io_rPort_2_en_0; // @[package.scala 94:16:@23562.4]
  assign RetimeWrapper_34_clock = clock; // @[:@23568.4]
  assign RetimeWrapper_34_reset = reset; // @[:@23569.4]
  assign RetimeWrapper_34_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23571.4]
  assign RetimeWrapper_34_io_in = _T_3121 & io_rPort_2_en_0; // @[package.scala 94:16:@23570.4]
  assign RetimeWrapper_35_clock = clock; // @[:@23576.4]
  assign RetimeWrapper_35_reset = reset; // @[:@23577.4]
  assign RetimeWrapper_35_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@23579.4]
  assign RetimeWrapper_35_io_in = _T_3305 & io_rPort_2_en_0; // @[package.scala 94:16:@23578.4]
  assign RetimeWrapper_36_clock = clock; // @[:@23632.4]
  assign RetimeWrapper_36_reset = reset; // @[:@23633.4]
  assign RetimeWrapper_36_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23635.4]
  assign RetimeWrapper_36_io_in = _T_1189 & io_rPort_3_en_0; // @[package.scala 94:16:@23634.4]
  assign RetimeWrapper_37_clock = clock; // @[:@23640.4]
  assign RetimeWrapper_37_reset = reset; // @[:@23641.4]
  assign RetimeWrapper_37_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23643.4]
  assign RetimeWrapper_37_io_in = _T_1373 & io_rPort_3_en_0; // @[package.scala 94:16:@23642.4]
  assign RetimeWrapper_38_clock = clock; // @[:@23648.4]
  assign RetimeWrapper_38_reset = reset; // @[:@23649.4]
  assign RetimeWrapper_38_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23651.4]
  assign RetimeWrapper_38_io_in = _T_1557 & io_rPort_3_en_0; // @[package.scala 94:16:@23650.4]
  assign RetimeWrapper_39_clock = clock; // @[:@23656.4]
  assign RetimeWrapper_39_reset = reset; // @[:@23657.4]
  assign RetimeWrapper_39_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23659.4]
  assign RetimeWrapper_39_io_in = _T_1741 & io_rPort_3_en_0; // @[package.scala 94:16:@23658.4]
  assign RetimeWrapper_40_clock = clock; // @[:@23664.4]
  assign RetimeWrapper_40_reset = reset; // @[:@23665.4]
  assign RetimeWrapper_40_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23667.4]
  assign RetimeWrapper_40_io_in = _T_1925 & io_rPort_3_en_0; // @[package.scala 94:16:@23666.4]
  assign RetimeWrapper_41_clock = clock; // @[:@23672.4]
  assign RetimeWrapper_41_reset = reset; // @[:@23673.4]
  assign RetimeWrapper_41_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23675.4]
  assign RetimeWrapper_41_io_in = _T_2109 & io_rPort_3_en_0; // @[package.scala 94:16:@23674.4]
  assign RetimeWrapper_42_clock = clock; // @[:@23680.4]
  assign RetimeWrapper_42_reset = reset; // @[:@23681.4]
  assign RetimeWrapper_42_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23683.4]
  assign RetimeWrapper_42_io_in = _T_2293 & io_rPort_3_en_0; // @[package.scala 94:16:@23682.4]
  assign RetimeWrapper_43_clock = clock; // @[:@23688.4]
  assign RetimeWrapper_43_reset = reset; // @[:@23689.4]
  assign RetimeWrapper_43_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23691.4]
  assign RetimeWrapper_43_io_in = _T_2477 & io_rPort_3_en_0; // @[package.scala 94:16:@23690.4]
  assign RetimeWrapper_44_clock = clock; // @[:@23696.4]
  assign RetimeWrapper_44_reset = reset; // @[:@23697.4]
  assign RetimeWrapper_44_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23699.4]
  assign RetimeWrapper_44_io_in = _T_2661 & io_rPort_3_en_0; // @[package.scala 94:16:@23698.4]
  assign RetimeWrapper_45_clock = clock; // @[:@23704.4]
  assign RetimeWrapper_45_reset = reset; // @[:@23705.4]
  assign RetimeWrapper_45_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23707.4]
  assign RetimeWrapper_45_io_in = _T_2845 & io_rPort_3_en_0; // @[package.scala 94:16:@23706.4]
  assign RetimeWrapper_46_clock = clock; // @[:@23712.4]
  assign RetimeWrapper_46_reset = reset; // @[:@23713.4]
  assign RetimeWrapper_46_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23715.4]
  assign RetimeWrapper_46_io_in = _T_3029 & io_rPort_3_en_0; // @[package.scala 94:16:@23714.4]
  assign RetimeWrapper_47_clock = clock; // @[:@23720.4]
  assign RetimeWrapper_47_reset = reset; // @[:@23721.4]
  assign RetimeWrapper_47_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@23723.4]
  assign RetimeWrapper_47_io_in = _T_3213 & io_rPort_3_en_0; // @[package.scala 94:16:@23722.4]
  assign RetimeWrapper_48_clock = clock; // @[:@23776.4]
  assign RetimeWrapper_48_reset = reset; // @[:@23777.4]
  assign RetimeWrapper_48_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23779.4]
  assign RetimeWrapper_48_io_in = _T_1287 & io_rPort_4_en_0; // @[package.scala 94:16:@23778.4]
  assign RetimeWrapper_49_clock = clock; // @[:@23784.4]
  assign RetimeWrapper_49_reset = reset; // @[:@23785.4]
  assign RetimeWrapper_49_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23787.4]
  assign RetimeWrapper_49_io_in = _T_1471 & io_rPort_4_en_0; // @[package.scala 94:16:@23786.4]
  assign RetimeWrapper_50_clock = clock; // @[:@23792.4]
  assign RetimeWrapper_50_reset = reset; // @[:@23793.4]
  assign RetimeWrapper_50_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23795.4]
  assign RetimeWrapper_50_io_in = _T_1655 & io_rPort_4_en_0; // @[package.scala 94:16:@23794.4]
  assign RetimeWrapper_51_clock = clock; // @[:@23800.4]
  assign RetimeWrapper_51_reset = reset; // @[:@23801.4]
  assign RetimeWrapper_51_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23803.4]
  assign RetimeWrapper_51_io_in = _T_1839 & io_rPort_4_en_0; // @[package.scala 94:16:@23802.4]
  assign RetimeWrapper_52_clock = clock; // @[:@23808.4]
  assign RetimeWrapper_52_reset = reset; // @[:@23809.4]
  assign RetimeWrapper_52_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23811.4]
  assign RetimeWrapper_52_io_in = _T_2023 & io_rPort_4_en_0; // @[package.scala 94:16:@23810.4]
  assign RetimeWrapper_53_clock = clock; // @[:@23816.4]
  assign RetimeWrapper_53_reset = reset; // @[:@23817.4]
  assign RetimeWrapper_53_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23819.4]
  assign RetimeWrapper_53_io_in = _T_2207 & io_rPort_4_en_0; // @[package.scala 94:16:@23818.4]
  assign RetimeWrapper_54_clock = clock; // @[:@23824.4]
  assign RetimeWrapper_54_reset = reset; // @[:@23825.4]
  assign RetimeWrapper_54_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23827.4]
  assign RetimeWrapper_54_io_in = _T_2391 & io_rPort_4_en_0; // @[package.scala 94:16:@23826.4]
  assign RetimeWrapper_55_clock = clock; // @[:@23832.4]
  assign RetimeWrapper_55_reset = reset; // @[:@23833.4]
  assign RetimeWrapper_55_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23835.4]
  assign RetimeWrapper_55_io_in = _T_2575 & io_rPort_4_en_0; // @[package.scala 94:16:@23834.4]
  assign RetimeWrapper_56_clock = clock; // @[:@23840.4]
  assign RetimeWrapper_56_reset = reset; // @[:@23841.4]
  assign RetimeWrapper_56_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23843.4]
  assign RetimeWrapper_56_io_in = _T_2759 & io_rPort_4_en_0; // @[package.scala 94:16:@23842.4]
  assign RetimeWrapper_57_clock = clock; // @[:@23848.4]
  assign RetimeWrapper_57_reset = reset; // @[:@23849.4]
  assign RetimeWrapper_57_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23851.4]
  assign RetimeWrapper_57_io_in = _T_2943 & io_rPort_4_en_0; // @[package.scala 94:16:@23850.4]
  assign RetimeWrapper_58_clock = clock; // @[:@23856.4]
  assign RetimeWrapper_58_reset = reset; // @[:@23857.4]
  assign RetimeWrapper_58_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23859.4]
  assign RetimeWrapper_58_io_in = _T_3127 & io_rPort_4_en_0; // @[package.scala 94:16:@23858.4]
  assign RetimeWrapper_59_clock = clock; // @[:@23864.4]
  assign RetimeWrapper_59_reset = reset; // @[:@23865.4]
  assign RetimeWrapper_59_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23867.4]
  assign RetimeWrapper_59_io_in = _T_3311 & io_rPort_4_en_0; // @[package.scala 94:16:@23866.4]
  assign RetimeWrapper_60_clock = clock; // @[:@23920.4]
  assign RetimeWrapper_60_reset = reset; // @[:@23921.4]
  assign RetimeWrapper_60_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23923.4]
  assign RetimeWrapper_60_io_in = _T_1293 & io_rPort_5_en_0; // @[package.scala 94:16:@23922.4]
  assign RetimeWrapper_61_clock = clock; // @[:@23928.4]
  assign RetimeWrapper_61_reset = reset; // @[:@23929.4]
  assign RetimeWrapper_61_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23931.4]
  assign RetimeWrapper_61_io_in = _T_1477 & io_rPort_5_en_0; // @[package.scala 94:16:@23930.4]
  assign RetimeWrapper_62_clock = clock; // @[:@23936.4]
  assign RetimeWrapper_62_reset = reset; // @[:@23937.4]
  assign RetimeWrapper_62_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23939.4]
  assign RetimeWrapper_62_io_in = _T_1661 & io_rPort_5_en_0; // @[package.scala 94:16:@23938.4]
  assign RetimeWrapper_63_clock = clock; // @[:@23944.4]
  assign RetimeWrapper_63_reset = reset; // @[:@23945.4]
  assign RetimeWrapper_63_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23947.4]
  assign RetimeWrapper_63_io_in = _T_1845 & io_rPort_5_en_0; // @[package.scala 94:16:@23946.4]
  assign RetimeWrapper_64_clock = clock; // @[:@23952.4]
  assign RetimeWrapper_64_reset = reset; // @[:@23953.4]
  assign RetimeWrapper_64_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23955.4]
  assign RetimeWrapper_64_io_in = _T_2029 & io_rPort_5_en_0; // @[package.scala 94:16:@23954.4]
  assign RetimeWrapper_65_clock = clock; // @[:@23960.4]
  assign RetimeWrapper_65_reset = reset; // @[:@23961.4]
  assign RetimeWrapper_65_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23963.4]
  assign RetimeWrapper_65_io_in = _T_2213 & io_rPort_5_en_0; // @[package.scala 94:16:@23962.4]
  assign RetimeWrapper_66_clock = clock; // @[:@23968.4]
  assign RetimeWrapper_66_reset = reset; // @[:@23969.4]
  assign RetimeWrapper_66_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23971.4]
  assign RetimeWrapper_66_io_in = _T_2397 & io_rPort_5_en_0; // @[package.scala 94:16:@23970.4]
  assign RetimeWrapper_67_clock = clock; // @[:@23976.4]
  assign RetimeWrapper_67_reset = reset; // @[:@23977.4]
  assign RetimeWrapper_67_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23979.4]
  assign RetimeWrapper_67_io_in = _T_2581 & io_rPort_5_en_0; // @[package.scala 94:16:@23978.4]
  assign RetimeWrapper_68_clock = clock; // @[:@23984.4]
  assign RetimeWrapper_68_reset = reset; // @[:@23985.4]
  assign RetimeWrapper_68_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23987.4]
  assign RetimeWrapper_68_io_in = _T_2765 & io_rPort_5_en_0; // @[package.scala 94:16:@23986.4]
  assign RetimeWrapper_69_clock = clock; // @[:@23992.4]
  assign RetimeWrapper_69_reset = reset; // @[:@23993.4]
  assign RetimeWrapper_69_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23995.4]
  assign RetimeWrapper_69_io_in = _T_2949 & io_rPort_5_en_0; // @[package.scala 94:16:@23994.4]
  assign RetimeWrapper_70_clock = clock; // @[:@24000.4]
  assign RetimeWrapper_70_reset = reset; // @[:@24001.4]
  assign RetimeWrapper_70_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@24003.4]
  assign RetimeWrapper_70_io_in = _T_3133 & io_rPort_5_en_0; // @[package.scala 94:16:@24002.4]
  assign RetimeWrapper_71_clock = clock; // @[:@24008.4]
  assign RetimeWrapper_71_reset = reset; // @[:@24009.4]
  assign RetimeWrapper_71_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@24011.4]
  assign RetimeWrapper_71_io_in = _T_3317 & io_rPort_5_en_0; // @[package.scala 94:16:@24010.4]
  assign RetimeWrapper_72_clock = clock; // @[:@24064.4]
  assign RetimeWrapper_72_reset = reset; // @[:@24065.4]
  assign RetimeWrapper_72_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24067.4]
  assign RetimeWrapper_72_io_in = _T_1195 & io_rPort_6_en_0; // @[package.scala 94:16:@24066.4]
  assign RetimeWrapper_73_clock = clock; // @[:@24072.4]
  assign RetimeWrapper_73_reset = reset; // @[:@24073.4]
  assign RetimeWrapper_73_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24075.4]
  assign RetimeWrapper_73_io_in = _T_1379 & io_rPort_6_en_0; // @[package.scala 94:16:@24074.4]
  assign RetimeWrapper_74_clock = clock; // @[:@24080.4]
  assign RetimeWrapper_74_reset = reset; // @[:@24081.4]
  assign RetimeWrapper_74_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24083.4]
  assign RetimeWrapper_74_io_in = _T_1563 & io_rPort_6_en_0; // @[package.scala 94:16:@24082.4]
  assign RetimeWrapper_75_clock = clock; // @[:@24088.4]
  assign RetimeWrapper_75_reset = reset; // @[:@24089.4]
  assign RetimeWrapper_75_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24091.4]
  assign RetimeWrapper_75_io_in = _T_1747 & io_rPort_6_en_0; // @[package.scala 94:16:@24090.4]
  assign RetimeWrapper_76_clock = clock; // @[:@24096.4]
  assign RetimeWrapper_76_reset = reset; // @[:@24097.4]
  assign RetimeWrapper_76_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24099.4]
  assign RetimeWrapper_76_io_in = _T_1931 & io_rPort_6_en_0; // @[package.scala 94:16:@24098.4]
  assign RetimeWrapper_77_clock = clock; // @[:@24104.4]
  assign RetimeWrapper_77_reset = reset; // @[:@24105.4]
  assign RetimeWrapper_77_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24107.4]
  assign RetimeWrapper_77_io_in = _T_2115 & io_rPort_6_en_0; // @[package.scala 94:16:@24106.4]
  assign RetimeWrapper_78_clock = clock; // @[:@24112.4]
  assign RetimeWrapper_78_reset = reset; // @[:@24113.4]
  assign RetimeWrapper_78_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24115.4]
  assign RetimeWrapper_78_io_in = _T_2299 & io_rPort_6_en_0; // @[package.scala 94:16:@24114.4]
  assign RetimeWrapper_79_clock = clock; // @[:@24120.4]
  assign RetimeWrapper_79_reset = reset; // @[:@24121.4]
  assign RetimeWrapper_79_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24123.4]
  assign RetimeWrapper_79_io_in = _T_2483 & io_rPort_6_en_0; // @[package.scala 94:16:@24122.4]
  assign RetimeWrapper_80_clock = clock; // @[:@24128.4]
  assign RetimeWrapper_80_reset = reset; // @[:@24129.4]
  assign RetimeWrapper_80_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24131.4]
  assign RetimeWrapper_80_io_in = _T_2667 & io_rPort_6_en_0; // @[package.scala 94:16:@24130.4]
  assign RetimeWrapper_81_clock = clock; // @[:@24136.4]
  assign RetimeWrapper_81_reset = reset; // @[:@24137.4]
  assign RetimeWrapper_81_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24139.4]
  assign RetimeWrapper_81_io_in = _T_2851 & io_rPort_6_en_0; // @[package.scala 94:16:@24138.4]
  assign RetimeWrapper_82_clock = clock; // @[:@24144.4]
  assign RetimeWrapper_82_reset = reset; // @[:@24145.4]
  assign RetimeWrapper_82_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24147.4]
  assign RetimeWrapper_82_io_in = _T_3035 & io_rPort_6_en_0; // @[package.scala 94:16:@24146.4]
  assign RetimeWrapper_83_clock = clock; // @[:@24152.4]
  assign RetimeWrapper_83_reset = reset; // @[:@24153.4]
  assign RetimeWrapper_83_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@24155.4]
  assign RetimeWrapper_83_io_in = _T_3219 & io_rPort_6_en_0; // @[package.scala 94:16:@24154.4]
  assign RetimeWrapper_84_clock = clock; // @[:@24208.4]
  assign RetimeWrapper_84_reset = reset; // @[:@24209.4]
  assign RetimeWrapper_84_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24211.4]
  assign RetimeWrapper_84_io_in = _T_1299 & io_rPort_7_en_0; // @[package.scala 94:16:@24210.4]
  assign RetimeWrapper_85_clock = clock; // @[:@24216.4]
  assign RetimeWrapper_85_reset = reset; // @[:@24217.4]
  assign RetimeWrapper_85_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24219.4]
  assign RetimeWrapper_85_io_in = _T_1483 & io_rPort_7_en_0; // @[package.scala 94:16:@24218.4]
  assign RetimeWrapper_86_clock = clock; // @[:@24224.4]
  assign RetimeWrapper_86_reset = reset; // @[:@24225.4]
  assign RetimeWrapper_86_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24227.4]
  assign RetimeWrapper_86_io_in = _T_1667 & io_rPort_7_en_0; // @[package.scala 94:16:@24226.4]
  assign RetimeWrapper_87_clock = clock; // @[:@24232.4]
  assign RetimeWrapper_87_reset = reset; // @[:@24233.4]
  assign RetimeWrapper_87_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24235.4]
  assign RetimeWrapper_87_io_in = _T_1851 & io_rPort_7_en_0; // @[package.scala 94:16:@24234.4]
  assign RetimeWrapper_88_clock = clock; // @[:@24240.4]
  assign RetimeWrapper_88_reset = reset; // @[:@24241.4]
  assign RetimeWrapper_88_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24243.4]
  assign RetimeWrapper_88_io_in = _T_2035 & io_rPort_7_en_0; // @[package.scala 94:16:@24242.4]
  assign RetimeWrapper_89_clock = clock; // @[:@24248.4]
  assign RetimeWrapper_89_reset = reset; // @[:@24249.4]
  assign RetimeWrapper_89_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24251.4]
  assign RetimeWrapper_89_io_in = _T_2219 & io_rPort_7_en_0; // @[package.scala 94:16:@24250.4]
  assign RetimeWrapper_90_clock = clock; // @[:@24256.4]
  assign RetimeWrapper_90_reset = reset; // @[:@24257.4]
  assign RetimeWrapper_90_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24259.4]
  assign RetimeWrapper_90_io_in = _T_2403 & io_rPort_7_en_0; // @[package.scala 94:16:@24258.4]
  assign RetimeWrapper_91_clock = clock; // @[:@24264.4]
  assign RetimeWrapper_91_reset = reset; // @[:@24265.4]
  assign RetimeWrapper_91_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24267.4]
  assign RetimeWrapper_91_io_in = _T_2587 & io_rPort_7_en_0; // @[package.scala 94:16:@24266.4]
  assign RetimeWrapper_92_clock = clock; // @[:@24272.4]
  assign RetimeWrapper_92_reset = reset; // @[:@24273.4]
  assign RetimeWrapper_92_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24275.4]
  assign RetimeWrapper_92_io_in = _T_2771 & io_rPort_7_en_0; // @[package.scala 94:16:@24274.4]
  assign RetimeWrapper_93_clock = clock; // @[:@24280.4]
  assign RetimeWrapper_93_reset = reset; // @[:@24281.4]
  assign RetimeWrapper_93_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24283.4]
  assign RetimeWrapper_93_io_in = _T_2955 & io_rPort_7_en_0; // @[package.scala 94:16:@24282.4]
  assign RetimeWrapper_94_clock = clock; // @[:@24288.4]
  assign RetimeWrapper_94_reset = reset; // @[:@24289.4]
  assign RetimeWrapper_94_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24291.4]
  assign RetimeWrapper_94_io_in = _T_3139 & io_rPort_7_en_0; // @[package.scala 94:16:@24290.4]
  assign RetimeWrapper_95_clock = clock; // @[:@24296.4]
  assign RetimeWrapper_95_reset = reset; // @[:@24297.4]
  assign RetimeWrapper_95_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@24299.4]
  assign RetimeWrapper_95_io_in = _T_3323 & io_rPort_7_en_0; // @[package.scala 94:16:@24298.4]
  assign RetimeWrapper_96_clock = clock; // @[:@24352.4]
  assign RetimeWrapper_96_reset = reset; // @[:@24353.4]
  assign RetimeWrapper_96_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24355.4]
  assign RetimeWrapper_96_io_in = _T_1201 & io_rPort_8_en_0; // @[package.scala 94:16:@24354.4]
  assign RetimeWrapper_97_clock = clock; // @[:@24360.4]
  assign RetimeWrapper_97_reset = reset; // @[:@24361.4]
  assign RetimeWrapper_97_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24363.4]
  assign RetimeWrapper_97_io_in = _T_1385 & io_rPort_8_en_0; // @[package.scala 94:16:@24362.4]
  assign RetimeWrapper_98_clock = clock; // @[:@24368.4]
  assign RetimeWrapper_98_reset = reset; // @[:@24369.4]
  assign RetimeWrapper_98_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24371.4]
  assign RetimeWrapper_98_io_in = _T_1569 & io_rPort_8_en_0; // @[package.scala 94:16:@24370.4]
  assign RetimeWrapper_99_clock = clock; // @[:@24376.4]
  assign RetimeWrapper_99_reset = reset; // @[:@24377.4]
  assign RetimeWrapper_99_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24379.4]
  assign RetimeWrapper_99_io_in = _T_1753 & io_rPort_8_en_0; // @[package.scala 94:16:@24378.4]
  assign RetimeWrapper_100_clock = clock; // @[:@24384.4]
  assign RetimeWrapper_100_reset = reset; // @[:@24385.4]
  assign RetimeWrapper_100_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24387.4]
  assign RetimeWrapper_100_io_in = _T_1937 & io_rPort_8_en_0; // @[package.scala 94:16:@24386.4]
  assign RetimeWrapper_101_clock = clock; // @[:@24392.4]
  assign RetimeWrapper_101_reset = reset; // @[:@24393.4]
  assign RetimeWrapper_101_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24395.4]
  assign RetimeWrapper_101_io_in = _T_2121 & io_rPort_8_en_0; // @[package.scala 94:16:@24394.4]
  assign RetimeWrapper_102_clock = clock; // @[:@24400.4]
  assign RetimeWrapper_102_reset = reset; // @[:@24401.4]
  assign RetimeWrapper_102_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24403.4]
  assign RetimeWrapper_102_io_in = _T_2305 & io_rPort_8_en_0; // @[package.scala 94:16:@24402.4]
  assign RetimeWrapper_103_clock = clock; // @[:@24408.4]
  assign RetimeWrapper_103_reset = reset; // @[:@24409.4]
  assign RetimeWrapper_103_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24411.4]
  assign RetimeWrapper_103_io_in = _T_2489 & io_rPort_8_en_0; // @[package.scala 94:16:@24410.4]
  assign RetimeWrapper_104_clock = clock; // @[:@24416.4]
  assign RetimeWrapper_104_reset = reset; // @[:@24417.4]
  assign RetimeWrapper_104_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24419.4]
  assign RetimeWrapper_104_io_in = _T_2673 & io_rPort_8_en_0; // @[package.scala 94:16:@24418.4]
  assign RetimeWrapper_105_clock = clock; // @[:@24424.4]
  assign RetimeWrapper_105_reset = reset; // @[:@24425.4]
  assign RetimeWrapper_105_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24427.4]
  assign RetimeWrapper_105_io_in = _T_2857 & io_rPort_8_en_0; // @[package.scala 94:16:@24426.4]
  assign RetimeWrapper_106_clock = clock; // @[:@24432.4]
  assign RetimeWrapper_106_reset = reset; // @[:@24433.4]
  assign RetimeWrapper_106_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24435.4]
  assign RetimeWrapper_106_io_in = _T_3041 & io_rPort_8_en_0; // @[package.scala 94:16:@24434.4]
  assign RetimeWrapper_107_clock = clock; // @[:@24440.4]
  assign RetimeWrapper_107_reset = reset; // @[:@24441.4]
  assign RetimeWrapper_107_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@24443.4]
  assign RetimeWrapper_107_io_in = _T_3225 & io_rPort_8_en_0; // @[package.scala 94:16:@24442.4]
  assign RetimeWrapper_108_clock = clock; // @[:@24496.4]
  assign RetimeWrapper_108_reset = reset; // @[:@24497.4]
  assign RetimeWrapper_108_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24499.4]
  assign RetimeWrapper_108_io_in = _T_1305 & io_rPort_9_en_0; // @[package.scala 94:16:@24498.4]
  assign RetimeWrapper_109_clock = clock; // @[:@24504.4]
  assign RetimeWrapper_109_reset = reset; // @[:@24505.4]
  assign RetimeWrapper_109_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24507.4]
  assign RetimeWrapper_109_io_in = _T_1489 & io_rPort_9_en_0; // @[package.scala 94:16:@24506.4]
  assign RetimeWrapper_110_clock = clock; // @[:@24512.4]
  assign RetimeWrapper_110_reset = reset; // @[:@24513.4]
  assign RetimeWrapper_110_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24515.4]
  assign RetimeWrapper_110_io_in = _T_1673 & io_rPort_9_en_0; // @[package.scala 94:16:@24514.4]
  assign RetimeWrapper_111_clock = clock; // @[:@24520.4]
  assign RetimeWrapper_111_reset = reset; // @[:@24521.4]
  assign RetimeWrapper_111_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24523.4]
  assign RetimeWrapper_111_io_in = _T_1857 & io_rPort_9_en_0; // @[package.scala 94:16:@24522.4]
  assign RetimeWrapper_112_clock = clock; // @[:@24528.4]
  assign RetimeWrapper_112_reset = reset; // @[:@24529.4]
  assign RetimeWrapper_112_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24531.4]
  assign RetimeWrapper_112_io_in = _T_2041 & io_rPort_9_en_0; // @[package.scala 94:16:@24530.4]
  assign RetimeWrapper_113_clock = clock; // @[:@24536.4]
  assign RetimeWrapper_113_reset = reset; // @[:@24537.4]
  assign RetimeWrapper_113_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24539.4]
  assign RetimeWrapper_113_io_in = _T_2225 & io_rPort_9_en_0; // @[package.scala 94:16:@24538.4]
  assign RetimeWrapper_114_clock = clock; // @[:@24544.4]
  assign RetimeWrapper_114_reset = reset; // @[:@24545.4]
  assign RetimeWrapper_114_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24547.4]
  assign RetimeWrapper_114_io_in = _T_2409 & io_rPort_9_en_0; // @[package.scala 94:16:@24546.4]
  assign RetimeWrapper_115_clock = clock; // @[:@24552.4]
  assign RetimeWrapper_115_reset = reset; // @[:@24553.4]
  assign RetimeWrapper_115_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24555.4]
  assign RetimeWrapper_115_io_in = _T_2593 & io_rPort_9_en_0; // @[package.scala 94:16:@24554.4]
  assign RetimeWrapper_116_clock = clock; // @[:@24560.4]
  assign RetimeWrapper_116_reset = reset; // @[:@24561.4]
  assign RetimeWrapper_116_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24563.4]
  assign RetimeWrapper_116_io_in = _T_2777 & io_rPort_9_en_0; // @[package.scala 94:16:@24562.4]
  assign RetimeWrapper_117_clock = clock; // @[:@24568.4]
  assign RetimeWrapper_117_reset = reset; // @[:@24569.4]
  assign RetimeWrapper_117_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24571.4]
  assign RetimeWrapper_117_io_in = _T_2961 & io_rPort_9_en_0; // @[package.scala 94:16:@24570.4]
  assign RetimeWrapper_118_clock = clock; // @[:@24576.4]
  assign RetimeWrapper_118_reset = reset; // @[:@24577.4]
  assign RetimeWrapper_118_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24579.4]
  assign RetimeWrapper_118_io_in = _T_3145 & io_rPort_9_en_0; // @[package.scala 94:16:@24578.4]
  assign RetimeWrapper_119_clock = clock; // @[:@24584.4]
  assign RetimeWrapper_119_reset = reset; // @[:@24585.4]
  assign RetimeWrapper_119_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@24587.4]
  assign RetimeWrapper_119_io_in = _T_3329 & io_rPort_9_en_0; // @[package.scala 94:16:@24586.4]
  assign RetimeWrapper_120_clock = clock; // @[:@24640.4]
  assign RetimeWrapper_120_reset = reset; // @[:@24641.4]
  assign RetimeWrapper_120_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24643.4]
  assign RetimeWrapper_120_io_in = _T_1207 & io_rPort_10_en_0; // @[package.scala 94:16:@24642.4]
  assign RetimeWrapper_121_clock = clock; // @[:@24648.4]
  assign RetimeWrapper_121_reset = reset; // @[:@24649.4]
  assign RetimeWrapper_121_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24651.4]
  assign RetimeWrapper_121_io_in = _T_1391 & io_rPort_10_en_0; // @[package.scala 94:16:@24650.4]
  assign RetimeWrapper_122_clock = clock; // @[:@24656.4]
  assign RetimeWrapper_122_reset = reset; // @[:@24657.4]
  assign RetimeWrapper_122_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24659.4]
  assign RetimeWrapper_122_io_in = _T_1575 & io_rPort_10_en_0; // @[package.scala 94:16:@24658.4]
  assign RetimeWrapper_123_clock = clock; // @[:@24664.4]
  assign RetimeWrapper_123_reset = reset; // @[:@24665.4]
  assign RetimeWrapper_123_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24667.4]
  assign RetimeWrapper_123_io_in = _T_1759 & io_rPort_10_en_0; // @[package.scala 94:16:@24666.4]
  assign RetimeWrapper_124_clock = clock; // @[:@24672.4]
  assign RetimeWrapper_124_reset = reset; // @[:@24673.4]
  assign RetimeWrapper_124_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24675.4]
  assign RetimeWrapper_124_io_in = _T_1943 & io_rPort_10_en_0; // @[package.scala 94:16:@24674.4]
  assign RetimeWrapper_125_clock = clock; // @[:@24680.4]
  assign RetimeWrapper_125_reset = reset; // @[:@24681.4]
  assign RetimeWrapper_125_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24683.4]
  assign RetimeWrapper_125_io_in = _T_2127 & io_rPort_10_en_0; // @[package.scala 94:16:@24682.4]
  assign RetimeWrapper_126_clock = clock; // @[:@24688.4]
  assign RetimeWrapper_126_reset = reset; // @[:@24689.4]
  assign RetimeWrapper_126_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24691.4]
  assign RetimeWrapper_126_io_in = _T_2311 & io_rPort_10_en_0; // @[package.scala 94:16:@24690.4]
  assign RetimeWrapper_127_clock = clock; // @[:@24696.4]
  assign RetimeWrapper_127_reset = reset; // @[:@24697.4]
  assign RetimeWrapper_127_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24699.4]
  assign RetimeWrapper_127_io_in = _T_2495 & io_rPort_10_en_0; // @[package.scala 94:16:@24698.4]
  assign RetimeWrapper_128_clock = clock; // @[:@24704.4]
  assign RetimeWrapper_128_reset = reset; // @[:@24705.4]
  assign RetimeWrapper_128_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24707.4]
  assign RetimeWrapper_128_io_in = _T_2679 & io_rPort_10_en_0; // @[package.scala 94:16:@24706.4]
  assign RetimeWrapper_129_clock = clock; // @[:@24712.4]
  assign RetimeWrapper_129_reset = reset; // @[:@24713.4]
  assign RetimeWrapper_129_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24715.4]
  assign RetimeWrapper_129_io_in = _T_2863 & io_rPort_10_en_0; // @[package.scala 94:16:@24714.4]
  assign RetimeWrapper_130_clock = clock; // @[:@24720.4]
  assign RetimeWrapper_130_reset = reset; // @[:@24721.4]
  assign RetimeWrapper_130_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24723.4]
  assign RetimeWrapper_130_io_in = _T_3047 & io_rPort_10_en_0; // @[package.scala 94:16:@24722.4]
  assign RetimeWrapper_131_clock = clock; // @[:@24728.4]
  assign RetimeWrapper_131_reset = reset; // @[:@24729.4]
  assign RetimeWrapper_131_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@24731.4]
  assign RetimeWrapper_131_io_in = _T_3231 & io_rPort_10_en_0; // @[package.scala 94:16:@24730.4]
  assign RetimeWrapper_132_clock = clock; // @[:@24784.4]
  assign RetimeWrapper_132_reset = reset; // @[:@24785.4]
  assign RetimeWrapper_132_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24787.4]
  assign RetimeWrapper_132_io_in = _T_1311 & io_rPort_11_en_0; // @[package.scala 94:16:@24786.4]
  assign RetimeWrapper_133_clock = clock; // @[:@24792.4]
  assign RetimeWrapper_133_reset = reset; // @[:@24793.4]
  assign RetimeWrapper_133_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24795.4]
  assign RetimeWrapper_133_io_in = _T_1495 & io_rPort_11_en_0; // @[package.scala 94:16:@24794.4]
  assign RetimeWrapper_134_clock = clock; // @[:@24800.4]
  assign RetimeWrapper_134_reset = reset; // @[:@24801.4]
  assign RetimeWrapper_134_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24803.4]
  assign RetimeWrapper_134_io_in = _T_1679 & io_rPort_11_en_0; // @[package.scala 94:16:@24802.4]
  assign RetimeWrapper_135_clock = clock; // @[:@24808.4]
  assign RetimeWrapper_135_reset = reset; // @[:@24809.4]
  assign RetimeWrapper_135_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24811.4]
  assign RetimeWrapper_135_io_in = _T_1863 & io_rPort_11_en_0; // @[package.scala 94:16:@24810.4]
  assign RetimeWrapper_136_clock = clock; // @[:@24816.4]
  assign RetimeWrapper_136_reset = reset; // @[:@24817.4]
  assign RetimeWrapper_136_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24819.4]
  assign RetimeWrapper_136_io_in = _T_2047 & io_rPort_11_en_0; // @[package.scala 94:16:@24818.4]
  assign RetimeWrapper_137_clock = clock; // @[:@24824.4]
  assign RetimeWrapper_137_reset = reset; // @[:@24825.4]
  assign RetimeWrapper_137_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24827.4]
  assign RetimeWrapper_137_io_in = _T_2231 & io_rPort_11_en_0; // @[package.scala 94:16:@24826.4]
  assign RetimeWrapper_138_clock = clock; // @[:@24832.4]
  assign RetimeWrapper_138_reset = reset; // @[:@24833.4]
  assign RetimeWrapper_138_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24835.4]
  assign RetimeWrapper_138_io_in = _T_2415 & io_rPort_11_en_0; // @[package.scala 94:16:@24834.4]
  assign RetimeWrapper_139_clock = clock; // @[:@24840.4]
  assign RetimeWrapper_139_reset = reset; // @[:@24841.4]
  assign RetimeWrapper_139_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24843.4]
  assign RetimeWrapper_139_io_in = _T_2599 & io_rPort_11_en_0; // @[package.scala 94:16:@24842.4]
  assign RetimeWrapper_140_clock = clock; // @[:@24848.4]
  assign RetimeWrapper_140_reset = reset; // @[:@24849.4]
  assign RetimeWrapper_140_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24851.4]
  assign RetimeWrapper_140_io_in = _T_2783 & io_rPort_11_en_0; // @[package.scala 94:16:@24850.4]
  assign RetimeWrapper_141_clock = clock; // @[:@24856.4]
  assign RetimeWrapper_141_reset = reset; // @[:@24857.4]
  assign RetimeWrapper_141_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24859.4]
  assign RetimeWrapper_141_io_in = _T_2967 & io_rPort_11_en_0; // @[package.scala 94:16:@24858.4]
  assign RetimeWrapper_142_clock = clock; // @[:@24864.4]
  assign RetimeWrapper_142_reset = reset; // @[:@24865.4]
  assign RetimeWrapper_142_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24867.4]
  assign RetimeWrapper_142_io_in = _T_3151 & io_rPort_11_en_0; // @[package.scala 94:16:@24866.4]
  assign RetimeWrapper_143_clock = clock; // @[:@24872.4]
  assign RetimeWrapper_143_reset = reset; // @[:@24873.4]
  assign RetimeWrapper_143_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24875.4]
  assign RetimeWrapper_143_io_in = _T_3335 & io_rPort_11_en_0; // @[package.scala 94:16:@24874.4]
  assign RetimeWrapper_144_clock = clock; // @[:@24928.4]
  assign RetimeWrapper_144_reset = reset; // @[:@24929.4]
  assign RetimeWrapper_144_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24931.4]
  assign RetimeWrapper_144_io_in = _T_1213 & io_rPort_12_en_0; // @[package.scala 94:16:@24930.4]
  assign RetimeWrapper_145_clock = clock; // @[:@24936.4]
  assign RetimeWrapper_145_reset = reset; // @[:@24937.4]
  assign RetimeWrapper_145_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24939.4]
  assign RetimeWrapper_145_io_in = _T_1397 & io_rPort_12_en_0; // @[package.scala 94:16:@24938.4]
  assign RetimeWrapper_146_clock = clock; // @[:@24944.4]
  assign RetimeWrapper_146_reset = reset; // @[:@24945.4]
  assign RetimeWrapper_146_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24947.4]
  assign RetimeWrapper_146_io_in = _T_1581 & io_rPort_12_en_0; // @[package.scala 94:16:@24946.4]
  assign RetimeWrapper_147_clock = clock; // @[:@24952.4]
  assign RetimeWrapper_147_reset = reset; // @[:@24953.4]
  assign RetimeWrapper_147_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24955.4]
  assign RetimeWrapper_147_io_in = _T_1765 & io_rPort_12_en_0; // @[package.scala 94:16:@24954.4]
  assign RetimeWrapper_148_clock = clock; // @[:@24960.4]
  assign RetimeWrapper_148_reset = reset; // @[:@24961.4]
  assign RetimeWrapper_148_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24963.4]
  assign RetimeWrapper_148_io_in = _T_1949 & io_rPort_12_en_0; // @[package.scala 94:16:@24962.4]
  assign RetimeWrapper_149_clock = clock; // @[:@24968.4]
  assign RetimeWrapper_149_reset = reset; // @[:@24969.4]
  assign RetimeWrapper_149_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24971.4]
  assign RetimeWrapper_149_io_in = _T_2133 & io_rPort_12_en_0; // @[package.scala 94:16:@24970.4]
  assign RetimeWrapper_150_clock = clock; // @[:@24976.4]
  assign RetimeWrapper_150_reset = reset; // @[:@24977.4]
  assign RetimeWrapper_150_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24979.4]
  assign RetimeWrapper_150_io_in = _T_2317 & io_rPort_12_en_0; // @[package.scala 94:16:@24978.4]
  assign RetimeWrapper_151_clock = clock; // @[:@24984.4]
  assign RetimeWrapper_151_reset = reset; // @[:@24985.4]
  assign RetimeWrapper_151_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24987.4]
  assign RetimeWrapper_151_io_in = _T_2501 & io_rPort_12_en_0; // @[package.scala 94:16:@24986.4]
  assign RetimeWrapper_152_clock = clock; // @[:@24992.4]
  assign RetimeWrapper_152_reset = reset; // @[:@24993.4]
  assign RetimeWrapper_152_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24995.4]
  assign RetimeWrapper_152_io_in = _T_2685 & io_rPort_12_en_0; // @[package.scala 94:16:@24994.4]
  assign RetimeWrapper_153_clock = clock; // @[:@25000.4]
  assign RetimeWrapper_153_reset = reset; // @[:@25001.4]
  assign RetimeWrapper_153_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@25003.4]
  assign RetimeWrapper_153_io_in = _T_2869 & io_rPort_12_en_0; // @[package.scala 94:16:@25002.4]
  assign RetimeWrapper_154_clock = clock; // @[:@25008.4]
  assign RetimeWrapper_154_reset = reset; // @[:@25009.4]
  assign RetimeWrapper_154_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@25011.4]
  assign RetimeWrapper_154_io_in = _T_3053 & io_rPort_12_en_0; // @[package.scala 94:16:@25010.4]
  assign RetimeWrapper_155_clock = clock; // @[:@25016.4]
  assign RetimeWrapper_155_reset = reset; // @[:@25017.4]
  assign RetimeWrapper_155_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@25019.4]
  assign RetimeWrapper_155_io_in = _T_3237 & io_rPort_12_en_0; // @[package.scala 94:16:@25018.4]
  assign RetimeWrapper_156_clock = clock; // @[:@25072.4]
  assign RetimeWrapper_156_reset = reset; // @[:@25073.4]
  assign RetimeWrapper_156_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25075.4]
  assign RetimeWrapper_156_io_in = _T_1317 & io_rPort_13_en_0; // @[package.scala 94:16:@25074.4]
  assign RetimeWrapper_157_clock = clock; // @[:@25080.4]
  assign RetimeWrapper_157_reset = reset; // @[:@25081.4]
  assign RetimeWrapper_157_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25083.4]
  assign RetimeWrapper_157_io_in = _T_1501 & io_rPort_13_en_0; // @[package.scala 94:16:@25082.4]
  assign RetimeWrapper_158_clock = clock; // @[:@25088.4]
  assign RetimeWrapper_158_reset = reset; // @[:@25089.4]
  assign RetimeWrapper_158_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25091.4]
  assign RetimeWrapper_158_io_in = _T_1685 & io_rPort_13_en_0; // @[package.scala 94:16:@25090.4]
  assign RetimeWrapper_159_clock = clock; // @[:@25096.4]
  assign RetimeWrapper_159_reset = reset; // @[:@25097.4]
  assign RetimeWrapper_159_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25099.4]
  assign RetimeWrapper_159_io_in = _T_1869 & io_rPort_13_en_0; // @[package.scala 94:16:@25098.4]
  assign RetimeWrapper_160_clock = clock; // @[:@25104.4]
  assign RetimeWrapper_160_reset = reset; // @[:@25105.4]
  assign RetimeWrapper_160_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25107.4]
  assign RetimeWrapper_160_io_in = _T_2053 & io_rPort_13_en_0; // @[package.scala 94:16:@25106.4]
  assign RetimeWrapper_161_clock = clock; // @[:@25112.4]
  assign RetimeWrapper_161_reset = reset; // @[:@25113.4]
  assign RetimeWrapper_161_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25115.4]
  assign RetimeWrapper_161_io_in = _T_2237 & io_rPort_13_en_0; // @[package.scala 94:16:@25114.4]
  assign RetimeWrapper_162_clock = clock; // @[:@25120.4]
  assign RetimeWrapper_162_reset = reset; // @[:@25121.4]
  assign RetimeWrapper_162_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25123.4]
  assign RetimeWrapper_162_io_in = _T_2421 & io_rPort_13_en_0; // @[package.scala 94:16:@25122.4]
  assign RetimeWrapper_163_clock = clock; // @[:@25128.4]
  assign RetimeWrapper_163_reset = reset; // @[:@25129.4]
  assign RetimeWrapper_163_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25131.4]
  assign RetimeWrapper_163_io_in = _T_2605 & io_rPort_13_en_0; // @[package.scala 94:16:@25130.4]
  assign RetimeWrapper_164_clock = clock; // @[:@25136.4]
  assign RetimeWrapper_164_reset = reset; // @[:@25137.4]
  assign RetimeWrapper_164_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25139.4]
  assign RetimeWrapper_164_io_in = _T_2789 & io_rPort_13_en_0; // @[package.scala 94:16:@25138.4]
  assign RetimeWrapper_165_clock = clock; // @[:@25144.4]
  assign RetimeWrapper_165_reset = reset; // @[:@25145.4]
  assign RetimeWrapper_165_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25147.4]
  assign RetimeWrapper_165_io_in = _T_2973 & io_rPort_13_en_0; // @[package.scala 94:16:@25146.4]
  assign RetimeWrapper_166_clock = clock; // @[:@25152.4]
  assign RetimeWrapper_166_reset = reset; // @[:@25153.4]
  assign RetimeWrapper_166_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25155.4]
  assign RetimeWrapper_166_io_in = _T_3157 & io_rPort_13_en_0; // @[package.scala 94:16:@25154.4]
  assign RetimeWrapper_167_clock = clock; // @[:@25160.4]
  assign RetimeWrapper_167_reset = reset; // @[:@25161.4]
  assign RetimeWrapper_167_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@25163.4]
  assign RetimeWrapper_167_io_in = _T_3341 & io_rPort_13_en_0; // @[package.scala 94:16:@25162.4]
  assign RetimeWrapper_168_clock = clock; // @[:@25216.4]
  assign RetimeWrapper_168_reset = reset; // @[:@25217.4]
  assign RetimeWrapper_168_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25219.4]
  assign RetimeWrapper_168_io_in = _T_1323 & io_rPort_14_en_0; // @[package.scala 94:16:@25218.4]
  assign RetimeWrapper_169_clock = clock; // @[:@25224.4]
  assign RetimeWrapper_169_reset = reset; // @[:@25225.4]
  assign RetimeWrapper_169_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25227.4]
  assign RetimeWrapper_169_io_in = _T_1507 & io_rPort_14_en_0; // @[package.scala 94:16:@25226.4]
  assign RetimeWrapper_170_clock = clock; // @[:@25232.4]
  assign RetimeWrapper_170_reset = reset; // @[:@25233.4]
  assign RetimeWrapper_170_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25235.4]
  assign RetimeWrapper_170_io_in = _T_1691 & io_rPort_14_en_0; // @[package.scala 94:16:@25234.4]
  assign RetimeWrapper_171_clock = clock; // @[:@25240.4]
  assign RetimeWrapper_171_reset = reset; // @[:@25241.4]
  assign RetimeWrapper_171_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25243.4]
  assign RetimeWrapper_171_io_in = _T_1875 & io_rPort_14_en_0; // @[package.scala 94:16:@25242.4]
  assign RetimeWrapper_172_clock = clock; // @[:@25248.4]
  assign RetimeWrapper_172_reset = reset; // @[:@25249.4]
  assign RetimeWrapper_172_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25251.4]
  assign RetimeWrapper_172_io_in = _T_2059 & io_rPort_14_en_0; // @[package.scala 94:16:@25250.4]
  assign RetimeWrapper_173_clock = clock; // @[:@25256.4]
  assign RetimeWrapper_173_reset = reset; // @[:@25257.4]
  assign RetimeWrapper_173_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25259.4]
  assign RetimeWrapper_173_io_in = _T_2243 & io_rPort_14_en_0; // @[package.scala 94:16:@25258.4]
  assign RetimeWrapper_174_clock = clock; // @[:@25264.4]
  assign RetimeWrapper_174_reset = reset; // @[:@25265.4]
  assign RetimeWrapper_174_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25267.4]
  assign RetimeWrapper_174_io_in = _T_2427 & io_rPort_14_en_0; // @[package.scala 94:16:@25266.4]
  assign RetimeWrapper_175_clock = clock; // @[:@25272.4]
  assign RetimeWrapper_175_reset = reset; // @[:@25273.4]
  assign RetimeWrapper_175_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25275.4]
  assign RetimeWrapper_175_io_in = _T_2611 & io_rPort_14_en_0; // @[package.scala 94:16:@25274.4]
  assign RetimeWrapper_176_clock = clock; // @[:@25280.4]
  assign RetimeWrapper_176_reset = reset; // @[:@25281.4]
  assign RetimeWrapper_176_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25283.4]
  assign RetimeWrapper_176_io_in = _T_2795 & io_rPort_14_en_0; // @[package.scala 94:16:@25282.4]
  assign RetimeWrapper_177_clock = clock; // @[:@25288.4]
  assign RetimeWrapper_177_reset = reset; // @[:@25289.4]
  assign RetimeWrapper_177_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25291.4]
  assign RetimeWrapper_177_io_in = _T_2979 & io_rPort_14_en_0; // @[package.scala 94:16:@25290.4]
  assign RetimeWrapper_178_clock = clock; // @[:@25296.4]
  assign RetimeWrapper_178_reset = reset; // @[:@25297.4]
  assign RetimeWrapper_178_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25299.4]
  assign RetimeWrapper_178_io_in = _T_3163 & io_rPort_14_en_0; // @[package.scala 94:16:@25298.4]
  assign RetimeWrapper_179_clock = clock; // @[:@25304.4]
  assign RetimeWrapper_179_reset = reset; // @[:@25305.4]
  assign RetimeWrapper_179_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@25307.4]
  assign RetimeWrapper_179_io_in = _T_3347 & io_rPort_14_en_0; // @[package.scala 94:16:@25306.4]
  assign RetimeWrapper_180_clock = clock; // @[:@25360.4]
  assign RetimeWrapper_180_reset = reset; // @[:@25361.4]
  assign RetimeWrapper_180_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25363.4]
  assign RetimeWrapper_180_io_in = _T_1219 & io_rPort_15_en_0; // @[package.scala 94:16:@25362.4]
  assign RetimeWrapper_181_clock = clock; // @[:@25368.4]
  assign RetimeWrapper_181_reset = reset; // @[:@25369.4]
  assign RetimeWrapper_181_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25371.4]
  assign RetimeWrapper_181_io_in = _T_1403 & io_rPort_15_en_0; // @[package.scala 94:16:@25370.4]
  assign RetimeWrapper_182_clock = clock; // @[:@25376.4]
  assign RetimeWrapper_182_reset = reset; // @[:@25377.4]
  assign RetimeWrapper_182_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25379.4]
  assign RetimeWrapper_182_io_in = _T_1587 & io_rPort_15_en_0; // @[package.scala 94:16:@25378.4]
  assign RetimeWrapper_183_clock = clock; // @[:@25384.4]
  assign RetimeWrapper_183_reset = reset; // @[:@25385.4]
  assign RetimeWrapper_183_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25387.4]
  assign RetimeWrapper_183_io_in = _T_1771 & io_rPort_15_en_0; // @[package.scala 94:16:@25386.4]
  assign RetimeWrapper_184_clock = clock; // @[:@25392.4]
  assign RetimeWrapper_184_reset = reset; // @[:@25393.4]
  assign RetimeWrapper_184_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25395.4]
  assign RetimeWrapper_184_io_in = _T_1955 & io_rPort_15_en_0; // @[package.scala 94:16:@25394.4]
  assign RetimeWrapper_185_clock = clock; // @[:@25400.4]
  assign RetimeWrapper_185_reset = reset; // @[:@25401.4]
  assign RetimeWrapper_185_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25403.4]
  assign RetimeWrapper_185_io_in = _T_2139 & io_rPort_15_en_0; // @[package.scala 94:16:@25402.4]
  assign RetimeWrapper_186_clock = clock; // @[:@25408.4]
  assign RetimeWrapper_186_reset = reset; // @[:@25409.4]
  assign RetimeWrapper_186_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25411.4]
  assign RetimeWrapper_186_io_in = _T_2323 & io_rPort_15_en_0; // @[package.scala 94:16:@25410.4]
  assign RetimeWrapper_187_clock = clock; // @[:@25416.4]
  assign RetimeWrapper_187_reset = reset; // @[:@25417.4]
  assign RetimeWrapper_187_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25419.4]
  assign RetimeWrapper_187_io_in = _T_2507 & io_rPort_15_en_0; // @[package.scala 94:16:@25418.4]
  assign RetimeWrapper_188_clock = clock; // @[:@25424.4]
  assign RetimeWrapper_188_reset = reset; // @[:@25425.4]
  assign RetimeWrapper_188_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25427.4]
  assign RetimeWrapper_188_io_in = _T_2691 & io_rPort_15_en_0; // @[package.scala 94:16:@25426.4]
  assign RetimeWrapper_189_clock = clock; // @[:@25432.4]
  assign RetimeWrapper_189_reset = reset; // @[:@25433.4]
  assign RetimeWrapper_189_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25435.4]
  assign RetimeWrapper_189_io_in = _T_2875 & io_rPort_15_en_0; // @[package.scala 94:16:@25434.4]
  assign RetimeWrapper_190_clock = clock; // @[:@25440.4]
  assign RetimeWrapper_190_reset = reset; // @[:@25441.4]
  assign RetimeWrapper_190_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25443.4]
  assign RetimeWrapper_190_io_in = _T_3059 & io_rPort_15_en_0; // @[package.scala 94:16:@25442.4]
  assign RetimeWrapper_191_clock = clock; // @[:@25448.4]
  assign RetimeWrapper_191_reset = reset; // @[:@25449.4]
  assign RetimeWrapper_191_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@25451.4]
  assign RetimeWrapper_191_io_in = _T_3243 & io_rPort_15_en_0; // @[package.scala 94:16:@25450.4]
  assign RetimeWrapper_192_clock = clock; // @[:@25504.4]
  assign RetimeWrapper_192_reset = reset; // @[:@25505.4]
  assign RetimeWrapper_192_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25507.4]
  assign RetimeWrapper_192_io_in = _T_1225 & io_rPort_16_en_0; // @[package.scala 94:16:@25506.4]
  assign RetimeWrapper_193_clock = clock; // @[:@25512.4]
  assign RetimeWrapper_193_reset = reset; // @[:@25513.4]
  assign RetimeWrapper_193_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25515.4]
  assign RetimeWrapper_193_io_in = _T_1409 & io_rPort_16_en_0; // @[package.scala 94:16:@25514.4]
  assign RetimeWrapper_194_clock = clock; // @[:@25520.4]
  assign RetimeWrapper_194_reset = reset; // @[:@25521.4]
  assign RetimeWrapper_194_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25523.4]
  assign RetimeWrapper_194_io_in = _T_1593 & io_rPort_16_en_0; // @[package.scala 94:16:@25522.4]
  assign RetimeWrapper_195_clock = clock; // @[:@25528.4]
  assign RetimeWrapper_195_reset = reset; // @[:@25529.4]
  assign RetimeWrapper_195_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25531.4]
  assign RetimeWrapper_195_io_in = _T_1777 & io_rPort_16_en_0; // @[package.scala 94:16:@25530.4]
  assign RetimeWrapper_196_clock = clock; // @[:@25536.4]
  assign RetimeWrapper_196_reset = reset; // @[:@25537.4]
  assign RetimeWrapper_196_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25539.4]
  assign RetimeWrapper_196_io_in = _T_1961 & io_rPort_16_en_0; // @[package.scala 94:16:@25538.4]
  assign RetimeWrapper_197_clock = clock; // @[:@25544.4]
  assign RetimeWrapper_197_reset = reset; // @[:@25545.4]
  assign RetimeWrapper_197_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25547.4]
  assign RetimeWrapper_197_io_in = _T_2145 & io_rPort_16_en_0; // @[package.scala 94:16:@25546.4]
  assign RetimeWrapper_198_clock = clock; // @[:@25552.4]
  assign RetimeWrapper_198_reset = reset; // @[:@25553.4]
  assign RetimeWrapper_198_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25555.4]
  assign RetimeWrapper_198_io_in = _T_2329 & io_rPort_16_en_0; // @[package.scala 94:16:@25554.4]
  assign RetimeWrapper_199_clock = clock; // @[:@25560.4]
  assign RetimeWrapper_199_reset = reset; // @[:@25561.4]
  assign RetimeWrapper_199_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25563.4]
  assign RetimeWrapper_199_io_in = _T_2513 & io_rPort_16_en_0; // @[package.scala 94:16:@25562.4]
  assign RetimeWrapper_200_clock = clock; // @[:@25568.4]
  assign RetimeWrapper_200_reset = reset; // @[:@25569.4]
  assign RetimeWrapper_200_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25571.4]
  assign RetimeWrapper_200_io_in = _T_2697 & io_rPort_16_en_0; // @[package.scala 94:16:@25570.4]
  assign RetimeWrapper_201_clock = clock; // @[:@25576.4]
  assign RetimeWrapper_201_reset = reset; // @[:@25577.4]
  assign RetimeWrapper_201_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25579.4]
  assign RetimeWrapper_201_io_in = _T_2881 & io_rPort_16_en_0; // @[package.scala 94:16:@25578.4]
  assign RetimeWrapper_202_clock = clock; // @[:@25584.4]
  assign RetimeWrapper_202_reset = reset; // @[:@25585.4]
  assign RetimeWrapper_202_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25587.4]
  assign RetimeWrapper_202_io_in = _T_3065 & io_rPort_16_en_0; // @[package.scala 94:16:@25586.4]
  assign RetimeWrapper_203_clock = clock; // @[:@25592.4]
  assign RetimeWrapper_203_reset = reset; // @[:@25593.4]
  assign RetimeWrapper_203_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@25595.4]
  assign RetimeWrapper_203_io_in = _T_3249 & io_rPort_16_en_0; // @[package.scala 94:16:@25594.4]
  assign RetimeWrapper_204_clock = clock; // @[:@25648.4]
  assign RetimeWrapper_204_reset = reset; // @[:@25649.4]
  assign RetimeWrapper_204_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25651.4]
  assign RetimeWrapper_204_io_in = _T_1231 & io_rPort_17_en_0; // @[package.scala 94:16:@25650.4]
  assign RetimeWrapper_205_clock = clock; // @[:@25656.4]
  assign RetimeWrapper_205_reset = reset; // @[:@25657.4]
  assign RetimeWrapper_205_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25659.4]
  assign RetimeWrapper_205_io_in = _T_1415 & io_rPort_17_en_0; // @[package.scala 94:16:@25658.4]
  assign RetimeWrapper_206_clock = clock; // @[:@25664.4]
  assign RetimeWrapper_206_reset = reset; // @[:@25665.4]
  assign RetimeWrapper_206_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25667.4]
  assign RetimeWrapper_206_io_in = _T_1599 & io_rPort_17_en_0; // @[package.scala 94:16:@25666.4]
  assign RetimeWrapper_207_clock = clock; // @[:@25672.4]
  assign RetimeWrapper_207_reset = reset; // @[:@25673.4]
  assign RetimeWrapper_207_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25675.4]
  assign RetimeWrapper_207_io_in = _T_1783 & io_rPort_17_en_0; // @[package.scala 94:16:@25674.4]
  assign RetimeWrapper_208_clock = clock; // @[:@25680.4]
  assign RetimeWrapper_208_reset = reset; // @[:@25681.4]
  assign RetimeWrapper_208_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25683.4]
  assign RetimeWrapper_208_io_in = _T_1967 & io_rPort_17_en_0; // @[package.scala 94:16:@25682.4]
  assign RetimeWrapper_209_clock = clock; // @[:@25688.4]
  assign RetimeWrapper_209_reset = reset; // @[:@25689.4]
  assign RetimeWrapper_209_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25691.4]
  assign RetimeWrapper_209_io_in = _T_2151 & io_rPort_17_en_0; // @[package.scala 94:16:@25690.4]
  assign RetimeWrapper_210_clock = clock; // @[:@25696.4]
  assign RetimeWrapper_210_reset = reset; // @[:@25697.4]
  assign RetimeWrapper_210_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25699.4]
  assign RetimeWrapper_210_io_in = _T_2335 & io_rPort_17_en_0; // @[package.scala 94:16:@25698.4]
  assign RetimeWrapper_211_clock = clock; // @[:@25704.4]
  assign RetimeWrapper_211_reset = reset; // @[:@25705.4]
  assign RetimeWrapper_211_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25707.4]
  assign RetimeWrapper_211_io_in = _T_2519 & io_rPort_17_en_0; // @[package.scala 94:16:@25706.4]
  assign RetimeWrapper_212_clock = clock; // @[:@25712.4]
  assign RetimeWrapper_212_reset = reset; // @[:@25713.4]
  assign RetimeWrapper_212_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25715.4]
  assign RetimeWrapper_212_io_in = _T_2703 & io_rPort_17_en_0; // @[package.scala 94:16:@25714.4]
  assign RetimeWrapper_213_clock = clock; // @[:@25720.4]
  assign RetimeWrapper_213_reset = reset; // @[:@25721.4]
  assign RetimeWrapper_213_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25723.4]
  assign RetimeWrapper_213_io_in = _T_2887 & io_rPort_17_en_0; // @[package.scala 94:16:@25722.4]
  assign RetimeWrapper_214_clock = clock; // @[:@25728.4]
  assign RetimeWrapper_214_reset = reset; // @[:@25729.4]
  assign RetimeWrapper_214_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25731.4]
  assign RetimeWrapper_214_io_in = _T_3071 & io_rPort_17_en_0; // @[package.scala 94:16:@25730.4]
  assign RetimeWrapper_215_clock = clock; // @[:@25736.4]
  assign RetimeWrapper_215_reset = reset; // @[:@25737.4]
  assign RetimeWrapper_215_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@25739.4]
  assign RetimeWrapper_215_io_in = _T_3255 & io_rPort_17_en_0; // @[package.scala 94:16:@25738.4]
endmodule
module Modulo( // @[:@25768.2]
  input         clock, // @[:@25769.4]
  input         io_flow, // @[:@25771.4]
  input  [31:0] io_dividend, // @[:@25771.4]
  input  [31:0] io_divisor, // @[:@25771.4]
  output [31:0] io_out // @[:@25771.4]
);
  wire [31:0] m_m_axis_dout_tdata; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  wire  m_m_axis_dout_tvalid; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  wire [31:0] m_s_axis_divisor_tdata; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  wire  m_s_axis_divisor_tvalid; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  wire [31:0] m_s_axis_dividend_tdata; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  wire  m_s_axis_dividend_tvalid; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  wire  m_aclken; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  wire  m_aclk; // @[ZynqBlackBoxes.scala 48:19:@25773.4]
  div_32_32_16_Unsigned_Remainder m ( // @[ZynqBlackBoxes.scala 48:19:@25773.4]
    .m_axis_dout_tdata(m_m_axis_dout_tdata),
    .m_axis_dout_tvalid(m_m_axis_dout_tvalid),
    .s_axis_divisor_tdata(m_s_axis_divisor_tdata),
    .s_axis_divisor_tvalid(m_s_axis_divisor_tvalid),
    .s_axis_dividend_tdata(m_s_axis_dividend_tdata),
    .s_axis_dividend_tvalid(m_s_axis_dividend_tvalid),
    .aclken(m_aclken),
    .aclk(m_aclk)
  );
  assign io_out = m_m_axis_dout_tdata; // @[ZynqBlackBoxes.scala 56:12:@25789.4]
  assign m_s_axis_divisor_tdata = io_divisor; // @[ZynqBlackBoxes.scala 54:31:@25787.4]
  assign m_s_axis_divisor_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 53:32:@25786.4]
  assign m_s_axis_dividend_tdata = io_dividend; // @[ZynqBlackBoxes.scala 52:32:@25785.4]
  assign m_s_axis_dividend_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 51:33:@25784.4]
  assign m_aclken = io_flow; // @[ZynqBlackBoxes.scala 50:17:@25783.4 ZynqBlackBoxes.scala 55:17:@25788.4]
  assign m_aclk = clock; // @[ZynqBlackBoxes.scala 49:15:@25782.4]
endmodule
module fix2fixBox_38( // @[:@25791.2]
  input  [63:0] io_a, // @[:@25794.4]
  output [31:0] io_b // @[:@25794.4]
);
  assign io_b = io_a[31:0]; // @[Converter.scala 95:38:@25807.4]
endmodule
module x339( // @[:@25809.2]
  input         clock, // @[:@25810.4]
  input  [31:0] io_a, // @[:@25812.4]
  input         io_flow, // @[:@25812.4]
  output [31:0] io_result // @[:@25812.4]
);
  wire  x339_clock; // @[BigIPZynq.scala 35:21:@25820.4]
  wire  x339_io_flow; // @[BigIPZynq.scala 35:21:@25820.4]
  wire [31:0] x339_io_dividend; // @[BigIPZynq.scala 35:21:@25820.4]
  wire [31:0] x339_io_divisor; // @[BigIPZynq.scala 35:21:@25820.4]
  wire [31:0] x339_io_out; // @[BigIPZynq.scala 35:21:@25820.4]
  wire [63:0] fix2fixBox_io_a; // @[Math.scala 357:30:@25827.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 357:30:@25827.4]
  Modulo x339 ( // @[BigIPZynq.scala 35:21:@25820.4]
    .clock(x339_clock),
    .io_flow(x339_io_flow),
    .io_dividend(x339_io_dividend),
    .io_divisor(x339_io_divisor),
    .io_out(x339_io_out)
  );
  fix2fixBox_38 fix2fixBox ( // @[Math.scala 357:30:@25827.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 363:17:@25835.4]
  assign x339_clock = clock; // @[:@25821.4]
  assign x339_io_flow = io_flow; // @[BigIPZynq.scala 38:17:@25825.4]
  assign x339_io_dividend = io_a; // @[BigIPZynq.scala 36:21:@25823.4]
  assign x339_io_divisor = 32'h6; // @[BigIPZynq.scala 37:20:@25824.4]
  assign fix2fixBox_io_a = {{32'd0}, x339_io_out}; // @[Math.scala 358:23:@25830.4]
endmodule
module Divider( // @[:@26029.2]
  input         clock, // @[:@26030.4]
  input         io_flow, // @[:@26032.4]
  input  [31:0] io_dividend, // @[:@26032.4]
  input  [31:0] io_divisor, // @[:@26032.4]
  output [31:0] io_out // @[:@26032.4]
);
  wire [31:0] m_m_axis_dout_tdata; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire  m_m_axis_dout_tvalid; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire [31:0] m_s_axis_divisor_tdata; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire  m_s_axis_divisor_tvalid; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire [31:0] m_s_axis_dividend_tdata; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire  m_s_axis_dividend_tvalid; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire  m_aclken; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire  m_aclk; // @[ZynqBlackBoxes.scala 26:19:@26034.4]
  wire [29:0] _T_15; // @[ZynqBlackBoxes.scala 34:37:@26050.4]
  div_32_32_20_Signed_Fractional m ( // @[ZynqBlackBoxes.scala 26:19:@26034.4]
    .m_axis_dout_tdata(m_m_axis_dout_tdata),
    .m_axis_dout_tvalid(m_m_axis_dout_tvalid),
    .s_axis_divisor_tdata(m_s_axis_divisor_tdata),
    .s_axis_divisor_tvalid(m_s_axis_divisor_tvalid),
    .s_axis_dividend_tdata(m_s_axis_dividend_tdata),
    .s_axis_dividend_tvalid(m_s_axis_dividend_tvalid),
    .aclken(m_aclken),
    .aclk(m_aclk)
  );
  assign _T_15 = m_m_axis_dout_tdata[31:2]; // @[ZynqBlackBoxes.scala 34:37:@26050.4]
  assign io_out = {{2'd0}, _T_15}; // @[ZynqBlackBoxes.scala 34:12:@26051.4]
  assign m_s_axis_divisor_tdata = io_divisor; // @[ZynqBlackBoxes.scala 32:31:@26048.4]
  assign m_s_axis_divisor_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 31:32:@26047.4]
  assign m_s_axis_dividend_tdata = io_dividend; // @[ZynqBlackBoxes.scala 30:32:@26046.4]
  assign m_s_axis_dividend_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 29:33:@26045.4]
  assign m_aclken = io_flow; // @[ZynqBlackBoxes.scala 28:17:@26044.4 ZynqBlackBoxes.scala 33:17:@26049.4]
  assign m_aclk = clock; // @[ZynqBlackBoxes.scala 27:15:@26043.4]
endmodule
module x342_div( // @[:@26089.2]
  input         clock, // @[:@26090.4]
  input  [31:0] io_a, // @[:@26092.4]
  input         io_flow, // @[:@26092.4]
  output [31:0] io_result // @[:@26092.4]
);
  wire  x342_div_clock; // @[BigIPZynq.scala 25:21:@26100.4]
  wire  x342_div_io_flow; // @[BigIPZynq.scala 25:21:@26100.4]
  wire [31:0] x342_div_io_dividend; // @[BigIPZynq.scala 25:21:@26100.4]
  wire [31:0] x342_div_io_divisor; // @[BigIPZynq.scala 25:21:@26100.4]
  wire [31:0] x342_div_io_out; // @[BigIPZynq.scala 25:21:@26100.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@26113.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@26113.4]
  wire [31:0] _T_15; // @[FixedPoint.scala 24:59:@26098.4]
  wire [31:0] _T_19; // @[BigIPZynq.scala 29:16:@26108.4]
  Divider x342_div ( // @[BigIPZynq.scala 25:21:@26100.4]
    .clock(x342_div_clock),
    .io_flow(x342_div_io_flow),
    .io_dividend(x342_div_io_dividend),
    .io_divisor(x342_div_io_divisor),
    .io_out(x342_div_io_out)
  );
  _ _ ( // @[Math.scala 720:24:@26113.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign _T_15 = $signed(io_a); // @[FixedPoint.scala 24:59:@26098.4]
  assign _T_19 = $signed(x342_div_io_out); // @[BigIPZynq.scala 29:16:@26108.4]
  assign io_result = __io_result; // @[Math.scala 290:34:@26121.4]
  assign x342_div_clock = clock; // @[:@26101.4]
  assign x342_div_io_flow = io_flow; // @[BigIPZynq.scala 28:17:@26107.4]
  assign x342_div_io_dividend = $unsigned(_T_15); // @[BigIPZynq.scala 26:21:@26104.4]
  assign x342_div_io_divisor = 32'h6; // @[BigIPZynq.scala 27:20:@26106.4]
  assign __io_b = $unsigned(_T_19); // @[Math.scala 721:17:@26116.4]
endmodule
module RetimeWrapper_298( // @[:@26135.2]
  input         clock, // @[:@26136.4]
  input         reset, // @[:@26137.4]
  input         io_flow, // @[:@26138.4]
  input  [31:0] io_in, // @[:@26138.4]
  output [31:0] io_out // @[:@26138.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26140.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26140.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26140.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26140.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26140.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26140.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(19)) sr ( // @[RetimeShiftRegister.scala 15:20:@26140.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26153.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26152.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26151.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26150.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26149.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26147.4]
endmodule
module RetimeWrapper_300( // @[:@26346.2]
  input         clock, // @[:@26347.4]
  input         reset, // @[:@26348.4]
  input         io_flow, // @[:@26349.4]
  input  [31:0] io_in, // @[:@26349.4]
  output [31:0] io_out // @[:@26349.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26351.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26351.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26351.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26351.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26351.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26351.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@26351.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26364.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26363.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26362.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26361.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26360.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26358.4]
endmodule
module RetimeWrapper_301( // @[:@26378.2]
  input         clock, // @[:@26379.4]
  input         reset, // @[:@26380.4]
  input         io_flow, // @[:@26381.4]
  input  [31:0] io_in, // @[:@26381.4]
  output [31:0] io_out // @[:@26381.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26383.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26383.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26383.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26383.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26383.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26383.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@26383.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26396.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26395.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26394.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26393.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26392.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26390.4]
endmodule
module RetimeWrapper_302( // @[:@26410.2]
  input         clock, // @[:@26411.4]
  input         reset, // @[:@26412.4]
  input         io_flow, // @[:@26413.4]
  input  [31:0] io_in, // @[:@26413.4]
  output [31:0] io_out // @[:@26413.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26415.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26415.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26415.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26415.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26415.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26415.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@26415.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26428.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26427.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26426.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26425.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26424.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26422.4]
endmodule
module RetimeWrapper_303( // @[:@26442.2]
  input   clock, // @[:@26443.4]
  input   reset, // @[:@26444.4]
  input   io_flow, // @[:@26445.4]
  input   io_in, // @[:@26445.4]
  output  io_out // @[:@26445.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@26447.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@26447.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@26447.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26447.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26447.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26447.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@26447.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26460.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26459.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@26458.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26457.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26456.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26454.4]
endmodule
module RetimeWrapper_305( // @[:@26506.2]
  input         clock, // @[:@26507.4]
  input         reset, // @[:@26508.4]
  input         io_flow, // @[:@26509.4]
  input  [31:0] io_in, // @[:@26509.4]
  output [31:0] io_out // @[:@26509.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26511.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26511.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26511.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26511.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26511.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26511.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@26511.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26524.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26523.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26522.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26521.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26520.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26518.4]
endmodule
module RetimeWrapper_308( // @[:@26938.2]
  input         clock, // @[:@26939.4]
  input         reset, // @[:@26940.4]
  input         io_flow, // @[:@26941.4]
  input  [31:0] io_in, // @[:@26941.4]
  output [31:0] io_out // @[:@26941.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26943.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26943.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26943.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26943.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26943.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26943.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@26943.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26956.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26955.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26954.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26953.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26952.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26950.4]
endmodule
module RetimeWrapper_310( // @[:@27149.2]
  input         clock, // @[:@27150.4]
  input         reset, // @[:@27151.4]
  input         io_flow, // @[:@27152.4]
  input  [31:0] io_in, // @[:@27152.4]
  output [31:0] io_out // @[:@27152.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@27154.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@27154.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@27154.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@27154.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@27154.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@27154.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@27154.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@27167.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@27166.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@27165.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@27164.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@27163.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@27161.4]
endmodule
module RetimeWrapper_311( // @[:@27181.2]
  input         clock, // @[:@27182.4]
  input         reset, // @[:@27183.4]
  input         io_flow, // @[:@27184.4]
  input  [31:0] io_in, // @[:@27184.4]
  output [31:0] io_out // @[:@27184.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@27186.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@27186.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@27186.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@27186.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@27186.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@27186.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@27186.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@27199.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@27198.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@27197.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@27196.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@27195.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@27193.4]
endmodule
module RetimeWrapper_326( // @[:@28627.2]
  input         clock, // @[:@28628.4]
  input         reset, // @[:@28629.4]
  input         io_flow, // @[:@28630.4]
  input  [31:0] io_in, // @[:@28630.4]
  output [31:0] io_out // @[:@28630.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@28632.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@28632.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@28632.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@28632.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@28632.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@28632.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(26)) sr ( // @[RetimeShiftRegister.scala 15:20:@28632.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@28645.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@28644.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@28643.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@28642.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@28641.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@28639.4]
endmodule
module RetimeWrapper_332( // @[:@28819.2]
  input         clock, // @[:@28820.4]
  input         reset, // @[:@28821.4]
  input         io_flow, // @[:@28822.4]
  input  [31:0] io_in, // @[:@28822.4]
  output [31:0] io_out // @[:@28822.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@28824.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@28824.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@28824.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@28824.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@28824.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@28824.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(48)) sr ( // @[RetimeShiftRegister.scala 15:20:@28824.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@28837.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@28836.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@28835.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@28834.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@28833.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@28831.4]
endmodule
module RetimeWrapper_333( // @[:@28851.2]
  input   clock, // @[:@28852.4]
  input   reset, // @[:@28853.4]
  input   io_flow, // @[:@28854.4]
  input   io_in, // @[:@28854.4]
  output  io_out // @[:@28854.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@28856.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@28856.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@28856.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@28856.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@28856.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@28856.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@28856.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@28869.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@28868.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@28867.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@28866.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@28865.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@28863.4]
endmodule
module RetimeWrapper_334( // @[:@28883.2]
  input   clock, // @[:@28884.4]
  input   reset, // @[:@28885.4]
  input   io_flow, // @[:@28886.4]
  input   io_in, // @[:@28886.4]
  output  io_out // @[:@28886.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@28888.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@28888.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@28888.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@28888.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@28888.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@28888.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(48)) sr ( // @[RetimeShiftRegister.scala 15:20:@28888.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@28901.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@28900.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@28899.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@28898.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@28897.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@28895.4]
endmodule
module RetimeWrapper_336( // @[:@28947.2]
  input         clock, // @[:@28948.4]
  input         reset, // @[:@28949.4]
  input         io_flow, // @[:@28950.4]
  input  [31:0] io_in, // @[:@28950.4]
  output [31:0] io_out // @[:@28950.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@28952.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@28952.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@28952.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@28952.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@28952.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@28952.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(31)) sr ( // @[RetimeShiftRegister.scala 15:20:@28952.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@28965.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@28964.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@28963.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@28962.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@28961.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@28959.4]
endmodule
module RetimeWrapper_352( // @[:@29459.2]
  input         clock, // @[:@29460.4]
  input         reset, // @[:@29461.4]
  input         io_flow, // @[:@29462.4]
  input  [31:0] io_in, // @[:@29462.4]
  output [31:0] io_out // @[:@29462.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@29464.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@29464.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@29464.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29464.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29464.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29464.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(32)) sr ( // @[RetimeShiftRegister.scala 15:20:@29464.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29477.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29476.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@29475.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29474.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29473.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29471.4]
endmodule
module RetimeWrapper_353( // @[:@29491.2]
  input         clock, // @[:@29492.4]
  input         reset, // @[:@29493.4]
  input         io_flow, // @[:@29494.4]
  input  [31:0] io_in, // @[:@29494.4]
  output [31:0] io_out // @[:@29494.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@29496.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@29496.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@29496.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29496.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29496.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29496.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(27)) sr ( // @[RetimeShiftRegister.scala 15:20:@29496.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29509.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29508.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@29507.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29506.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29505.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29503.4]
endmodule
module RetimeWrapper_354( // @[:@29523.2]
  input   clock, // @[:@29524.4]
  input   reset, // @[:@29525.4]
  input   io_flow, // @[:@29526.4]
  input   io_in, // @[:@29526.4]
  output  io_out // @[:@29526.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@29528.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@29528.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@29528.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29528.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29528.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29528.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@29528.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29541.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29540.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@29539.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29538.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29537.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29535.4]
endmodule
module RetimeWrapper_358( // @[:@29987.2]
  input         clock, // @[:@29988.4]
  input         reset, // @[:@29989.4]
  input         io_flow, // @[:@29990.4]
  input  [31:0] io_in, // @[:@29990.4]
  output [31:0] io_out // @[:@29990.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@29992.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@29992.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@29992.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29992.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29992.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29992.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(46)) sr ( // @[RetimeShiftRegister.scala 15:20:@29992.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30005.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30004.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30003.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30002.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30001.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29999.4]
endmodule
module RetimeWrapper_360( // @[:@30198.2]
  input         clock, // @[:@30199.4]
  input         reset, // @[:@30200.4]
  input         io_flow, // @[:@30201.4]
  input  [31:0] io_in, // @[:@30201.4]
  output [31:0] io_out // @[:@30201.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30203.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30203.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30203.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30203.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30203.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30203.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@30203.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30216.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30215.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30214.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30213.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30212.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30210.4]
endmodule
module RetimeWrapper_374( // @[:@31424.2]
  input         clock, // @[:@31425.4]
  input         reset, // @[:@31426.4]
  input         io_flow, // @[:@31427.4]
  input  [31:0] io_in, // @[:@31427.4]
  output [31:0] io_out // @[:@31427.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31429.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31429.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31429.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31429.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31429.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31429.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@31429.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31442.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31441.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31440.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31439.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31438.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31436.4]
endmodule
module RetimeWrapper_390( // @[:@32377.2]
  input         clock, // @[:@32378.4]
  input         reset, // @[:@32379.4]
  input         io_flow, // @[:@32380.4]
  input  [31:0] io_in, // @[:@32380.4]
  output [31:0] io_out // @[:@32380.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@32382.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@32382.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@32382.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@32382.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@32382.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@32382.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(17)) sr ( // @[RetimeShiftRegister.scala 15:20:@32382.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@32395.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@32394.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@32393.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@32392.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@32391.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@32389.4]
endmodule
module Multiplier( // @[:@35209.2]
  input         clock, // @[:@35210.4]
  input         io_flow, // @[:@35212.4]
  input  [31:0] io_a, // @[:@35212.4]
  input  [31:0] io_b, // @[:@35212.4]
  output [31:0] io_out // @[:@35212.4]
);
  wire [31:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@35214.4]
  wire [31:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@35214.4]
  wire [31:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@35214.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@35214.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@35214.4]
  mul_32_32_32_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@35214.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@35224.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@35222.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@35221.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@35223.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@35220.4]
endmodule
module x475( // @[:@35244.2]
  input         clock, // @[:@35245.4]
  input  [31:0] io_a, // @[:@35247.4]
  input  [31:0] io_b, // @[:@35247.4]
  input         io_flow, // @[:@35247.4]
  output [31:0] io_result // @[:@35247.4]
);
  wire  x475_clock; // @[BigIPZynq.scala 63:21:@35254.4]
  wire  x475_io_flow; // @[BigIPZynq.scala 63:21:@35254.4]
  wire [31:0] x475_io_a; // @[BigIPZynq.scala 63:21:@35254.4]
  wire [31:0] x475_io_b; // @[BigIPZynq.scala 63:21:@35254.4]
  wire [31:0] x475_io_out; // @[BigIPZynq.scala 63:21:@35254.4]
  wire [31:0] fix2fixBox_io_a; // @[Math.scala 253:30:@35263.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@35263.4]
  Multiplier x475 ( // @[BigIPZynq.scala 63:21:@35254.4]
    .clock(x475_clock),
    .io_flow(x475_io_flow),
    .io_a(x475_io_a),
    .io_b(x475_io_b),
    .io_out(x475_io_out)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 253:30:@35263.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@35271.4]
  assign x475_clock = clock; // @[:@35255.4]
  assign x475_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@35259.4]
  assign x475_io_a = io_a; // @[BigIPZynq.scala 64:14:@35257.4]
  assign x475_io_b = io_b; // @[BigIPZynq.scala 65:14:@35258.4]
  assign fix2fixBox_io_a = x475_io_out; // @[Math.scala 254:23:@35266.4]
endmodule
module fix2fixBox_143( // @[:@35865.2]
  input  [31:0] io_a, // @[:@35868.4]
  output [32:0] io_b // @[:@35868.4]
);
  assign io_b = {1'h0,io_a}; // @[Converter.scala 95:38:@35882.4]
endmodule
module __86( // @[:@35884.2]
  input  [31:0] io_b, // @[:@35887.4]
  output [32:0] io_result // @[:@35887.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@35892.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@35892.4]
  fix2fixBox_143 fix2fixBox ( // @[BigIPZynq.scala 219:30:@35892.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@35900.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@35895.4]
endmodule
module x484_x3( // @[:@35996.2]
  input         clock, // @[:@35997.4]
  input         reset, // @[:@35998.4]
  input  [31:0] io_a, // @[:@35999.4]
  input  [31:0] io_b, // @[:@35999.4]
  input         io_flow, // @[:@35999.4]
  output [31:0] io_result // @[:@35999.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@36007.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@36007.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@36014.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@36014.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@36024.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@36024.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@36024.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@36024.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@36024.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@36012.4 Math.scala 724:14:@36013.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@36019.4 Math.scala 724:14:@36020.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@36021.4]
  __86 _ ( // @[Math.scala 720:24:@36007.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __86 __1 ( // @[Math.scala 720:24:@36014.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@36024.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@36012.4 Math.scala 724:14:@36013.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@36019.4 Math.scala 724:14:@36020.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@36021.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@36032.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@36010.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@36017.4]
  assign fix2fixBox_clock = clock; // @[:@36025.4]
  assign fix2fixBox_reset = reset; // @[:@36026.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@36027.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@36030.4]
endmodule
module fix2fixBox_167( // @[:@37249.2]
  input  [31:0] io_a, // @[:@37252.4]
  output [31:0] io_b // @[:@37252.4]
);
  wire [24:0] new_dec; // @[Converter.scala 63:26:@37262.4]
  assign new_dec = io_a[24:0]; // @[Converter.scala 63:26:@37262.4]
  assign io_b = {new_dec,7'h0}; // @[Converter.scala 94:38:@37265.4]
endmodule
module x492( // @[:@37267.2]
  input  [31:0] io_b, // @[:@37270.4]
  output [31:0] io_result // @[:@37270.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@37275.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@37275.4]
  fix2fixBox_167 fix2fixBox ( // @[BigIPZynq.scala 219:30:@37275.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@37283.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@37278.4]
endmodule
module Multiplier_9( // @[:@37295.2]
  input         clock, // @[:@37296.4]
  input         io_flow, // @[:@37298.4]
  input  [38:0] io_a, // @[:@37298.4]
  input  [38:0] io_b, // @[:@37298.4]
  output [38:0] io_out // @[:@37298.4]
);
  wire [38:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@37300.4]
  wire [38:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@37300.4]
  wire [38:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@37300.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@37300.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@37300.4]
  mul_39_39_39_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@37300.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@37310.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@37308.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@37307.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@37309.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@37306.4]
endmodule
module fix2fixBox_168( // @[:@37312.2]
  input  [38:0] io_a, // @[:@37315.4]
  output [31:0] io_b // @[:@37315.4]
);
  wire [6:0] tmp_frac; // @[Converter.scala 38:42:@37323.4]
  wire [24:0] new_dec; // @[Converter.scala 88:34:@37326.4]
  assign tmp_frac = io_a[13:7]; // @[Converter.scala 38:42:@37323.4]
  assign new_dec = io_a[38:14]; // @[Converter.scala 88:34:@37326.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@37329.4]
endmodule
module x493_mul( // @[:@37331.2]
  input         clock, // @[:@37332.4]
  input  [31:0] io_a, // @[:@37334.4]
  input         io_flow, // @[:@37334.4]
  output [31:0] io_result // @[:@37334.4]
);
  wire  x493_mul_clock; // @[BigIPZynq.scala 63:21:@37349.4]
  wire  x493_mul_io_flow; // @[BigIPZynq.scala 63:21:@37349.4]
  wire [38:0] x493_mul_io_a; // @[BigIPZynq.scala 63:21:@37349.4]
  wire [38:0] x493_mul_io_b; // @[BigIPZynq.scala 63:21:@37349.4]
  wire [38:0] x493_mul_io_out; // @[BigIPZynq.scala 63:21:@37349.4]
  wire [38:0] fix2fixBox_io_a; // @[Math.scala 253:30:@37357.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@37357.4]
  wire  _T_16; // @[FixedPoint.scala 50:25:@37341.4]
  wire [6:0] _T_20; // @[Bitwise.scala 72:12:@37343.4]
  Multiplier_9 x493_mul ( // @[BigIPZynq.scala 63:21:@37349.4]
    .clock(x493_mul_clock),
    .io_flow(x493_mul_io_flow),
    .io_a(x493_mul_io_a),
    .io_b(x493_mul_io_b),
    .io_out(x493_mul_io_out)
  );
  fix2fixBox_168 fix2fixBox ( // @[Math.scala 253:30:@37357.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_16 = io_a[31]; // @[FixedPoint.scala 50:25:@37341.4]
  assign _T_20 = _T_16 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@37343.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@37365.4]
  assign x493_mul_clock = clock; // @[:@37350.4]
  assign x493_mul_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@37354.4]
  assign x493_mul_io_a = {_T_20,io_a}; // @[BigIPZynq.scala 64:14:@37352.4]
  assign x493_mul_io_b = 39'h8; // @[BigIPZynq.scala 65:14:@37353.4]
  assign fix2fixBox_io_a = x493_mul_io_out; // @[Math.scala 254:23:@37360.4]
endmodule
module fix2fixBox_169( // @[:@37367.2]
  input  [31:0] io_a, // @[:@37370.4]
  output [31:0] io_b // @[:@37370.4]
);
  wire [24:0] _T_25; // @[Converter.scala 84:75:@37382.4]
  assign _T_25 = io_a[31:7]; // @[Converter.scala 84:75:@37382.4]
  assign io_b = {7'h0,_T_25}; // @[Converter.scala 95:38:@37385.4]
endmodule
module x494( // @[:@37387.2]
  input  [31:0] io_b, // @[:@37390.4]
  output [31:0] io_result // @[:@37390.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@37395.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@37395.4]
  fix2fixBox_169 fix2fixBox ( // @[BigIPZynq.scala 219:30:@37395.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@37403.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@37398.4]
endmodule
module RetimeWrapper_464( // @[:@43591.2]
  input          clock, // @[:@43592.4]
  input          reset, // @[:@43593.4]
  input          io_flow, // @[:@43594.4]
  input  [127:0] io_in, // @[:@43594.4]
  output [127:0] io_out // @[:@43594.4]
);
  wire [127:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@43596.4]
  wire [127:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@43596.4]
  wire [127:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@43596.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@43596.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@43596.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@43596.4]
  RetimeShiftRegister #(.WIDTH(128), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@43596.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@43609.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@43608.4]
  assign sr_init = 128'h0; // @[RetimeShiftRegister.scala 19:16:@43607.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@43606.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@43605.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@43603.4]
endmodule
module x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@43707.2]
  input          clock, // @[:@43708.4]
  input          reset, // @[:@43709.4]
  output         io_in_x289_TREADY, // @[:@43710.4]
  input  [255:0] io_in_x289_TDATA, // @[:@43710.4]
  input  [7:0]   io_in_x289_TID, // @[:@43710.4]
  input  [7:0]   io_in_x289_TDEST, // @[:@43710.4]
  output         io_in_x290_TVALID, // @[:@43710.4]
  input          io_in_x290_TREADY, // @[:@43710.4]
  output [255:0] io_in_x290_TDATA, // @[:@43710.4]
  input          io_sigsIn_backpressure, // @[:@43710.4]
  input          io_sigsIn_datapathEn, // @[:@43710.4]
  input          io_sigsIn_break, // @[:@43710.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@43710.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@43710.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@43710.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@43710.4]
  input          io_rr // @[:@43710.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@43724.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@43724.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@43736.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@43736.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@43759.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@43759.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@43759.4]
  wire [127:0] RetimeWrapper_io_in; // @[package.scala 93:22:@43759.4]
  wire [127:0] RetimeWrapper_io_out; // @[package.scala 93:22:@43759.4]
  wire  x334_lb_0_clock; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_reset; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_17_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_17_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_17_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_17_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_17_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_17_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_16_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_16_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_16_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_16_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_16_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_16_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_15_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_15_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_15_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_15_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_15_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_15_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_14_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_14_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_14_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_14_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_14_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_14_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_13_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_13_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_13_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_13_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_13_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_13_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_12_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_12_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_12_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_12_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_12_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_12_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_11_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_11_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_11_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_11_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_11_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_11_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_10_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_10_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_10_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_10_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_10_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_10_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_9_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_9_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_9_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_9_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_9_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_9_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_8_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_8_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_8_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_8_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_8_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_8_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_7_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_7_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_7_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_7_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_7_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_7_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_6_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_6_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_6_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_6_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_6_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_6_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_5_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_5_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_5_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_5_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_5_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_5_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_4_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_4_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_4_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_4_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_4_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_4_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_3_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_3_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_3_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_3_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_3_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_3_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_2_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_2_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_2_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_2_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_2_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_2_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_1_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_1_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_1_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_1_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_1_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_1_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_0_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_rPort_0_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_rPort_0_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_0_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_rPort_0_backpressure; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_rPort_0_output_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_wPort_3_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_wPort_3_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_wPort_3_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_wPort_3_data_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_wPort_3_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_wPort_2_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_wPort_2_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_wPort_2_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_wPort_2_data_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_wPort_2_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_wPort_1_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_wPort_1_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_wPort_1_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_wPort_1_data_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_wPort_1_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_wPort_0_banks_1; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [2:0] x334_lb_0_io_wPort_0_banks_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [8:0] x334_lb_0_io_wPort_0_ofs_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire [31:0] x334_lb_0_io_wPort_0_data_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x334_lb_0_io_wPort_0_en_0; // @[m_x334_lb_0.scala 47:17:@43769.4]
  wire  x339_1_clock; // @[Math.scala 366:24:@43952.4]
  wire [31:0] x339_1_io_a; // @[Math.scala 366:24:@43952.4]
  wire  x339_1_io_flow; // @[Math.scala 366:24:@43952.4]
  wire [31:0] x339_1_io_result; // @[Math.scala 366:24:@43952.4]
  wire  x621_sum_1_clock; // @[Math.scala 150:24:@43989.4]
  wire  x621_sum_1_reset; // @[Math.scala 150:24:@43989.4]
  wire [31:0] x621_sum_1_io_a; // @[Math.scala 150:24:@43989.4]
  wire [31:0] x621_sum_1_io_b; // @[Math.scala 150:24:@43989.4]
  wire  x621_sum_1_io_flow; // @[Math.scala 150:24:@43989.4]
  wire [31:0] x621_sum_1_io_result; // @[Math.scala 150:24:@43989.4]
  wire  x342_div_1_clock; // @[Math.scala 327:24:@44001.4]
  wire [31:0] x342_div_1_io_a; // @[Math.scala 327:24:@44001.4]
  wire  x342_div_1_io_flow; // @[Math.scala 327:24:@44001.4]
  wire [31:0] x342_div_1_io_result; // @[Math.scala 327:24:@44001.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@44011.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@44011.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@44011.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@44011.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@44011.4]
  wire  x343_sum_1_clock; // @[Math.scala 150:24:@44020.4]
  wire  x343_sum_1_reset; // @[Math.scala 150:24:@44020.4]
  wire [31:0] x343_sum_1_io_a; // @[Math.scala 150:24:@44020.4]
  wire [31:0] x343_sum_1_io_b; // @[Math.scala 150:24:@44020.4]
  wire  x343_sum_1_io_flow; // @[Math.scala 150:24:@44020.4]
  wire [31:0] x343_sum_1_io_result; // @[Math.scala 150:24:@44020.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@44030.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@44030.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@44030.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@44030.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@44030.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@44039.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@44039.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@44039.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@44039.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@44039.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@44048.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@44048.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@44048.4]
  wire [31:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@44048.4]
  wire [31:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@44048.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@44057.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@44057.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@44057.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@44057.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@44057.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@44066.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@44066.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@44066.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@44066.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@44066.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@44075.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@44075.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@44075.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@44075.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@44075.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@44086.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@44086.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@44086.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@44086.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@44086.4]
  wire  x345_rdcol_1_clock; // @[Math.scala 150:24:@44109.4]
  wire  x345_rdcol_1_reset; // @[Math.scala 150:24:@44109.4]
  wire [31:0] x345_rdcol_1_io_a; // @[Math.scala 150:24:@44109.4]
  wire [31:0] x345_rdcol_1_io_b; // @[Math.scala 150:24:@44109.4]
  wire  x345_rdcol_1_io_flow; // @[Math.scala 150:24:@44109.4]
  wire [31:0] x345_rdcol_1_io_result; // @[Math.scala 150:24:@44109.4]
  wire  x347_1_clock; // @[Math.scala 366:24:@44123.4]
  wire [31:0] x347_1_io_a; // @[Math.scala 366:24:@44123.4]
  wire  x347_1_io_flow; // @[Math.scala 366:24:@44123.4]
  wire [31:0] x347_1_io_result; // @[Math.scala 366:24:@44123.4]
  wire  x348_div_1_clock; // @[Math.scala 327:24:@44135.4]
  wire [31:0] x348_div_1_io_a; // @[Math.scala 327:24:@44135.4]
  wire  x348_div_1_io_flow; // @[Math.scala 327:24:@44135.4]
  wire [31:0] x348_div_1_io_result; // @[Math.scala 327:24:@44135.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@44145.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@44145.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@44145.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@44145.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@44145.4]
  wire  x349_sum_1_clock; // @[Math.scala 150:24:@44154.4]
  wire  x349_sum_1_reset; // @[Math.scala 150:24:@44154.4]
  wire [31:0] x349_sum_1_io_a; // @[Math.scala 150:24:@44154.4]
  wire [31:0] x349_sum_1_io_b; // @[Math.scala 150:24:@44154.4]
  wire  x349_sum_1_io_flow; // @[Math.scala 150:24:@44154.4]
  wire [31:0] x349_sum_1_io_result; // @[Math.scala 150:24:@44154.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@44164.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@44164.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@44164.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@44164.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@44164.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@44173.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@44173.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@44173.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@44173.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@44173.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@44182.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@44182.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@44182.4]
  wire [31:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@44182.4]
  wire [31:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@44182.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@44193.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@44193.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@44193.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@44193.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@44193.4]
  wire  x351_rdcol_1_clock; // @[Math.scala 150:24:@44216.4]
  wire  x351_rdcol_1_reset; // @[Math.scala 150:24:@44216.4]
  wire [31:0] x351_rdcol_1_io_a; // @[Math.scala 150:24:@44216.4]
  wire [31:0] x351_rdcol_1_io_b; // @[Math.scala 150:24:@44216.4]
  wire  x351_rdcol_1_io_flow; // @[Math.scala 150:24:@44216.4]
  wire [31:0] x351_rdcol_1_io_result; // @[Math.scala 150:24:@44216.4]
  wire  x353_1_clock; // @[Math.scala 366:24:@44230.4]
  wire [31:0] x353_1_io_a; // @[Math.scala 366:24:@44230.4]
  wire  x353_1_io_flow; // @[Math.scala 366:24:@44230.4]
  wire [31:0] x353_1_io_result; // @[Math.scala 366:24:@44230.4]
  wire  x354_div_1_clock; // @[Math.scala 327:24:@44242.4]
  wire [31:0] x354_div_1_io_a; // @[Math.scala 327:24:@44242.4]
  wire  x354_div_1_io_flow; // @[Math.scala 327:24:@44242.4]
  wire [31:0] x354_div_1_io_result; // @[Math.scala 327:24:@44242.4]
  wire  x355_sum_1_clock; // @[Math.scala 150:24:@44252.4]
  wire  x355_sum_1_reset; // @[Math.scala 150:24:@44252.4]
  wire [31:0] x355_sum_1_io_a; // @[Math.scala 150:24:@44252.4]
  wire [31:0] x355_sum_1_io_b; // @[Math.scala 150:24:@44252.4]
  wire  x355_sum_1_io_flow; // @[Math.scala 150:24:@44252.4]
  wire [31:0] x355_sum_1_io_result; // @[Math.scala 150:24:@44252.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@44262.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@44262.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@44262.4]
  wire [31:0] RetimeWrapper_14_io_in; // @[package.scala 93:22:@44262.4]
  wire [31:0] RetimeWrapper_14_io_out; // @[package.scala 93:22:@44262.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@44271.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@44271.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@44271.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@44271.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@44271.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@44280.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@44280.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@44280.4]
  wire [31:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@44280.4]
  wire [31:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@44280.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@44291.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@44291.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@44291.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@44291.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@44291.4]
  wire  x357_rdcol_1_clock; // @[Math.scala 150:24:@44314.4]
  wire  x357_rdcol_1_reset; // @[Math.scala 150:24:@44314.4]
  wire [31:0] x357_rdcol_1_io_a; // @[Math.scala 150:24:@44314.4]
  wire [31:0] x357_rdcol_1_io_b; // @[Math.scala 150:24:@44314.4]
  wire  x357_rdcol_1_io_flow; // @[Math.scala 150:24:@44314.4]
  wire [31:0] x357_rdcol_1_io_result; // @[Math.scala 150:24:@44314.4]
  wire  x359_1_clock; // @[Math.scala 366:24:@44328.4]
  wire [31:0] x359_1_io_a; // @[Math.scala 366:24:@44328.4]
  wire  x359_1_io_flow; // @[Math.scala 366:24:@44328.4]
  wire [31:0] x359_1_io_result; // @[Math.scala 366:24:@44328.4]
  wire  x360_div_1_clock; // @[Math.scala 327:24:@44340.4]
  wire [31:0] x360_div_1_io_a; // @[Math.scala 327:24:@44340.4]
  wire  x360_div_1_io_flow; // @[Math.scala 327:24:@44340.4]
  wire [31:0] x360_div_1_io_result; // @[Math.scala 327:24:@44340.4]
  wire  x361_sum_1_clock; // @[Math.scala 150:24:@44350.4]
  wire  x361_sum_1_reset; // @[Math.scala 150:24:@44350.4]
  wire [31:0] x361_sum_1_io_a; // @[Math.scala 150:24:@44350.4]
  wire [31:0] x361_sum_1_io_b; // @[Math.scala 150:24:@44350.4]
  wire  x361_sum_1_io_flow; // @[Math.scala 150:24:@44350.4]
  wire [31:0] x361_sum_1_io_result; // @[Math.scala 150:24:@44350.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@44360.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@44360.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@44360.4]
  wire [31:0] RetimeWrapper_18_io_in; // @[package.scala 93:22:@44360.4]
  wire [31:0] RetimeWrapper_18_io_out; // @[package.scala 93:22:@44360.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@44369.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@44369.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@44369.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@44369.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@44369.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@44378.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@44378.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@44378.4]
  wire [31:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@44378.4]
  wire [31:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@44378.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@44389.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@44389.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@44389.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@44389.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@44389.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@44410.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@44410.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@44410.4]
  wire [31:0] RetimeWrapper_22_io_in; // @[package.scala 93:22:@44410.4]
  wire [31:0] RetimeWrapper_22_io_out; // @[package.scala 93:22:@44410.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@44426.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@44426.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@44426.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@44426.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@44426.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@44435.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@44435.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@44435.4]
  wire [31:0] RetimeWrapper_24_io_in; // @[package.scala 93:22:@44435.4]
  wire [31:0] RetimeWrapper_24_io_out; // @[package.scala 93:22:@44435.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@44449.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@44449.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@44449.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@44449.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@44449.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@44458.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@44458.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@44458.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@44458.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@44458.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@44473.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@44473.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@44473.4]
  wire [31:0] RetimeWrapper_27_io_in; // @[package.scala 93:22:@44473.4]
  wire [31:0] RetimeWrapper_27_io_out; // @[package.scala 93:22:@44473.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@44482.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@44482.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@44482.4]
  wire [31:0] RetimeWrapper_28_io_in; // @[package.scala 93:22:@44482.4]
  wire [31:0] RetimeWrapper_28_io_out; // @[package.scala 93:22:@44482.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@44491.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@44491.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@44491.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@44491.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@44491.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@44500.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@44500.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@44500.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@44500.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@44500.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@44509.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@44509.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@44509.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@44509.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@44509.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@44518.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@44518.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@44518.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@44518.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@44518.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@44530.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@44530.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@44530.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@44530.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@44530.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@44551.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@44551.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@44551.4]
  wire [31:0] RetimeWrapper_34_io_in; // @[package.scala 93:22:@44551.4]
  wire [31:0] RetimeWrapper_34_io_out; // @[package.scala 93:22:@44551.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@44565.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@44565.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@44565.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@44565.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@44565.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@44580.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@44580.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@44580.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@44580.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@44580.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@44589.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@44589.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@44589.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@44589.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@44589.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@44598.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@44598.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@44598.4]
  wire [31:0] RetimeWrapper_38_io_in; // @[package.scala 93:22:@44598.4]
  wire [31:0] RetimeWrapper_38_io_out; // @[package.scala 93:22:@44598.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@44610.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@44610.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@44610.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@44610.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@44610.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@44631.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@44631.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@44631.4]
  wire [31:0] RetimeWrapper_40_io_in; // @[package.scala 93:22:@44631.4]
  wire [31:0] RetimeWrapper_40_io_out; // @[package.scala 93:22:@44631.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@44645.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@44645.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@44645.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@44645.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@44645.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@44660.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@44660.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@44660.4]
  wire [31:0] RetimeWrapper_42_io_in; // @[package.scala 93:22:@44660.4]
  wire [31:0] RetimeWrapper_42_io_out; // @[package.scala 93:22:@44660.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@44669.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@44669.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@44669.4]
  wire [31:0] RetimeWrapper_43_io_in; // @[package.scala 93:22:@44669.4]
  wire [31:0] RetimeWrapper_43_io_out; // @[package.scala 93:22:@44669.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@44678.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@44678.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@44678.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@44678.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@44678.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@44690.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@44690.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@44690.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@44690.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@44690.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@44711.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@44711.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@44711.4]
  wire [31:0] RetimeWrapper_46_io_in; // @[package.scala 93:22:@44711.4]
  wire [31:0] RetimeWrapper_46_io_out; // @[package.scala 93:22:@44711.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@44725.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@44725.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@44725.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@44725.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@44725.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@44740.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@44740.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@44740.4]
  wire [31:0] RetimeWrapper_48_io_in; // @[package.scala 93:22:@44740.4]
  wire [31:0] RetimeWrapper_48_io_out; // @[package.scala 93:22:@44740.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@44749.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@44749.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@44749.4]
  wire [31:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@44749.4]
  wire [31:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@44749.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@44758.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@44758.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@44758.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@44758.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@44758.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@44770.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@44770.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@44770.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@44770.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@44770.4]
  wire  x385_rdcol_1_clock; // @[Math.scala 150:24:@44793.4]
  wire  x385_rdcol_1_reset; // @[Math.scala 150:24:@44793.4]
  wire [31:0] x385_rdcol_1_io_a; // @[Math.scala 150:24:@44793.4]
  wire [31:0] x385_rdcol_1_io_b; // @[Math.scala 150:24:@44793.4]
  wire  x385_rdcol_1_io_flow; // @[Math.scala 150:24:@44793.4]
  wire [31:0] x385_rdcol_1_io_result; // @[Math.scala 150:24:@44793.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@44808.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@44808.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@44808.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@44808.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@44808.4]
  wire  x389_1_clock; // @[Math.scala 366:24:@44827.4]
  wire [31:0] x389_1_io_a; // @[Math.scala 366:24:@44827.4]
  wire  x389_1_io_flow; // @[Math.scala 366:24:@44827.4]
  wire [31:0] x389_1_io_result; // @[Math.scala 366:24:@44827.4]
  wire  x390_div_1_clock; // @[Math.scala 327:24:@44839.4]
  wire [31:0] x390_div_1_io_a; // @[Math.scala 327:24:@44839.4]
  wire  x390_div_1_io_flow; // @[Math.scala 327:24:@44839.4]
  wire [31:0] x390_div_1_io_result; // @[Math.scala 327:24:@44839.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@44849.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@44849.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@44849.4]
  wire [31:0] RetimeWrapper_53_io_in; // @[package.scala 93:22:@44849.4]
  wire [31:0] RetimeWrapper_53_io_out; // @[package.scala 93:22:@44849.4]
  wire  x391_sum_1_clock; // @[Math.scala 150:24:@44858.4]
  wire  x391_sum_1_reset; // @[Math.scala 150:24:@44858.4]
  wire [31:0] x391_sum_1_io_a; // @[Math.scala 150:24:@44858.4]
  wire [31:0] x391_sum_1_io_b; // @[Math.scala 150:24:@44858.4]
  wire  x391_sum_1_io_flow; // @[Math.scala 150:24:@44858.4]
  wire [31:0] x391_sum_1_io_result; // @[Math.scala 150:24:@44858.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@44868.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@44868.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@44868.4]
  wire [31:0] RetimeWrapper_54_io_in; // @[package.scala 93:22:@44868.4]
  wire [31:0] RetimeWrapper_54_io_out; // @[package.scala 93:22:@44868.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@44877.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@44877.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@44877.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@44877.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@44877.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@44889.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@44889.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@44889.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@44889.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@44889.4]
  wire  x394_rdcol_1_clock; // @[Math.scala 150:24:@44912.4]
  wire  x394_rdcol_1_reset; // @[Math.scala 150:24:@44912.4]
  wire [31:0] x394_rdcol_1_io_a; // @[Math.scala 150:24:@44912.4]
  wire [31:0] x394_rdcol_1_io_b; // @[Math.scala 150:24:@44912.4]
  wire  x394_rdcol_1_io_flow; // @[Math.scala 150:24:@44912.4]
  wire [31:0] x394_rdcol_1_io_result; // @[Math.scala 150:24:@44912.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@44927.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@44927.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@44927.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@44927.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@44927.4]
  wire  x398_1_clock; // @[Math.scala 366:24:@44944.4]
  wire [31:0] x398_1_io_a; // @[Math.scala 366:24:@44944.4]
  wire  x398_1_io_flow; // @[Math.scala 366:24:@44944.4]
  wire [31:0] x398_1_io_result; // @[Math.scala 366:24:@44944.4]
  wire  x399_div_1_clock; // @[Math.scala 327:24:@44956.4]
  wire [31:0] x399_div_1_io_a; // @[Math.scala 327:24:@44956.4]
  wire  x399_div_1_io_flow; // @[Math.scala 327:24:@44956.4]
  wire [31:0] x399_div_1_io_result; // @[Math.scala 327:24:@44956.4]
  wire  x400_sum_1_clock; // @[Math.scala 150:24:@44966.4]
  wire  x400_sum_1_reset; // @[Math.scala 150:24:@44966.4]
  wire [31:0] x400_sum_1_io_a; // @[Math.scala 150:24:@44966.4]
  wire [31:0] x400_sum_1_io_b; // @[Math.scala 150:24:@44966.4]
  wire  x400_sum_1_io_flow; // @[Math.scala 150:24:@44966.4]
  wire [31:0] x400_sum_1_io_result; // @[Math.scala 150:24:@44966.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@44976.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@44976.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@44976.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@44976.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@44976.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@44985.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@44985.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@44985.4]
  wire [31:0] RetimeWrapper_59_io_in; // @[package.scala 93:22:@44985.4]
  wire [31:0] RetimeWrapper_59_io_out; // @[package.scala 93:22:@44985.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@44997.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@44997.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@44997.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@44997.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@44997.4]
  wire  x403_rdrow_1_clock; // @[Math.scala 191:24:@45020.4]
  wire  x403_rdrow_1_reset; // @[Math.scala 191:24:@45020.4]
  wire [31:0] x403_rdrow_1_io_a; // @[Math.scala 191:24:@45020.4]
  wire [31:0] x403_rdrow_1_io_b; // @[Math.scala 191:24:@45020.4]
  wire  x403_rdrow_1_io_flow; // @[Math.scala 191:24:@45020.4]
  wire [31:0] x403_rdrow_1_io_result; // @[Math.scala 191:24:@45020.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@45046.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@45046.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@45046.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@45046.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@45046.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@45068.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@45068.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@45068.4]
  wire [31:0] RetimeWrapper_62_io_in; // @[package.scala 93:22:@45068.4]
  wire [31:0] RetimeWrapper_62_io_out; // @[package.scala 93:22:@45068.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@45094.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@45094.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@45094.4]
  wire [31:0] RetimeWrapper_63_io_in; // @[package.scala 93:22:@45094.4]
  wire [31:0] RetimeWrapper_63_io_out; // @[package.scala 93:22:@45094.4]
  wire  x626_sum_1_clock; // @[Math.scala 150:24:@45115.4]
  wire  x626_sum_1_reset; // @[Math.scala 150:24:@45115.4]
  wire [31:0] x626_sum_1_io_a; // @[Math.scala 150:24:@45115.4]
  wire [31:0] x626_sum_1_io_b; // @[Math.scala 150:24:@45115.4]
  wire  x626_sum_1_io_flow; // @[Math.scala 150:24:@45115.4]
  wire [31:0] x626_sum_1_io_result; // @[Math.scala 150:24:@45115.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@45125.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@45125.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@45125.4]
  wire [31:0] RetimeWrapper_64_io_in; // @[package.scala 93:22:@45125.4]
  wire [31:0] RetimeWrapper_64_io_out; // @[package.scala 93:22:@45125.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@45134.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@45134.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@45134.4]
  wire [31:0] RetimeWrapper_65_io_in; // @[package.scala 93:22:@45134.4]
  wire [31:0] RetimeWrapper_65_io_out; // @[package.scala 93:22:@45134.4]
  wire  x411_sum_1_clock; // @[Math.scala 150:24:@45143.4]
  wire  x411_sum_1_reset; // @[Math.scala 150:24:@45143.4]
  wire [31:0] x411_sum_1_io_a; // @[Math.scala 150:24:@45143.4]
  wire [31:0] x411_sum_1_io_b; // @[Math.scala 150:24:@45143.4]
  wire  x411_sum_1_io_flow; // @[Math.scala 150:24:@45143.4]
  wire [31:0] x411_sum_1_io_result; // @[Math.scala 150:24:@45143.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@45153.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@45153.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@45153.4]
  wire [31:0] RetimeWrapper_66_io_in; // @[package.scala 93:22:@45153.4]
  wire [31:0] RetimeWrapper_66_io_out; // @[package.scala 93:22:@45153.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@45162.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@45162.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@45162.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@45162.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@45162.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@45174.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@45174.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@45174.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@45174.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@45174.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@45201.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@45201.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@45201.4]
  wire [31:0] RetimeWrapper_69_io_in; // @[package.scala 93:22:@45201.4]
  wire [31:0] RetimeWrapper_69_io_out; // @[package.scala 93:22:@45201.4]
  wire  x416_sum_1_clock; // @[Math.scala 150:24:@45210.4]
  wire  x416_sum_1_reset; // @[Math.scala 150:24:@45210.4]
  wire [31:0] x416_sum_1_io_a; // @[Math.scala 150:24:@45210.4]
  wire [31:0] x416_sum_1_io_b; // @[Math.scala 150:24:@45210.4]
  wire  x416_sum_1_io_flow; // @[Math.scala 150:24:@45210.4]
  wire [31:0] x416_sum_1_io_result; // @[Math.scala 150:24:@45210.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@45220.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@45220.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@45220.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@45220.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@45220.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@45232.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@45232.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@45232.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@45232.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@45232.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@45259.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@45259.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@45259.4]
  wire [31:0] RetimeWrapper_72_io_in; // @[package.scala 93:22:@45259.4]
  wire [31:0] RetimeWrapper_72_io_out; // @[package.scala 93:22:@45259.4]
  wire  x421_sum_1_clock; // @[Math.scala 150:24:@45268.4]
  wire  x421_sum_1_reset; // @[Math.scala 150:24:@45268.4]
  wire [31:0] x421_sum_1_io_a; // @[Math.scala 150:24:@45268.4]
  wire [31:0] x421_sum_1_io_b; // @[Math.scala 150:24:@45268.4]
  wire  x421_sum_1_io_flow; // @[Math.scala 150:24:@45268.4]
  wire [31:0] x421_sum_1_io_result; // @[Math.scala 150:24:@45268.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@45278.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@45278.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@45278.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@45278.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@45278.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@45290.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@45290.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@45290.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@45290.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@45290.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@45311.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@45311.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@45311.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@45311.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@45311.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@45326.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@45326.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@45326.4]
  wire [31:0] RetimeWrapper_76_io_in; // @[package.scala 93:22:@45326.4]
  wire [31:0] RetimeWrapper_76_io_out; // @[package.scala 93:22:@45326.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@45335.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@45335.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@45335.4]
  wire [31:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@45335.4]
  wire [31:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@45335.4]
  wire  x426_sum_1_clock; // @[Math.scala 150:24:@45346.4]
  wire  x426_sum_1_reset; // @[Math.scala 150:24:@45346.4]
  wire [31:0] x426_sum_1_io_a; // @[Math.scala 150:24:@45346.4]
  wire [31:0] x426_sum_1_io_b; // @[Math.scala 150:24:@45346.4]
  wire  x426_sum_1_io_flow; // @[Math.scala 150:24:@45346.4]
  wire [31:0] x426_sum_1_io_result; // @[Math.scala 150:24:@45346.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@45356.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@45356.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@45356.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@45356.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@45356.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@45365.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@45365.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@45365.4]
  wire [31:0] RetimeWrapper_79_io_in; // @[package.scala 93:22:@45365.4]
  wire [31:0] RetimeWrapper_79_io_out; // @[package.scala 93:22:@45365.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@45377.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@45377.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@45377.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@45377.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@45377.4]
  wire  x431_sum_1_clock; // @[Math.scala 150:24:@45404.4]
  wire  x431_sum_1_reset; // @[Math.scala 150:24:@45404.4]
  wire [31:0] x431_sum_1_io_a; // @[Math.scala 150:24:@45404.4]
  wire [31:0] x431_sum_1_io_b; // @[Math.scala 150:24:@45404.4]
  wire  x431_sum_1_io_flow; // @[Math.scala 150:24:@45404.4]
  wire [31:0] x431_sum_1_io_result; // @[Math.scala 150:24:@45404.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@45414.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@45414.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@45414.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@45414.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@45414.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@45426.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@45426.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@45426.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@45426.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@45426.4]
  wire  x436_sum_1_clock; // @[Math.scala 150:24:@45453.4]
  wire  x436_sum_1_reset; // @[Math.scala 150:24:@45453.4]
  wire [31:0] x436_sum_1_io_a; // @[Math.scala 150:24:@45453.4]
  wire [31:0] x436_sum_1_io_b; // @[Math.scala 150:24:@45453.4]
  wire  x436_sum_1_io_flow; // @[Math.scala 150:24:@45453.4]
  wire [31:0] x436_sum_1_io_result; // @[Math.scala 150:24:@45453.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@45463.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@45463.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@45463.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@45463.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@45463.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@45475.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@45475.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@45475.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@45475.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@45475.4]
  wire  x439_rdrow_1_clock; // @[Math.scala 191:24:@45498.4]
  wire  x439_rdrow_1_reset; // @[Math.scala 191:24:@45498.4]
  wire [31:0] x439_rdrow_1_io_a; // @[Math.scala 191:24:@45498.4]
  wire [31:0] x439_rdrow_1_io_b; // @[Math.scala 191:24:@45498.4]
  wire  x439_rdrow_1_io_flow; // @[Math.scala 191:24:@45498.4]
  wire [31:0] x439_rdrow_1_io_result; // @[Math.scala 191:24:@45498.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@45524.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@45524.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@45524.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@45524.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@45524.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@45546.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@45546.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@45546.4]
  wire [31:0] RetimeWrapper_86_io_in; // @[package.scala 93:22:@45546.4]
  wire [31:0] RetimeWrapper_86_io_out; // @[package.scala 93:22:@45546.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@45572.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@45572.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@45572.4]
  wire [31:0] RetimeWrapper_87_io_in; // @[package.scala 93:22:@45572.4]
  wire [31:0] RetimeWrapper_87_io_out; // @[package.scala 93:22:@45572.4]
  wire  x631_sum_1_clock; // @[Math.scala 150:24:@45593.4]
  wire  x631_sum_1_reset; // @[Math.scala 150:24:@45593.4]
  wire [31:0] x631_sum_1_io_a; // @[Math.scala 150:24:@45593.4]
  wire [31:0] x631_sum_1_io_b; // @[Math.scala 150:24:@45593.4]
  wire  x631_sum_1_io_flow; // @[Math.scala 150:24:@45593.4]
  wire [31:0] x631_sum_1_io_result; // @[Math.scala 150:24:@45593.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@45603.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@45603.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@45603.4]
  wire [31:0] RetimeWrapper_88_io_in; // @[package.scala 93:22:@45603.4]
  wire [31:0] RetimeWrapper_88_io_out; // @[package.scala 93:22:@45603.4]
  wire  x447_sum_1_clock; // @[Math.scala 150:24:@45612.4]
  wire  x447_sum_1_reset; // @[Math.scala 150:24:@45612.4]
  wire [31:0] x447_sum_1_io_a; // @[Math.scala 150:24:@45612.4]
  wire [31:0] x447_sum_1_io_b; // @[Math.scala 150:24:@45612.4]
  wire  x447_sum_1_io_flow; // @[Math.scala 150:24:@45612.4]
  wire [31:0] x447_sum_1_io_result; // @[Math.scala 150:24:@45612.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@45622.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@45622.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@45622.4]
  wire [31:0] RetimeWrapper_89_io_in; // @[package.scala 93:22:@45622.4]
  wire [31:0] RetimeWrapper_89_io_out; // @[package.scala 93:22:@45622.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@45631.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@45631.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@45631.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@45631.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@45631.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@45643.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@45643.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@45643.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@45643.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@45643.4]
  wire  x452_sum_1_clock; // @[Math.scala 150:24:@45670.4]
  wire  x452_sum_1_reset; // @[Math.scala 150:24:@45670.4]
  wire [31:0] x452_sum_1_io_a; // @[Math.scala 150:24:@45670.4]
  wire [31:0] x452_sum_1_io_b; // @[Math.scala 150:24:@45670.4]
  wire  x452_sum_1_io_flow; // @[Math.scala 150:24:@45670.4]
  wire [31:0] x452_sum_1_io_result; // @[Math.scala 150:24:@45670.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@45680.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@45680.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@45680.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@45680.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@45680.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@45692.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@45692.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@45692.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@45692.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@45692.4]
  wire  x457_sum_1_clock; // @[Math.scala 150:24:@45719.4]
  wire  x457_sum_1_reset; // @[Math.scala 150:24:@45719.4]
  wire [31:0] x457_sum_1_io_a; // @[Math.scala 150:24:@45719.4]
  wire [31:0] x457_sum_1_io_b; // @[Math.scala 150:24:@45719.4]
  wire  x457_sum_1_io_flow; // @[Math.scala 150:24:@45719.4]
  wire [31:0] x457_sum_1_io_result; // @[Math.scala 150:24:@45719.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@45729.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@45729.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@45729.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@45729.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@45729.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@45741.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@45741.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@45741.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@45741.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@45741.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@45768.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@45768.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@45768.4]
  wire [31:0] RetimeWrapper_96_io_in; // @[package.scala 93:22:@45768.4]
  wire [31:0] RetimeWrapper_96_io_out; // @[package.scala 93:22:@45768.4]
  wire  x462_sum_1_clock; // @[Math.scala 150:24:@45779.4]
  wire  x462_sum_1_reset; // @[Math.scala 150:24:@45779.4]
  wire [31:0] x462_sum_1_io_a; // @[Math.scala 150:24:@45779.4]
  wire [31:0] x462_sum_1_io_b; // @[Math.scala 150:24:@45779.4]
  wire  x462_sum_1_io_flow; // @[Math.scala 150:24:@45779.4]
  wire [31:0] x462_sum_1_io_result; // @[Math.scala 150:24:@45779.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@45789.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@45789.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@45789.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@45789.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@45789.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@45798.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@45798.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@45798.4]
  wire [31:0] RetimeWrapper_98_io_in; // @[package.scala 93:22:@45798.4]
  wire [31:0] RetimeWrapper_98_io_out; // @[package.scala 93:22:@45798.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@45810.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@45810.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@45810.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@45810.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@45810.4]
  wire  x467_sum_1_clock; // @[Math.scala 150:24:@45837.4]
  wire  x467_sum_1_reset; // @[Math.scala 150:24:@45837.4]
  wire [31:0] x467_sum_1_io_a; // @[Math.scala 150:24:@45837.4]
  wire [31:0] x467_sum_1_io_b; // @[Math.scala 150:24:@45837.4]
  wire  x467_sum_1_io_flow; // @[Math.scala 150:24:@45837.4]
  wire [31:0] x467_sum_1_io_result; // @[Math.scala 150:24:@45837.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@45847.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@45847.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@45847.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@45847.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@45847.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@45859.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@45859.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@45859.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@45859.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@45859.4]
  wire  x472_sum_1_clock; // @[Math.scala 150:24:@45886.4]
  wire  x472_sum_1_reset; // @[Math.scala 150:24:@45886.4]
  wire [31:0] x472_sum_1_io_a; // @[Math.scala 150:24:@45886.4]
  wire [31:0] x472_sum_1_io_b; // @[Math.scala 150:24:@45886.4]
  wire  x472_sum_1_io_flow; // @[Math.scala 150:24:@45886.4]
  wire [31:0] x472_sum_1_io_result; // @[Math.scala 150:24:@45886.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@45896.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@45896.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@45896.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@45896.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@45896.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@45908.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@45908.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@45908.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@45908.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@45908.4]
  wire  x475_1_clock; // @[Math.scala 262:24:@45931.4]
  wire [31:0] x475_1_io_a; // @[Math.scala 262:24:@45931.4]
  wire [31:0] x475_1_io_b; // @[Math.scala 262:24:@45931.4]
  wire  x475_1_io_flow; // @[Math.scala 262:24:@45931.4]
  wire [31:0] x475_1_io_result; // @[Math.scala 262:24:@45931.4]
  wire  x476_1_clock; // @[Math.scala 262:24:@45943.4]
  wire [31:0] x476_1_io_a; // @[Math.scala 262:24:@45943.4]
  wire [31:0] x476_1_io_b; // @[Math.scala 262:24:@45943.4]
  wire  x476_1_io_flow; // @[Math.scala 262:24:@45943.4]
  wire [31:0] x476_1_io_result; // @[Math.scala 262:24:@45943.4]
  wire  x477_1_clock; // @[Math.scala 262:24:@45955.4]
  wire [31:0] x477_1_io_a; // @[Math.scala 262:24:@45955.4]
  wire [31:0] x477_1_io_b; // @[Math.scala 262:24:@45955.4]
  wire  x477_1_io_flow; // @[Math.scala 262:24:@45955.4]
  wire [31:0] x477_1_io_result; // @[Math.scala 262:24:@45955.4]
  wire  x478_1_clock; // @[Math.scala 262:24:@45967.4]
  wire [31:0] x478_1_io_a; // @[Math.scala 262:24:@45967.4]
  wire [31:0] x478_1_io_b; // @[Math.scala 262:24:@45967.4]
  wire  x478_1_io_flow; // @[Math.scala 262:24:@45967.4]
  wire [31:0] x478_1_io_result; // @[Math.scala 262:24:@45967.4]
  wire  x479_1_clock; // @[Math.scala 262:24:@45979.4]
  wire [31:0] x479_1_io_a; // @[Math.scala 262:24:@45979.4]
  wire [31:0] x479_1_io_b; // @[Math.scala 262:24:@45979.4]
  wire  x479_1_io_flow; // @[Math.scala 262:24:@45979.4]
  wire [31:0] x479_1_io_result; // @[Math.scala 262:24:@45979.4]
  wire  x480_1_clock; // @[Math.scala 262:24:@45991.4]
  wire [31:0] x480_1_io_a; // @[Math.scala 262:24:@45991.4]
  wire [31:0] x480_1_io_b; // @[Math.scala 262:24:@45991.4]
  wire  x480_1_io_flow; // @[Math.scala 262:24:@45991.4]
  wire [31:0] x480_1_io_result; // @[Math.scala 262:24:@45991.4]
  wire  x481_1_clock; // @[Math.scala 262:24:@46003.4]
  wire [31:0] x481_1_io_a; // @[Math.scala 262:24:@46003.4]
  wire [31:0] x481_1_io_b; // @[Math.scala 262:24:@46003.4]
  wire  x481_1_io_flow; // @[Math.scala 262:24:@46003.4]
  wire [31:0] x481_1_io_result; // @[Math.scala 262:24:@46003.4]
  wire  x482_1_clock; // @[Math.scala 262:24:@46015.4]
  wire [31:0] x482_1_io_a; // @[Math.scala 262:24:@46015.4]
  wire [31:0] x482_1_io_b; // @[Math.scala 262:24:@46015.4]
  wire  x482_1_io_flow; // @[Math.scala 262:24:@46015.4]
  wire [31:0] x482_1_io_result; // @[Math.scala 262:24:@46015.4]
  wire  x483_1_clock; // @[Math.scala 262:24:@46027.4]
  wire [31:0] x483_1_io_a; // @[Math.scala 262:24:@46027.4]
  wire [31:0] x483_1_io_b; // @[Math.scala 262:24:@46027.4]
  wire  x483_1_io_flow; // @[Math.scala 262:24:@46027.4]
  wire [31:0] x483_1_io_result; // @[Math.scala 262:24:@46027.4]
  wire  x484_x3_1_clock; // @[Math.scala 150:24:@46037.4]
  wire  x484_x3_1_reset; // @[Math.scala 150:24:@46037.4]
  wire [31:0] x484_x3_1_io_a; // @[Math.scala 150:24:@46037.4]
  wire [31:0] x484_x3_1_io_b; // @[Math.scala 150:24:@46037.4]
  wire  x484_x3_1_io_flow; // @[Math.scala 150:24:@46037.4]
  wire [31:0] x484_x3_1_io_result; // @[Math.scala 150:24:@46037.4]
  wire  x485_x4_1_clock; // @[Math.scala 150:24:@46047.4]
  wire  x485_x4_1_reset; // @[Math.scala 150:24:@46047.4]
  wire [31:0] x485_x4_1_io_a; // @[Math.scala 150:24:@46047.4]
  wire [31:0] x485_x4_1_io_b; // @[Math.scala 150:24:@46047.4]
  wire  x485_x4_1_io_flow; // @[Math.scala 150:24:@46047.4]
  wire [31:0] x485_x4_1_io_result; // @[Math.scala 150:24:@46047.4]
  wire  x486_x3_1_clock; // @[Math.scala 150:24:@46057.4]
  wire  x486_x3_1_reset; // @[Math.scala 150:24:@46057.4]
  wire [31:0] x486_x3_1_io_a; // @[Math.scala 150:24:@46057.4]
  wire [31:0] x486_x3_1_io_b; // @[Math.scala 150:24:@46057.4]
  wire  x486_x3_1_io_flow; // @[Math.scala 150:24:@46057.4]
  wire [31:0] x486_x3_1_io_result; // @[Math.scala 150:24:@46057.4]
  wire  x487_x4_1_clock; // @[Math.scala 150:24:@46067.4]
  wire  x487_x4_1_reset; // @[Math.scala 150:24:@46067.4]
  wire [31:0] x487_x4_1_io_a; // @[Math.scala 150:24:@46067.4]
  wire [31:0] x487_x4_1_io_b; // @[Math.scala 150:24:@46067.4]
  wire  x487_x4_1_io_flow; // @[Math.scala 150:24:@46067.4]
  wire [31:0] x487_x4_1_io_result; // @[Math.scala 150:24:@46067.4]
  wire  x488_x3_1_clock; // @[Math.scala 150:24:@46077.4]
  wire  x488_x3_1_reset; // @[Math.scala 150:24:@46077.4]
  wire [31:0] x488_x3_1_io_a; // @[Math.scala 150:24:@46077.4]
  wire [31:0] x488_x3_1_io_b; // @[Math.scala 150:24:@46077.4]
  wire  x488_x3_1_io_flow; // @[Math.scala 150:24:@46077.4]
  wire [31:0] x488_x3_1_io_result; // @[Math.scala 150:24:@46077.4]
  wire  x489_x4_1_clock; // @[Math.scala 150:24:@46087.4]
  wire  x489_x4_1_reset; // @[Math.scala 150:24:@46087.4]
  wire [31:0] x489_x4_1_io_a; // @[Math.scala 150:24:@46087.4]
  wire [31:0] x489_x4_1_io_b; // @[Math.scala 150:24:@46087.4]
  wire  x489_x4_1_io_flow; // @[Math.scala 150:24:@46087.4]
  wire [31:0] x489_x4_1_io_result; // @[Math.scala 150:24:@46087.4]
  wire  x490_x3_1_clock; // @[Math.scala 150:24:@46097.4]
  wire  x490_x3_1_reset; // @[Math.scala 150:24:@46097.4]
  wire [31:0] x490_x3_1_io_a; // @[Math.scala 150:24:@46097.4]
  wire [31:0] x490_x3_1_io_b; // @[Math.scala 150:24:@46097.4]
  wire  x490_x3_1_io_flow; // @[Math.scala 150:24:@46097.4]
  wire [31:0] x490_x3_1_io_result; // @[Math.scala 150:24:@46097.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@46107.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@46107.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@46107.4]
  wire [31:0] RetimeWrapper_104_io_in; // @[package.scala 93:22:@46107.4]
  wire [31:0] RetimeWrapper_104_io_out; // @[package.scala 93:22:@46107.4]
  wire  x491_sum_1_clock; // @[Math.scala 150:24:@46116.4]
  wire  x491_sum_1_reset; // @[Math.scala 150:24:@46116.4]
  wire [31:0] x491_sum_1_io_a; // @[Math.scala 150:24:@46116.4]
  wire [31:0] x491_sum_1_io_b; // @[Math.scala 150:24:@46116.4]
  wire  x491_sum_1_io_flow; // @[Math.scala 150:24:@46116.4]
  wire [31:0] x491_sum_1_io_result; // @[Math.scala 150:24:@46116.4]
  wire [31:0] x492_1_io_b; // @[Math.scala 720:24:@46126.4]
  wire [31:0] x492_1_io_result; // @[Math.scala 720:24:@46126.4]
  wire  x493_mul_1_clock; // @[Math.scala 262:24:@46137.4]
  wire [31:0] x493_mul_1_io_a; // @[Math.scala 262:24:@46137.4]
  wire  x493_mul_1_io_flow; // @[Math.scala 262:24:@46137.4]
  wire [31:0] x493_mul_1_io_result; // @[Math.scala 262:24:@46137.4]
  wire [31:0] x494_1_io_b; // @[Math.scala 720:24:@46147.4]
  wire [31:0] x494_1_io_result; // @[Math.scala 720:24:@46147.4]
  wire  x495_1_clock; // @[Math.scala 262:24:@46158.4]
  wire [31:0] x495_1_io_a; // @[Math.scala 262:24:@46158.4]
  wire [31:0] x495_1_io_b; // @[Math.scala 262:24:@46158.4]
  wire  x495_1_io_flow; // @[Math.scala 262:24:@46158.4]
  wire [31:0] x495_1_io_result; // @[Math.scala 262:24:@46158.4]
  wire  x496_1_clock; // @[Math.scala 262:24:@46170.4]
  wire [31:0] x496_1_io_a; // @[Math.scala 262:24:@46170.4]
  wire [31:0] x496_1_io_b; // @[Math.scala 262:24:@46170.4]
  wire  x496_1_io_flow; // @[Math.scala 262:24:@46170.4]
  wire [31:0] x496_1_io_result; // @[Math.scala 262:24:@46170.4]
  wire  x497_1_clock; // @[Math.scala 262:24:@46182.4]
  wire [31:0] x497_1_io_a; // @[Math.scala 262:24:@46182.4]
  wire [31:0] x497_1_io_b; // @[Math.scala 262:24:@46182.4]
  wire  x497_1_io_flow; // @[Math.scala 262:24:@46182.4]
  wire [31:0] x497_1_io_result; // @[Math.scala 262:24:@46182.4]
  wire  x498_1_clock; // @[Math.scala 262:24:@46194.4]
  wire [31:0] x498_1_io_a; // @[Math.scala 262:24:@46194.4]
  wire [31:0] x498_1_io_b; // @[Math.scala 262:24:@46194.4]
  wire  x498_1_io_flow; // @[Math.scala 262:24:@46194.4]
  wire [31:0] x498_1_io_result; // @[Math.scala 262:24:@46194.4]
  wire  x499_1_clock; // @[Math.scala 262:24:@46206.4]
  wire [31:0] x499_1_io_a; // @[Math.scala 262:24:@46206.4]
  wire [31:0] x499_1_io_b; // @[Math.scala 262:24:@46206.4]
  wire  x499_1_io_flow; // @[Math.scala 262:24:@46206.4]
  wire [31:0] x499_1_io_result; // @[Math.scala 262:24:@46206.4]
  wire  x500_1_clock; // @[Math.scala 262:24:@46218.4]
  wire [31:0] x500_1_io_a; // @[Math.scala 262:24:@46218.4]
  wire [31:0] x500_1_io_b; // @[Math.scala 262:24:@46218.4]
  wire  x500_1_io_flow; // @[Math.scala 262:24:@46218.4]
  wire [31:0] x500_1_io_result; // @[Math.scala 262:24:@46218.4]
  wire  x501_1_clock; // @[Math.scala 262:24:@46232.4]
  wire [31:0] x501_1_io_a; // @[Math.scala 262:24:@46232.4]
  wire [31:0] x501_1_io_b; // @[Math.scala 262:24:@46232.4]
  wire  x501_1_io_flow; // @[Math.scala 262:24:@46232.4]
  wire [31:0] x501_1_io_result; // @[Math.scala 262:24:@46232.4]
  wire  x502_1_clock; // @[Math.scala 262:24:@46244.4]
  wire [31:0] x502_1_io_a; // @[Math.scala 262:24:@46244.4]
  wire [31:0] x502_1_io_b; // @[Math.scala 262:24:@46244.4]
  wire  x502_1_io_flow; // @[Math.scala 262:24:@46244.4]
  wire [31:0] x502_1_io_result; // @[Math.scala 262:24:@46244.4]
  wire  x503_1_clock; // @[Math.scala 262:24:@46256.4]
  wire [31:0] x503_1_io_a; // @[Math.scala 262:24:@46256.4]
  wire [31:0] x503_1_io_b; // @[Math.scala 262:24:@46256.4]
  wire  x503_1_io_flow; // @[Math.scala 262:24:@46256.4]
  wire [31:0] x503_1_io_result; // @[Math.scala 262:24:@46256.4]
  wire  x504_x3_1_clock; // @[Math.scala 150:24:@46266.4]
  wire  x504_x3_1_reset; // @[Math.scala 150:24:@46266.4]
  wire [31:0] x504_x3_1_io_a; // @[Math.scala 150:24:@46266.4]
  wire [31:0] x504_x3_1_io_b; // @[Math.scala 150:24:@46266.4]
  wire  x504_x3_1_io_flow; // @[Math.scala 150:24:@46266.4]
  wire [31:0] x504_x3_1_io_result; // @[Math.scala 150:24:@46266.4]
  wire  x505_x4_1_clock; // @[Math.scala 150:24:@46276.4]
  wire  x505_x4_1_reset; // @[Math.scala 150:24:@46276.4]
  wire [31:0] x505_x4_1_io_a; // @[Math.scala 150:24:@46276.4]
  wire [31:0] x505_x4_1_io_b; // @[Math.scala 150:24:@46276.4]
  wire  x505_x4_1_io_flow; // @[Math.scala 150:24:@46276.4]
  wire [31:0] x505_x4_1_io_result; // @[Math.scala 150:24:@46276.4]
  wire  x506_x3_1_clock; // @[Math.scala 150:24:@46286.4]
  wire  x506_x3_1_reset; // @[Math.scala 150:24:@46286.4]
  wire [31:0] x506_x3_1_io_a; // @[Math.scala 150:24:@46286.4]
  wire [31:0] x506_x3_1_io_b; // @[Math.scala 150:24:@46286.4]
  wire  x506_x3_1_io_flow; // @[Math.scala 150:24:@46286.4]
  wire [31:0] x506_x3_1_io_result; // @[Math.scala 150:24:@46286.4]
  wire  x507_x4_1_clock; // @[Math.scala 150:24:@46296.4]
  wire  x507_x4_1_reset; // @[Math.scala 150:24:@46296.4]
  wire [31:0] x507_x4_1_io_a; // @[Math.scala 150:24:@46296.4]
  wire [31:0] x507_x4_1_io_b; // @[Math.scala 150:24:@46296.4]
  wire  x507_x4_1_io_flow; // @[Math.scala 150:24:@46296.4]
  wire [31:0] x507_x4_1_io_result; // @[Math.scala 150:24:@46296.4]
  wire  x508_x3_1_clock; // @[Math.scala 150:24:@46306.4]
  wire  x508_x3_1_reset; // @[Math.scala 150:24:@46306.4]
  wire [31:0] x508_x3_1_io_a; // @[Math.scala 150:24:@46306.4]
  wire [31:0] x508_x3_1_io_b; // @[Math.scala 150:24:@46306.4]
  wire  x508_x3_1_io_flow; // @[Math.scala 150:24:@46306.4]
  wire [31:0] x508_x3_1_io_result; // @[Math.scala 150:24:@46306.4]
  wire  x509_x4_1_clock; // @[Math.scala 150:24:@46316.4]
  wire  x509_x4_1_reset; // @[Math.scala 150:24:@46316.4]
  wire [31:0] x509_x4_1_io_a; // @[Math.scala 150:24:@46316.4]
  wire [31:0] x509_x4_1_io_b; // @[Math.scala 150:24:@46316.4]
  wire  x509_x4_1_io_flow; // @[Math.scala 150:24:@46316.4]
  wire [31:0] x509_x4_1_io_result; // @[Math.scala 150:24:@46316.4]
  wire  x510_x3_1_clock; // @[Math.scala 150:24:@46326.4]
  wire  x510_x3_1_reset; // @[Math.scala 150:24:@46326.4]
  wire [31:0] x510_x3_1_io_a; // @[Math.scala 150:24:@46326.4]
  wire [31:0] x510_x3_1_io_b; // @[Math.scala 150:24:@46326.4]
  wire  x510_x3_1_io_flow; // @[Math.scala 150:24:@46326.4]
  wire [31:0] x510_x3_1_io_result; // @[Math.scala 150:24:@46326.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@46336.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@46336.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@46336.4]
  wire [31:0] RetimeWrapper_105_io_in; // @[package.scala 93:22:@46336.4]
  wire [31:0] RetimeWrapper_105_io_out; // @[package.scala 93:22:@46336.4]
  wire  x511_sum_1_clock; // @[Math.scala 150:24:@46345.4]
  wire  x511_sum_1_reset; // @[Math.scala 150:24:@46345.4]
  wire [31:0] x511_sum_1_io_a; // @[Math.scala 150:24:@46345.4]
  wire [31:0] x511_sum_1_io_b; // @[Math.scala 150:24:@46345.4]
  wire  x511_sum_1_io_flow; // @[Math.scala 150:24:@46345.4]
  wire [31:0] x511_sum_1_io_result; // @[Math.scala 150:24:@46345.4]
  wire [31:0] x512_1_io_b; // @[Math.scala 720:24:@46355.4]
  wire [31:0] x512_1_io_result; // @[Math.scala 720:24:@46355.4]
  wire  x513_mul_1_clock; // @[Math.scala 262:24:@46366.4]
  wire [31:0] x513_mul_1_io_a; // @[Math.scala 262:24:@46366.4]
  wire  x513_mul_1_io_flow; // @[Math.scala 262:24:@46366.4]
  wire [31:0] x513_mul_1_io_result; // @[Math.scala 262:24:@46366.4]
  wire [31:0] x514_1_io_b; // @[Math.scala 720:24:@46376.4]
  wire [31:0] x514_1_io_result; // @[Math.scala 720:24:@46376.4]
  wire  x515_1_clock; // @[Math.scala 262:24:@46387.4]
  wire [31:0] x515_1_io_a; // @[Math.scala 262:24:@46387.4]
  wire [31:0] x515_1_io_b; // @[Math.scala 262:24:@46387.4]
  wire  x515_1_io_flow; // @[Math.scala 262:24:@46387.4]
  wire [31:0] x515_1_io_result; // @[Math.scala 262:24:@46387.4]
  wire  x516_1_clock; // @[Math.scala 262:24:@46399.4]
  wire [31:0] x516_1_io_a; // @[Math.scala 262:24:@46399.4]
  wire [31:0] x516_1_io_b; // @[Math.scala 262:24:@46399.4]
  wire  x516_1_io_flow; // @[Math.scala 262:24:@46399.4]
  wire [31:0] x516_1_io_result; // @[Math.scala 262:24:@46399.4]
  wire  x517_1_clock; // @[Math.scala 262:24:@46411.4]
  wire [31:0] x517_1_io_a; // @[Math.scala 262:24:@46411.4]
  wire [31:0] x517_1_io_b; // @[Math.scala 262:24:@46411.4]
  wire  x517_1_io_flow; // @[Math.scala 262:24:@46411.4]
  wire [31:0] x517_1_io_result; // @[Math.scala 262:24:@46411.4]
  wire  x518_1_clock; // @[Math.scala 262:24:@46423.4]
  wire [31:0] x518_1_io_a; // @[Math.scala 262:24:@46423.4]
  wire [31:0] x518_1_io_b; // @[Math.scala 262:24:@46423.4]
  wire  x518_1_io_flow; // @[Math.scala 262:24:@46423.4]
  wire [31:0] x518_1_io_result; // @[Math.scala 262:24:@46423.4]
  wire  x519_1_clock; // @[Math.scala 262:24:@46435.4]
  wire [31:0] x519_1_io_a; // @[Math.scala 262:24:@46435.4]
  wire [31:0] x519_1_io_b; // @[Math.scala 262:24:@46435.4]
  wire  x519_1_io_flow; // @[Math.scala 262:24:@46435.4]
  wire [31:0] x519_1_io_result; // @[Math.scala 262:24:@46435.4]
  wire  x520_1_clock; // @[Math.scala 262:24:@46447.4]
  wire [31:0] x520_1_io_a; // @[Math.scala 262:24:@46447.4]
  wire [31:0] x520_1_io_b; // @[Math.scala 262:24:@46447.4]
  wire  x520_1_io_flow; // @[Math.scala 262:24:@46447.4]
  wire [31:0] x520_1_io_result; // @[Math.scala 262:24:@46447.4]
  wire  x521_x3_1_clock; // @[Math.scala 150:24:@46457.4]
  wire  x521_x3_1_reset; // @[Math.scala 150:24:@46457.4]
  wire [31:0] x521_x3_1_io_a; // @[Math.scala 150:24:@46457.4]
  wire [31:0] x521_x3_1_io_b; // @[Math.scala 150:24:@46457.4]
  wire  x521_x3_1_io_flow; // @[Math.scala 150:24:@46457.4]
  wire [31:0] x521_x3_1_io_result; // @[Math.scala 150:24:@46457.4]
  wire  x522_x4_1_clock; // @[Math.scala 150:24:@46467.4]
  wire  x522_x4_1_reset; // @[Math.scala 150:24:@46467.4]
  wire [31:0] x522_x4_1_io_a; // @[Math.scala 150:24:@46467.4]
  wire [31:0] x522_x4_1_io_b; // @[Math.scala 150:24:@46467.4]
  wire  x522_x4_1_io_flow; // @[Math.scala 150:24:@46467.4]
  wire [31:0] x522_x4_1_io_result; // @[Math.scala 150:24:@46467.4]
  wire  x523_x3_1_clock; // @[Math.scala 150:24:@46477.4]
  wire  x523_x3_1_reset; // @[Math.scala 150:24:@46477.4]
  wire [31:0] x523_x3_1_io_a; // @[Math.scala 150:24:@46477.4]
  wire [31:0] x523_x3_1_io_b; // @[Math.scala 150:24:@46477.4]
  wire  x523_x3_1_io_flow; // @[Math.scala 150:24:@46477.4]
  wire [31:0] x523_x3_1_io_result; // @[Math.scala 150:24:@46477.4]
  wire  x524_x4_1_clock; // @[Math.scala 150:24:@46487.4]
  wire  x524_x4_1_reset; // @[Math.scala 150:24:@46487.4]
  wire [31:0] x524_x4_1_io_a; // @[Math.scala 150:24:@46487.4]
  wire [31:0] x524_x4_1_io_b; // @[Math.scala 150:24:@46487.4]
  wire  x524_x4_1_io_flow; // @[Math.scala 150:24:@46487.4]
  wire [31:0] x524_x4_1_io_result; // @[Math.scala 150:24:@46487.4]
  wire  x525_x3_1_clock; // @[Math.scala 150:24:@46497.4]
  wire  x525_x3_1_reset; // @[Math.scala 150:24:@46497.4]
  wire [31:0] x525_x3_1_io_a; // @[Math.scala 150:24:@46497.4]
  wire [31:0] x525_x3_1_io_b; // @[Math.scala 150:24:@46497.4]
  wire  x525_x3_1_io_flow; // @[Math.scala 150:24:@46497.4]
  wire [31:0] x525_x3_1_io_result; // @[Math.scala 150:24:@46497.4]
  wire  x526_x4_1_clock; // @[Math.scala 150:24:@46507.4]
  wire  x526_x4_1_reset; // @[Math.scala 150:24:@46507.4]
  wire [31:0] x526_x4_1_io_a; // @[Math.scala 150:24:@46507.4]
  wire [31:0] x526_x4_1_io_b; // @[Math.scala 150:24:@46507.4]
  wire  x526_x4_1_io_flow; // @[Math.scala 150:24:@46507.4]
  wire [31:0] x526_x4_1_io_result; // @[Math.scala 150:24:@46507.4]
  wire  x527_x3_1_clock; // @[Math.scala 150:24:@46517.4]
  wire  x527_x3_1_reset; // @[Math.scala 150:24:@46517.4]
  wire [31:0] x527_x3_1_io_a; // @[Math.scala 150:24:@46517.4]
  wire [31:0] x527_x3_1_io_b; // @[Math.scala 150:24:@46517.4]
  wire  x527_x3_1_io_flow; // @[Math.scala 150:24:@46517.4]
  wire [31:0] x527_x3_1_io_result; // @[Math.scala 150:24:@46517.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@46527.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@46527.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@46527.4]
  wire [31:0] RetimeWrapper_106_io_in; // @[package.scala 93:22:@46527.4]
  wire [31:0] RetimeWrapper_106_io_out; // @[package.scala 93:22:@46527.4]
  wire  x528_sum_1_clock; // @[Math.scala 150:24:@46536.4]
  wire  x528_sum_1_reset; // @[Math.scala 150:24:@46536.4]
  wire [31:0] x528_sum_1_io_a; // @[Math.scala 150:24:@46536.4]
  wire [31:0] x528_sum_1_io_b; // @[Math.scala 150:24:@46536.4]
  wire  x528_sum_1_io_flow; // @[Math.scala 150:24:@46536.4]
  wire [31:0] x528_sum_1_io_result; // @[Math.scala 150:24:@46536.4]
  wire [31:0] x529_1_io_b; // @[Math.scala 720:24:@46546.4]
  wire [31:0] x529_1_io_result; // @[Math.scala 720:24:@46546.4]
  wire  x530_mul_1_clock; // @[Math.scala 262:24:@46557.4]
  wire [31:0] x530_mul_1_io_a; // @[Math.scala 262:24:@46557.4]
  wire  x530_mul_1_io_flow; // @[Math.scala 262:24:@46557.4]
  wire [31:0] x530_mul_1_io_result; // @[Math.scala 262:24:@46557.4]
  wire [31:0] x531_1_io_b; // @[Math.scala 720:24:@46567.4]
  wire [31:0] x531_1_io_result; // @[Math.scala 720:24:@46567.4]
  wire  x532_1_clock; // @[Math.scala 262:24:@46578.4]
  wire [31:0] x532_1_io_a; // @[Math.scala 262:24:@46578.4]
  wire [31:0] x532_1_io_b; // @[Math.scala 262:24:@46578.4]
  wire  x532_1_io_flow; // @[Math.scala 262:24:@46578.4]
  wire [31:0] x532_1_io_result; // @[Math.scala 262:24:@46578.4]
  wire  x533_1_clock; // @[Math.scala 262:24:@46590.4]
  wire [31:0] x533_1_io_a; // @[Math.scala 262:24:@46590.4]
  wire [31:0] x533_1_io_b; // @[Math.scala 262:24:@46590.4]
  wire  x533_1_io_flow; // @[Math.scala 262:24:@46590.4]
  wire [31:0] x533_1_io_result; // @[Math.scala 262:24:@46590.4]
  wire  x534_1_clock; // @[Math.scala 262:24:@46602.4]
  wire [31:0] x534_1_io_a; // @[Math.scala 262:24:@46602.4]
  wire [31:0] x534_1_io_b; // @[Math.scala 262:24:@46602.4]
  wire  x534_1_io_flow; // @[Math.scala 262:24:@46602.4]
  wire [31:0] x534_1_io_result; // @[Math.scala 262:24:@46602.4]
  wire  x535_1_clock; // @[Math.scala 262:24:@46614.4]
  wire [31:0] x535_1_io_a; // @[Math.scala 262:24:@46614.4]
  wire [31:0] x535_1_io_b; // @[Math.scala 262:24:@46614.4]
  wire  x535_1_io_flow; // @[Math.scala 262:24:@46614.4]
  wire [31:0] x535_1_io_result; // @[Math.scala 262:24:@46614.4]
  wire  x536_1_clock; // @[Math.scala 262:24:@46626.4]
  wire [31:0] x536_1_io_a; // @[Math.scala 262:24:@46626.4]
  wire [31:0] x536_1_io_b; // @[Math.scala 262:24:@46626.4]
  wire  x536_1_io_flow; // @[Math.scala 262:24:@46626.4]
  wire [31:0] x536_1_io_result; // @[Math.scala 262:24:@46626.4]
  wire  x537_1_clock; // @[Math.scala 262:24:@46638.4]
  wire [31:0] x537_1_io_a; // @[Math.scala 262:24:@46638.4]
  wire [31:0] x537_1_io_b; // @[Math.scala 262:24:@46638.4]
  wire  x537_1_io_flow; // @[Math.scala 262:24:@46638.4]
  wire [31:0] x537_1_io_result; // @[Math.scala 262:24:@46638.4]
  wire  x538_x3_1_clock; // @[Math.scala 150:24:@46648.4]
  wire  x538_x3_1_reset; // @[Math.scala 150:24:@46648.4]
  wire [31:0] x538_x3_1_io_a; // @[Math.scala 150:24:@46648.4]
  wire [31:0] x538_x3_1_io_b; // @[Math.scala 150:24:@46648.4]
  wire  x538_x3_1_io_flow; // @[Math.scala 150:24:@46648.4]
  wire [31:0] x538_x3_1_io_result; // @[Math.scala 150:24:@46648.4]
  wire  x539_x4_1_clock; // @[Math.scala 150:24:@46658.4]
  wire  x539_x4_1_reset; // @[Math.scala 150:24:@46658.4]
  wire [31:0] x539_x4_1_io_a; // @[Math.scala 150:24:@46658.4]
  wire [31:0] x539_x4_1_io_b; // @[Math.scala 150:24:@46658.4]
  wire  x539_x4_1_io_flow; // @[Math.scala 150:24:@46658.4]
  wire [31:0] x539_x4_1_io_result; // @[Math.scala 150:24:@46658.4]
  wire  x540_x3_1_clock; // @[Math.scala 150:24:@46668.4]
  wire  x540_x3_1_reset; // @[Math.scala 150:24:@46668.4]
  wire [31:0] x540_x3_1_io_a; // @[Math.scala 150:24:@46668.4]
  wire [31:0] x540_x3_1_io_b; // @[Math.scala 150:24:@46668.4]
  wire  x540_x3_1_io_flow; // @[Math.scala 150:24:@46668.4]
  wire [31:0] x540_x3_1_io_result; // @[Math.scala 150:24:@46668.4]
  wire  x541_x4_1_clock; // @[Math.scala 150:24:@46678.4]
  wire  x541_x4_1_reset; // @[Math.scala 150:24:@46678.4]
  wire [31:0] x541_x4_1_io_a; // @[Math.scala 150:24:@46678.4]
  wire [31:0] x541_x4_1_io_b; // @[Math.scala 150:24:@46678.4]
  wire  x541_x4_1_io_flow; // @[Math.scala 150:24:@46678.4]
  wire [31:0] x541_x4_1_io_result; // @[Math.scala 150:24:@46678.4]
  wire  x542_x3_1_clock; // @[Math.scala 150:24:@46688.4]
  wire  x542_x3_1_reset; // @[Math.scala 150:24:@46688.4]
  wire [31:0] x542_x3_1_io_a; // @[Math.scala 150:24:@46688.4]
  wire [31:0] x542_x3_1_io_b; // @[Math.scala 150:24:@46688.4]
  wire  x542_x3_1_io_flow; // @[Math.scala 150:24:@46688.4]
  wire [31:0] x542_x3_1_io_result; // @[Math.scala 150:24:@46688.4]
  wire  x543_x4_1_clock; // @[Math.scala 150:24:@46698.4]
  wire  x543_x4_1_reset; // @[Math.scala 150:24:@46698.4]
  wire [31:0] x543_x4_1_io_a; // @[Math.scala 150:24:@46698.4]
  wire [31:0] x543_x4_1_io_b; // @[Math.scala 150:24:@46698.4]
  wire  x543_x4_1_io_flow; // @[Math.scala 150:24:@46698.4]
  wire [31:0] x543_x4_1_io_result; // @[Math.scala 150:24:@46698.4]
  wire  x544_x3_1_clock; // @[Math.scala 150:24:@46708.4]
  wire  x544_x3_1_reset; // @[Math.scala 150:24:@46708.4]
  wire [31:0] x544_x3_1_io_a; // @[Math.scala 150:24:@46708.4]
  wire [31:0] x544_x3_1_io_b; // @[Math.scala 150:24:@46708.4]
  wire  x544_x3_1_io_flow; // @[Math.scala 150:24:@46708.4]
  wire [31:0] x544_x3_1_io_result; // @[Math.scala 150:24:@46708.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@46718.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@46718.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@46718.4]
  wire [31:0] RetimeWrapper_107_io_in; // @[package.scala 93:22:@46718.4]
  wire [31:0] RetimeWrapper_107_io_out; // @[package.scala 93:22:@46718.4]
  wire  x545_sum_1_clock; // @[Math.scala 150:24:@46727.4]
  wire  x545_sum_1_reset; // @[Math.scala 150:24:@46727.4]
  wire [31:0] x545_sum_1_io_a; // @[Math.scala 150:24:@46727.4]
  wire [31:0] x545_sum_1_io_b; // @[Math.scala 150:24:@46727.4]
  wire  x545_sum_1_io_flow; // @[Math.scala 150:24:@46727.4]
  wire [31:0] x545_sum_1_io_result; // @[Math.scala 150:24:@46727.4]
  wire [31:0] x546_1_io_b; // @[Math.scala 720:24:@46737.4]
  wire [31:0] x546_1_io_result; // @[Math.scala 720:24:@46737.4]
  wire  x547_mul_1_clock; // @[Math.scala 262:24:@46750.4]
  wire [31:0] x547_mul_1_io_a; // @[Math.scala 262:24:@46750.4]
  wire  x547_mul_1_io_flow; // @[Math.scala 262:24:@46750.4]
  wire [31:0] x547_mul_1_io_result; // @[Math.scala 262:24:@46750.4]
  wire [31:0] x548_1_io_b; // @[Math.scala 720:24:@46760.4]
  wire [31:0] x548_1_io_result; // @[Math.scala 720:24:@46760.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@46779.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@46779.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@46779.4]
  wire [127:0] RetimeWrapper_108_io_in; // @[package.scala 93:22:@46779.4]
  wire [127:0] RetimeWrapper_108_io_out; // @[package.scala 93:22:@46779.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@46788.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@46788.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@46788.4]
  wire  RetimeWrapper_109_io_in; // @[package.scala 93:22:@46788.4]
  wire  RetimeWrapper_109_io_out; // @[package.scala 93:22:@46788.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@46797.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@46797.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@46797.4]
  wire  RetimeWrapper_110_io_in; // @[package.scala 93:22:@46797.4]
  wire  RetimeWrapper_110_io_out; // @[package.scala 93:22:@46797.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@46806.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@46806.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@46806.4]
  wire  RetimeWrapper_111_io_in; // @[package.scala 93:22:@46806.4]
  wire  RetimeWrapper_111_io_out; // @[package.scala 93:22:@46806.4]
  wire  b330; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 62:18:@43744.4]
  wire  b331; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 63:18:@43745.4]
  wire  _T_205; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 67:30:@43747.4]
  wire  _T_206; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 67:37:@43748.4]
  wire  _T_210; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 69:76:@43753.4]
  wire  _T_211; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 69:62:@43754.4]
  wire  _T_213; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 69:101:@43755.4]
  wire [127:0] x637_x332_D1_0_number; // @[package.scala 96:25:@43764.4 package.scala 96:25:@43765.4]
  wire [31:0] b328_number; // @[Math.scala 723:22:@43729.4 Math.scala 724:14:@43730.4]
  wire [31:0] _T_247; // @[Math.scala 406:49:@43929.4]
  wire [31:0] _T_249; // @[Math.scala 406:56:@43931.4]
  wire [31:0] _T_250; // @[Math.scala 406:56:@43932.4]
  wire [31:0] x617_number; // @[implicits.scala 133:21:@43933.4]
  wire [31:0] _T_260; // @[Math.scala 406:49:@43942.4]
  wire [31:0] _T_262; // @[Math.scala 406:56:@43944.4]
  wire [31:0] _T_263; // @[Math.scala 406:56:@43945.4]
  wire  _T_274; // @[FixedPoint.scala 50:25:@43963.4]
  wire [1:0] _T_278; // @[Bitwise.scala 72:12:@43965.4]
  wire [29:0] _T_279; // @[FixedPoint.scala 18:52:@43966.4]
  wire  _T_285; // @[Math.scala 451:55:@43968.4]
  wire [1:0] _T_286; // @[FixedPoint.scala 18:52:@43969.4]
  wire  _T_292; // @[Math.scala 451:110:@43971.4]
  wire  _T_293; // @[Math.scala 451:94:@43972.4]
  wire [31:0] _T_295; // @[Cat.scala 30:58:@43974.4]
  wire [31:0] x340_1_number; // @[Math.scala 454:20:@43975.4]
  wire [39:0] _GEN_0; // @[Math.scala 461:32:@43980.4]
  wire [39:0] _T_300; // @[Math.scala 461:32:@43980.4]
  wire [37:0] _GEN_1; // @[Math.scala 461:32:@43985.4]
  wire [37:0] _T_303; // @[Math.scala 461:32:@43985.4]
  wire  _T_339; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 117:101:@44083.4]
  wire  _T_343; // @[package.scala 96:25:@44091.4 package.scala 96:25:@44092.4]
  wire  _T_345; // @[implicits.scala 55:10:@44093.4]
  wire  _T_346; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 117:118:@44094.4]
  wire  _T_348; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 117:207:@44096.4]
  wire  _T_349; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 117:226:@44097.4]
  wire  x642_b330_D24; // @[package.scala 96:25:@44062.4 package.scala 96:25:@44063.4]
  wire  _T_350; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 117:252:@44098.4]
  wire  x643_b331_D24; // @[package.scala 96:25:@44071.4 package.scala 96:25:@44072.4]
  wire  _T_394; // @[package.scala 96:25:@44198.4 package.scala 96:25:@44199.4]
  wire  _T_396; // @[implicits.scala 55:10:@44200.4]
  wire  _T_397; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 140:118:@44201.4]
  wire  _T_399; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 140:207:@44203.4]
  wire  _T_400; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 140:226:@44204.4]
  wire  _T_401; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 140:252:@44205.4]
  wire  _T_442; // @[package.scala 96:25:@44296.4 package.scala 96:25:@44297.4]
  wire  _T_444; // @[implicits.scala 55:10:@44298.4]
  wire  _T_445; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 161:118:@44299.4]
  wire  _T_447; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 161:207:@44301.4]
  wire  _T_448; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 161:226:@44302.4]
  wire  _T_449; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 161:252:@44303.4]
  wire  _T_490; // @[package.scala 96:25:@44394.4 package.scala 96:25:@44395.4]
  wire  _T_492; // @[implicits.scala 55:10:@44396.4]
  wire  _T_493; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 188:166:@44397.4]
  wire  _T_495; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 188:255:@44399.4]
  wire  _T_496; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 188:274:@44400.4]
  wire  _T_497; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 188:300:@44401.4]
  wire [31:0] x655_b328_D26_number; // @[package.scala 96:25:@44415.4 package.scala 96:25:@44416.4]
  wire [31:0] _T_509; // @[Math.scala 476:37:@44423.4]
  wire [31:0] x656_x357_rdcol_D26_number; // @[package.scala 96:25:@44440.4 package.scala 96:25:@44441.4]
  wire [31:0] _T_522; // @[Math.scala 476:37:@44446.4]
  wire  x657_x364_D1; // @[package.scala 96:25:@44463.4 package.scala 96:25:@44464.4]
  wire  x365; // @[package.scala 96:25:@44454.4 package.scala 96:25:@44455.4]
  wire  x366; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 203:24:@44467.4]
  wire  _T_563; // @[package.scala 96:25:@44535.4 package.scala 96:25:@44536.4]
  wire  _T_565; // @[implicits.scala 55:10:@44537.4]
  wire  _T_566; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 222:194:@44538.4]
  wire  x660_x367_D20; // @[package.scala 96:25:@44496.4 package.scala 96:25:@44497.4]
  wire  _T_567; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 222:283:@44539.4]
  wire  x661_b330_D48; // @[package.scala 96:25:@44505.4 package.scala 96:25:@44506.4]
  wire  _T_568; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 222:291:@44540.4]
  wire  x662_b331_D48; // @[package.scala 96:25:@44514.4 package.scala 96:25:@44515.4]
  wire [31:0] x664_x351_rdcol_D26_number; // @[package.scala 96:25:@44556.4 package.scala 96:25:@44557.4]
  wire [31:0] _T_579; // @[Math.scala 476:37:@44562.4]
  wire  x370; // @[package.scala 96:25:@44570.4 package.scala 96:25:@44571.4]
  wire  x371; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 230:24:@44574.4]
  wire  _T_608; // @[package.scala 96:25:@44615.4 package.scala 96:25:@44616.4]
  wire  _T_610; // @[implicits.scala 55:10:@44617.4]
  wire  _T_611; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 243:194:@44618.4]
  wire  x665_x372_D20; // @[package.scala 96:25:@44585.4 package.scala 96:25:@44586.4]
  wire  _T_612; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 243:283:@44619.4]
  wire  _T_613; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 243:291:@44620.4]
  wire [31:0] x668_x345_rdcol_D26_number; // @[package.scala 96:25:@44636.4 package.scala 96:25:@44637.4]
  wire [31:0] _T_624; // @[Math.scala 476:37:@44642.4]
  wire  x375; // @[package.scala 96:25:@44650.4 package.scala 96:25:@44651.4]
  wire  x376; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 251:24:@44654.4]
  wire  _T_653; // @[package.scala 96:25:@44695.4 package.scala 96:25:@44696.4]
  wire  _T_655; // @[implicits.scala 55:10:@44697.4]
  wire  _T_656; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 264:194:@44698.4]
  wire  x671_x377_D20; // @[package.scala 96:25:@44683.4 package.scala 96:25:@44684.4]
  wire  _T_657; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 264:283:@44699.4]
  wire  _T_658; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 264:291:@44700.4]
  wire [31:0] x672_b329_D26_number; // @[package.scala 96:25:@44716.4 package.scala 96:25:@44717.4]
  wire [31:0] _T_669; // @[Math.scala 476:37:@44722.4]
  wire  x364; // @[package.scala 96:25:@44431.4 package.scala 96:25:@44432.4]
  wire  x380; // @[package.scala 96:25:@44730.4 package.scala 96:25:@44731.4]
  wire  x381; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 272:24:@44734.4]
  wire  _T_698; // @[package.scala 96:25:@44775.4 package.scala 96:25:@44776.4]
  wire  _T_700; // @[implicits.scala 55:10:@44777.4]
  wire  _T_701; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 285:194:@44778.4]
  wire  x675_x382_D21; // @[package.scala 96:25:@44763.4 package.scala 96:25:@44764.4]
  wire  _T_702; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 285:283:@44779.4]
  wire  _T_703; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 285:291:@44780.4]
  wire [31:0] x385_rdcol_number; // @[Math.scala 154:22:@44799.4 Math.scala 155:14:@44800.4]
  wire [31:0] _T_718; // @[Math.scala 476:37:@44805.4]
  wire  x386; // @[package.scala 96:25:@44813.4 package.scala 96:25:@44814.4]
  wire  x387; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 293:24:@44817.4]
  wire  _T_766; // @[package.scala 96:25:@44894.4 package.scala 96:25:@44895.4]
  wire  _T_768; // @[implicits.scala 55:10:@44896.4]
  wire  _T_769; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 320:194:@44897.4]
  wire  x678_x388_D20; // @[package.scala 96:25:@44882.4 package.scala 96:25:@44883.4]
  wire  _T_770; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 320:283:@44898.4]
  wire  _T_771; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 320:291:@44899.4]
  wire [31:0] x394_rdcol_number; // @[Math.scala 154:22:@44918.4 Math.scala 155:14:@44919.4]
  wire [31:0] _T_786; // @[Math.scala 476:37:@44924.4]
  wire  x395; // @[package.scala 96:25:@44932.4 package.scala 96:25:@44933.4]
  wire  x396; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 328:59:@44936.4]
  wire  _T_829; // @[package.scala 96:25:@45002.4 package.scala 96:25:@45003.4]
  wire  _T_831; // @[implicits.scala 55:10:@45004.4]
  wire  _T_832; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 345:194:@45005.4]
  wire  x679_x397_D20; // @[package.scala 96:25:@44981.4 package.scala 96:25:@44982.4]
  wire  _T_833; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 345:283:@45006.4]
  wire  _T_834; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 345:291:@45007.4]
  wire [31:0] x403_rdrow_number; // @[Math.scala 195:22:@45026.4 Math.scala 196:14:@45027.4]
  wire [31:0] _T_851; // @[Math.scala 406:49:@45033.4]
  wire [31:0] _T_853; // @[Math.scala 406:56:@45035.4]
  wire [31:0] _T_854; // @[Math.scala 406:56:@45036.4]
  wire [31:0] x622_number; // @[implicits.scala 133:21:@45037.4]
  wire  x405; // @[package.scala 96:25:@45051.4 package.scala 96:25:@45052.4]
  wire  x406; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 355:24:@45055.4]
  wire [31:0] _T_877; // @[Math.scala 406:49:@45064.4]
  wire [31:0] _T_879; // @[Math.scala 406:56:@45066.4]
  wire [31:0] _T_880; // @[Math.scala 406:56:@45067.4]
  wire [31:0] _T_884; // @[package.scala 96:25:@45075.4]
  wire  _T_888; // @[FixedPoint.scala 50:25:@45082.4]
  wire [1:0] _T_892; // @[Bitwise.scala 72:12:@45084.4]
  wire [29:0] _T_893; // @[FixedPoint.scala 18:52:@45085.4]
  wire  _T_899; // @[Math.scala 451:55:@45087.4]
  wire [1:0] _T_900; // @[FixedPoint.scala 18:52:@45088.4]
  wire  _T_906; // @[Math.scala 451:110:@45090.4]
  wire  _T_907; // @[Math.scala 451:94:@45091.4]
  wire [31:0] _T_911; // @[package.scala 96:25:@45099.4 package.scala 96:25:@45100.4]
  wire [31:0] x409_1_number; // @[Math.scala 454:20:@45101.4]
  wire [39:0] _GEN_2; // @[Math.scala 461:32:@45106.4]
  wire [39:0] _T_916; // @[Math.scala 461:32:@45106.4]
  wire [37:0] _GEN_3; // @[Math.scala 461:32:@45111.4]
  wire [37:0] _T_919; // @[Math.scala 461:32:@45111.4]
  wire  _T_949; // @[package.scala 96:25:@45179.4 package.scala 96:25:@45180.4]
  wire  _T_951; // @[implicits.scala 55:10:@45181.4]
  wire  _T_952; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 382:194:@45182.4]
  wire  x684_x407_D20; // @[package.scala 96:25:@45167.4 package.scala 96:25:@45168.4]
  wire  _T_953; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 382:283:@45183.4]
  wire  _T_954; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 382:291:@45184.4]
  wire  x414; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 386:24:@45195.4]
  wire  _T_981; // @[package.scala 96:25:@45237.4 package.scala 96:25:@45238.4]
  wire  _T_983; // @[implicits.scala 55:10:@45239.4]
  wire  _T_984; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 399:194:@45240.4]
  wire  x686_x415_D20; // @[package.scala 96:25:@45225.4 package.scala 96:25:@45226.4]
  wire  _T_985; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 399:283:@45241.4]
  wire  _T_986; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 399:291:@45242.4]
  wire  x419; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 403:24:@45253.4]
  wire  _T_1013; // @[package.scala 96:25:@45295.4 package.scala 96:25:@45296.4]
  wire  _T_1015; // @[implicits.scala 55:10:@45297.4]
  wire  _T_1016; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 416:194:@45298.4]
  wire  x688_x420_D20; // @[package.scala 96:25:@45283.4 package.scala 96:25:@45284.4]
  wire  _T_1017; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 416:283:@45299.4]
  wire  _T_1018; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 416:291:@45300.4]
  wire  x689_x380_D1; // @[package.scala 96:25:@45316.4 package.scala 96:25:@45317.4]
  wire  x424; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 428:59:@45320.4]
  wire  _T_1056; // @[package.scala 96:25:@45382.4 package.scala 96:25:@45383.4]
  wire  _T_1058; // @[implicits.scala 55:10:@45384.4]
  wire  _T_1059; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 447:194:@45385.4]
  wire  x692_x425_D20; // @[package.scala 96:25:@45361.4 package.scala 96:25:@45362.4]
  wire  _T_1060; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 447:283:@45386.4]
  wire  _T_1061; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 447:291:@45387.4]
  wire  x429; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 451:59:@45398.4]
  wire  _T_1085; // @[package.scala 96:25:@45431.4 package.scala 96:25:@45432.4]
  wire  _T_1087; // @[implicits.scala 55:10:@45433.4]
  wire  _T_1088; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 462:194:@45434.4]
  wire  x694_x430_D20; // @[package.scala 96:25:@45419.4 package.scala 96:25:@45420.4]
  wire  _T_1089; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 462:283:@45435.4]
  wire  _T_1090; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 462:291:@45436.4]
  wire  x434; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 466:59:@45447.4]
  wire  _T_1114; // @[package.scala 96:25:@45480.4 package.scala 96:25:@45481.4]
  wire  _T_1116; // @[implicits.scala 55:10:@45482.4]
  wire  _T_1117; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 477:194:@45483.4]
  wire  x695_x435_D20; // @[package.scala 96:25:@45468.4 package.scala 96:25:@45469.4]
  wire  _T_1118; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 477:283:@45484.4]
  wire  _T_1119; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 477:291:@45485.4]
  wire [31:0] x439_rdrow_number; // @[Math.scala 195:22:@45504.4 Math.scala 196:14:@45505.4]
  wire [31:0] _T_1136; // @[Math.scala 406:49:@45511.4]
  wire [31:0] _T_1138; // @[Math.scala 406:56:@45513.4]
  wire [31:0] _T_1139; // @[Math.scala 406:56:@45514.4]
  wire [31:0] x627_number; // @[implicits.scala 133:21:@45515.4]
  wire  x441; // @[package.scala 96:25:@45529.4 package.scala 96:25:@45530.4]
  wire  x442; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 487:24:@45533.4]
  wire [31:0] _T_1162; // @[Math.scala 406:49:@45542.4]
  wire [31:0] _T_1164; // @[Math.scala 406:56:@45544.4]
  wire [31:0] _T_1165; // @[Math.scala 406:56:@45545.4]
  wire [31:0] _T_1169; // @[package.scala 96:25:@45553.4]
  wire  _T_1173; // @[FixedPoint.scala 50:25:@45560.4]
  wire [1:0] _T_1177; // @[Bitwise.scala 72:12:@45562.4]
  wire [29:0] _T_1178; // @[FixedPoint.scala 18:52:@45563.4]
  wire  _T_1184; // @[Math.scala 451:55:@45565.4]
  wire [1:0] _T_1185; // @[FixedPoint.scala 18:52:@45566.4]
  wire  _T_1191; // @[Math.scala 451:110:@45568.4]
  wire  _T_1192; // @[Math.scala 451:94:@45569.4]
  wire [31:0] _T_1196; // @[package.scala 96:25:@45577.4 package.scala 96:25:@45578.4]
  wire [31:0] x445_1_number; // @[Math.scala 454:20:@45579.4]
  wire [39:0] _GEN_4; // @[Math.scala 461:32:@45584.4]
  wire [39:0] _T_1201; // @[Math.scala 461:32:@45584.4]
  wire [37:0] _GEN_5; // @[Math.scala 461:32:@45589.4]
  wire [37:0] _T_1204; // @[Math.scala 461:32:@45589.4]
  wire  _T_1231; // @[package.scala 96:25:@45648.4 package.scala 96:25:@45649.4]
  wire  _T_1233; // @[implicits.scala 55:10:@45650.4]
  wire  _T_1234; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 512:194:@45651.4]
  wire  x698_x443_D20; // @[package.scala 96:25:@45636.4 package.scala 96:25:@45637.4]
  wire  _T_1235; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 512:283:@45652.4]
  wire  _T_1236; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 512:291:@45653.4]
  wire  x450; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 516:24:@45664.4]
  wire  _T_1260; // @[package.scala 96:25:@45697.4 package.scala 96:25:@45698.4]
  wire  _T_1262; // @[implicits.scala 55:10:@45699.4]
  wire  _T_1263; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 527:194:@45700.4]
  wire  x699_x451_D20; // @[package.scala 96:25:@45685.4 package.scala 96:25:@45686.4]
  wire  _T_1264; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 527:283:@45701.4]
  wire  _T_1265; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 527:291:@45702.4]
  wire  x455; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 531:24:@45713.4]
  wire  _T_1289; // @[package.scala 96:25:@45746.4 package.scala 96:25:@45747.4]
  wire  _T_1291; // @[implicits.scala 55:10:@45748.4]
  wire  _T_1292; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 548:194:@45749.4]
  wire  x700_x456_D20; // @[package.scala 96:25:@45734.4 package.scala 96:25:@45735.4]
  wire  _T_1293; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 548:283:@45750.4]
  wire  _T_1294; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 548:326:@45751.4]
  wire  x460; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 552:59:@45762.4]
  wire  _T_1326; // @[package.scala 96:25:@45815.4 package.scala 96:25:@45816.4]
  wire  _T_1328; // @[implicits.scala 55:10:@45817.4]
  wire  _T_1329; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 569:194:@45818.4]
  wire  x702_x461_D20; // @[package.scala 96:25:@45794.4 package.scala 96:25:@45795.4]
  wire  _T_1330; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 569:283:@45819.4]
  wire  _T_1331; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 569:291:@45820.4]
  wire  x465; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 573:59:@45831.4]
  wire  _T_1355; // @[package.scala 96:25:@45864.4 package.scala 96:25:@45865.4]
  wire  _T_1357; // @[implicits.scala 55:10:@45866.4]
  wire  _T_1358; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 584:194:@45867.4]
  wire  x704_x466_D20; // @[package.scala 96:25:@45852.4 package.scala 96:25:@45853.4]
  wire  _T_1359; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 584:283:@45868.4]
  wire  _T_1360; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 584:291:@45869.4]
  wire  x470; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 588:59:@45880.4]
  wire  _T_1384; // @[package.scala 96:25:@45913.4 package.scala 96:25:@45914.4]
  wire  _T_1386; // @[implicits.scala 55:10:@45915.4]
  wire  _T_1387; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 599:194:@45916.4]
  wire  x705_x471_D20; // @[package.scala 96:25:@45901.4 package.scala 96:25:@45902.4]
  wire  _T_1388; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 599:283:@45917.4]
  wire  _T_1389; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 599:291:@45918.4]
  wire [31:0] x531_number; // @[Math.scala 723:22:@46572.4 Math.scala 724:14:@46573.4]
  wire [31:0] x548_number; // @[Math.scala 723:22:@46765.4 Math.scala 724:14:@46766.4]
  wire [63:0] _T_1777; // @[Cat.scala 30:58:@46774.4]
  wire [31:0] x494_number; // @[Math.scala 723:22:@46152.4 Math.scala 724:14:@46153.4]
  wire [31:0] x514_number; // @[Math.scala 723:22:@46381.4 Math.scala 724:14:@46382.4]
  wire [63:0] _T_1778; // @[Cat.scala 30:58:@46775.4]
  wire  _T_1791; // @[package.scala 96:25:@46811.4 package.scala 96:25:@46812.4]
  wire  _T_1793; // @[implicits.scala 55:10:@46813.4]
  wire  x711_b330_D69; // @[package.scala 96:25:@46802.4 package.scala 96:25:@46803.4]
  wire  _T_1794; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 783:117:@46814.4]
  wire  x710_b331_D69; // @[package.scala 96:25:@46793.4 package.scala 96:25:@46794.4]
  wire  _T_1795; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 783:123:@46815.4]
  wire [31:0] x639_x339_D8_number; // @[package.scala 96:25:@44035.4 package.scala 96:25:@44036.4]
  wire [31:0] x640_x343_sum_D3_number; // @[package.scala 96:25:@44044.4 package.scala 96:25:@44045.4]
  wire [31:0] x641_x618_D24_number; // @[package.scala 96:25:@44053.4 package.scala 96:25:@44054.4]
  wire [31:0] x646_x347_D7_number; // @[package.scala 96:25:@44169.4 package.scala 96:25:@44170.4]
  wire [31:0] x647_x349_sum_D2_number; // @[package.scala 96:25:@44178.4 package.scala 96:25:@44179.4]
  wire [31:0] x650_x353_D7_number; // @[package.scala 96:25:@44276.4 package.scala 96:25:@44277.4]
  wire [31:0] x651_x355_sum_D2_number; // @[package.scala 96:25:@44285.4 package.scala 96:25:@44286.4]
  wire [31:0] x652_x361_sum_D2_number; // @[package.scala 96:25:@44365.4 package.scala 96:25:@44366.4]
  wire [31:0] x653_x359_D7_number; // @[package.scala 96:25:@44374.4 package.scala 96:25:@44375.4]
  wire [31:0] x658_x361_sum_D26_number; // @[package.scala 96:25:@44478.4 package.scala 96:25:@44479.4]
  wire [31:0] x659_x618_D48_number; // @[package.scala 96:25:@44487.4 package.scala 96:25:@44488.4]
  wire [31:0] x663_x359_D31_number; // @[package.scala 96:25:@44523.4 package.scala 96:25:@44524.4]
  wire [31:0] x666_x353_D31_number; // @[package.scala 96:25:@44594.4 package.scala 96:25:@44595.4]
  wire [31:0] x667_x355_sum_D26_number; // @[package.scala 96:25:@44603.4 package.scala 96:25:@44604.4]
  wire [31:0] x669_x347_D31_number; // @[package.scala 96:25:@44665.4 package.scala 96:25:@44666.4]
  wire [31:0] x670_x349_sum_D26_number; // @[package.scala 96:25:@44674.4 package.scala 96:25:@44675.4]
  wire [31:0] x673_x339_D32_number; // @[package.scala 96:25:@44745.4 package.scala 96:25:@44746.4]
  wire [31:0] x674_x343_sum_D27_number; // @[package.scala 96:25:@44754.4 package.scala 96:25:@44755.4]
  wire [31:0] x391_sum_number; // @[Math.scala 154:22:@44864.4 Math.scala 155:14:@44865.4]
  wire [31:0] x677_x389_D5_number; // @[package.scala 96:25:@44873.4 package.scala 96:25:@44874.4]
  wire [31:0] x400_sum_number; // @[Math.scala 154:22:@44972.4 Math.scala 155:14:@44973.4]
  wire [31:0] x680_x398_D5_number; // @[package.scala 96:25:@44990.4 package.scala 96:25:@44991.4]
  wire [31:0] x411_sum_number; // @[Math.scala 154:22:@45149.4 Math.scala 155:14:@45150.4]
  wire [31:0] x683_x623_D20_number; // @[package.scala 96:25:@45158.4 package.scala 96:25:@45159.4]
  wire [31:0] x416_sum_number; // @[Math.scala 154:22:@45216.4 Math.scala 155:14:@45217.4]
  wire [31:0] x421_sum_number; // @[Math.scala 154:22:@45274.4 Math.scala 155:14:@45275.4]
  wire [31:0] x693_x426_sum_D1_number; // @[package.scala 96:25:@45370.4 package.scala 96:25:@45371.4]
  wire [31:0] x431_sum_number; // @[Math.scala 154:22:@45410.4 Math.scala 155:14:@45411.4]
  wire [31:0] x436_sum_number; // @[Math.scala 154:22:@45459.4 Math.scala 155:14:@45460.4]
  wire [31:0] x447_sum_number; // @[Math.scala 154:22:@45618.4 Math.scala 155:14:@45619.4]
  wire [31:0] x697_x628_D20_number; // @[package.scala 96:25:@45627.4 package.scala 96:25:@45628.4]
  wire [31:0] x452_sum_number; // @[Math.scala 154:22:@45676.4 Math.scala 155:14:@45677.4]
  wire [31:0] x457_sum_number; // @[Math.scala 154:22:@45725.4 Math.scala 155:14:@45726.4]
  wire [31:0] x703_x462_sum_D1_number; // @[package.scala 96:25:@45803.4 package.scala 96:25:@45804.4]
  wire [31:0] x467_sum_number; // @[Math.scala 154:22:@45843.4 Math.scala 155:14:@45844.4]
  wire [31:0] x472_sum_number; // @[Math.scala 154:22:@45892.4 Math.scala 155:14:@45893.4]
  _ _ ( // @[Math.scala 720:24:@43724.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@43736.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_56 RetimeWrapper ( // @[package.scala 93:22:@43759.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x334_lb_0 x334_lb_0 ( // @[m_x334_lb_0.scala 47:17:@43769.4]
    .clock(x334_lb_0_clock),
    .reset(x334_lb_0_reset),
    .io_rPort_17_banks_1(x334_lb_0_io_rPort_17_banks_1),
    .io_rPort_17_banks_0(x334_lb_0_io_rPort_17_banks_0),
    .io_rPort_17_ofs_0(x334_lb_0_io_rPort_17_ofs_0),
    .io_rPort_17_en_0(x334_lb_0_io_rPort_17_en_0),
    .io_rPort_17_backpressure(x334_lb_0_io_rPort_17_backpressure),
    .io_rPort_17_output_0(x334_lb_0_io_rPort_17_output_0),
    .io_rPort_16_banks_1(x334_lb_0_io_rPort_16_banks_1),
    .io_rPort_16_banks_0(x334_lb_0_io_rPort_16_banks_0),
    .io_rPort_16_ofs_0(x334_lb_0_io_rPort_16_ofs_0),
    .io_rPort_16_en_0(x334_lb_0_io_rPort_16_en_0),
    .io_rPort_16_backpressure(x334_lb_0_io_rPort_16_backpressure),
    .io_rPort_16_output_0(x334_lb_0_io_rPort_16_output_0),
    .io_rPort_15_banks_1(x334_lb_0_io_rPort_15_banks_1),
    .io_rPort_15_banks_0(x334_lb_0_io_rPort_15_banks_0),
    .io_rPort_15_ofs_0(x334_lb_0_io_rPort_15_ofs_0),
    .io_rPort_15_en_0(x334_lb_0_io_rPort_15_en_0),
    .io_rPort_15_backpressure(x334_lb_0_io_rPort_15_backpressure),
    .io_rPort_15_output_0(x334_lb_0_io_rPort_15_output_0),
    .io_rPort_14_banks_1(x334_lb_0_io_rPort_14_banks_1),
    .io_rPort_14_banks_0(x334_lb_0_io_rPort_14_banks_0),
    .io_rPort_14_ofs_0(x334_lb_0_io_rPort_14_ofs_0),
    .io_rPort_14_en_0(x334_lb_0_io_rPort_14_en_0),
    .io_rPort_14_backpressure(x334_lb_0_io_rPort_14_backpressure),
    .io_rPort_14_output_0(x334_lb_0_io_rPort_14_output_0),
    .io_rPort_13_banks_1(x334_lb_0_io_rPort_13_banks_1),
    .io_rPort_13_banks_0(x334_lb_0_io_rPort_13_banks_0),
    .io_rPort_13_ofs_0(x334_lb_0_io_rPort_13_ofs_0),
    .io_rPort_13_en_0(x334_lb_0_io_rPort_13_en_0),
    .io_rPort_13_backpressure(x334_lb_0_io_rPort_13_backpressure),
    .io_rPort_13_output_0(x334_lb_0_io_rPort_13_output_0),
    .io_rPort_12_banks_1(x334_lb_0_io_rPort_12_banks_1),
    .io_rPort_12_banks_0(x334_lb_0_io_rPort_12_banks_0),
    .io_rPort_12_ofs_0(x334_lb_0_io_rPort_12_ofs_0),
    .io_rPort_12_en_0(x334_lb_0_io_rPort_12_en_0),
    .io_rPort_12_backpressure(x334_lb_0_io_rPort_12_backpressure),
    .io_rPort_12_output_0(x334_lb_0_io_rPort_12_output_0),
    .io_rPort_11_banks_1(x334_lb_0_io_rPort_11_banks_1),
    .io_rPort_11_banks_0(x334_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x334_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x334_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x334_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x334_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_1(x334_lb_0_io_rPort_10_banks_1),
    .io_rPort_10_banks_0(x334_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x334_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x334_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x334_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x334_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_1(x334_lb_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x334_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x334_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x334_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x334_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x334_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x334_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x334_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x334_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x334_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x334_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x334_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x334_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x334_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x334_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x334_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x334_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x334_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x334_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x334_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x334_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x334_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x334_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x334_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x334_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x334_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x334_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x334_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x334_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x334_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x334_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x334_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x334_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x334_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x334_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x334_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x334_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x334_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x334_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x334_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x334_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x334_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x334_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x334_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x334_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x334_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x334_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x334_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x334_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x334_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x334_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x334_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x334_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x334_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x334_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x334_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x334_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x334_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x334_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x334_lb_0_io_rPort_0_output_0),
    .io_wPort_3_banks_1(x334_lb_0_io_wPort_3_banks_1),
    .io_wPort_3_banks_0(x334_lb_0_io_wPort_3_banks_0),
    .io_wPort_3_ofs_0(x334_lb_0_io_wPort_3_ofs_0),
    .io_wPort_3_data_0(x334_lb_0_io_wPort_3_data_0),
    .io_wPort_3_en_0(x334_lb_0_io_wPort_3_en_0),
    .io_wPort_2_banks_1(x334_lb_0_io_wPort_2_banks_1),
    .io_wPort_2_banks_0(x334_lb_0_io_wPort_2_banks_0),
    .io_wPort_2_ofs_0(x334_lb_0_io_wPort_2_ofs_0),
    .io_wPort_2_data_0(x334_lb_0_io_wPort_2_data_0),
    .io_wPort_2_en_0(x334_lb_0_io_wPort_2_en_0),
    .io_wPort_1_banks_1(x334_lb_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x334_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x334_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x334_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x334_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x334_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x334_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x334_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x334_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x334_lb_0_io_wPort_0_en_0)
  );
  x339 x339_1 ( // @[Math.scala 366:24:@43952.4]
    .clock(x339_1_clock),
    .io_a(x339_1_io_a),
    .io_flow(x339_1_io_flow),
    .io_result(x339_1_io_result)
  );
  x303_sum x621_sum_1 ( // @[Math.scala 150:24:@43989.4]
    .clock(x621_sum_1_clock),
    .reset(x621_sum_1_reset),
    .io_a(x621_sum_1_io_a),
    .io_b(x621_sum_1_io_b),
    .io_flow(x621_sum_1_io_flow),
    .io_result(x621_sum_1_io_result)
  );
  x342_div x342_div_1 ( // @[Math.scala 327:24:@44001.4]
    .clock(x342_div_1_clock),
    .io_a(x342_div_1_io_a),
    .io_flow(x342_div_1_io_flow),
    .io_result(x342_div_1_io_result)
  );
  RetimeWrapper_298 RetimeWrapper_1 ( // @[package.scala 93:22:@44011.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x303_sum x343_sum_1 ( // @[Math.scala 150:24:@44020.4]
    .clock(x343_sum_1_clock),
    .reset(x343_sum_1_reset),
    .io_a(x343_sum_1_io_a),
    .io_b(x343_sum_1_io_b),
    .io_flow(x343_sum_1_io_flow),
    .io_result(x343_sum_1_io_result)
  );
  RetimeWrapper_300 RetimeWrapper_2 ( // @[package.scala 93:22:@44030.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_301 RetimeWrapper_3 ( // @[package.scala 93:22:@44039.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_302 RetimeWrapper_4 ( // @[package.scala 93:22:@44048.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_303 RetimeWrapper_5 ( // @[package.scala 93:22:@44057.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_303 RetimeWrapper_6 ( // @[package.scala 93:22:@44066.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_305 RetimeWrapper_7 ( // @[package.scala 93:22:@44075.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_303 RetimeWrapper_8 ( // @[package.scala 93:22:@44086.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  x303_sum x345_rdcol_1 ( // @[Math.scala 150:24:@44109.4]
    .clock(x345_rdcol_1_clock),
    .reset(x345_rdcol_1_reset),
    .io_a(x345_rdcol_1_io_a),
    .io_b(x345_rdcol_1_io_b),
    .io_flow(x345_rdcol_1_io_flow),
    .io_result(x345_rdcol_1_io_result)
  );
  x339 x347_1 ( // @[Math.scala 366:24:@44123.4]
    .clock(x347_1_clock),
    .io_a(x347_1_io_a),
    .io_flow(x347_1_io_flow),
    .io_result(x347_1_io_result)
  );
  x342_div x348_div_1 ( // @[Math.scala 327:24:@44135.4]
    .clock(x348_div_1_clock),
    .io_a(x348_div_1_io_a),
    .io_flow(x348_div_1_io_flow),
    .io_result(x348_div_1_io_result)
  );
  RetimeWrapper_308 RetimeWrapper_9 ( // @[package.scala 93:22:@44145.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  x303_sum x349_sum_1 ( // @[Math.scala 150:24:@44154.4]
    .clock(x349_sum_1_clock),
    .reset(x349_sum_1_reset),
    .io_a(x349_sum_1_io_a),
    .io_b(x349_sum_1_io_b),
    .io_flow(x349_sum_1_io_flow),
    .io_result(x349_sum_1_io_result)
  );
  RetimeWrapper_310 RetimeWrapper_10 ( // @[package.scala 93:22:@44164.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_11 ( // @[package.scala 93:22:@44173.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_305 RetimeWrapper_12 ( // @[package.scala 93:22:@44182.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_303 RetimeWrapper_13 ( // @[package.scala 93:22:@44193.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  x303_sum x351_rdcol_1 ( // @[Math.scala 150:24:@44216.4]
    .clock(x351_rdcol_1_clock),
    .reset(x351_rdcol_1_reset),
    .io_a(x351_rdcol_1_io_a),
    .io_b(x351_rdcol_1_io_b),
    .io_flow(x351_rdcol_1_io_flow),
    .io_result(x351_rdcol_1_io_result)
  );
  x339 x353_1 ( // @[Math.scala 366:24:@44230.4]
    .clock(x353_1_clock),
    .io_a(x353_1_io_a),
    .io_flow(x353_1_io_flow),
    .io_result(x353_1_io_result)
  );
  x342_div x354_div_1 ( // @[Math.scala 327:24:@44242.4]
    .clock(x354_div_1_clock),
    .io_a(x354_div_1_io_a),
    .io_flow(x354_div_1_io_flow),
    .io_result(x354_div_1_io_result)
  );
  x303_sum x355_sum_1 ( // @[Math.scala 150:24:@44252.4]
    .clock(x355_sum_1_clock),
    .reset(x355_sum_1_reset),
    .io_a(x355_sum_1_io_a),
    .io_b(x355_sum_1_io_b),
    .io_flow(x355_sum_1_io_flow),
    .io_result(x355_sum_1_io_result)
  );
  RetimeWrapper_305 RetimeWrapper_14 ( // @[package.scala 93:22:@44262.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_310 RetimeWrapper_15 ( // @[package.scala 93:22:@44271.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_311 RetimeWrapper_16 ( // @[package.scala 93:22:@44280.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_303 RetimeWrapper_17 ( // @[package.scala 93:22:@44291.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  x303_sum x357_rdcol_1 ( // @[Math.scala 150:24:@44314.4]
    .clock(x357_rdcol_1_clock),
    .reset(x357_rdcol_1_reset),
    .io_a(x357_rdcol_1_io_a),
    .io_b(x357_rdcol_1_io_b),
    .io_flow(x357_rdcol_1_io_flow),
    .io_result(x357_rdcol_1_io_result)
  );
  x339 x359_1 ( // @[Math.scala 366:24:@44328.4]
    .clock(x359_1_clock),
    .io_a(x359_1_io_a),
    .io_flow(x359_1_io_flow),
    .io_result(x359_1_io_result)
  );
  x342_div x360_div_1 ( // @[Math.scala 327:24:@44340.4]
    .clock(x360_div_1_clock),
    .io_a(x360_div_1_io_a),
    .io_flow(x360_div_1_io_flow),
    .io_result(x360_div_1_io_result)
  );
  x303_sum x361_sum_1 ( // @[Math.scala 150:24:@44350.4]
    .clock(x361_sum_1_clock),
    .reset(x361_sum_1_reset),
    .io_a(x361_sum_1_io_a),
    .io_b(x361_sum_1_io_b),
    .io_flow(x361_sum_1_io_flow),
    .io_result(x361_sum_1_io_result)
  );
  RetimeWrapper_311 RetimeWrapper_18 ( // @[package.scala 93:22:@44360.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_310 RetimeWrapper_19 ( // @[package.scala 93:22:@44369.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_305 RetimeWrapper_20 ( // @[package.scala 93:22:@44378.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_303 RetimeWrapper_21 ( // @[package.scala 93:22:@44389.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_22 ( // @[package.scala 93:22:@44410.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper RetimeWrapper_23 ( // @[package.scala 93:22:@44426.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_24 ( // @[package.scala 93:22:@44435.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@44449.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper RetimeWrapper_26 ( // @[package.scala 93:22:@44458.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_27 ( // @[package.scala 93:22:@44473.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_332 RetimeWrapper_28 ( // @[package.scala 93:22:@44482.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_29 ( // @[package.scala 93:22:@44491.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_30 ( // @[package.scala 93:22:@44500.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_31 ( // @[package.scala 93:22:@44509.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_336 RetimeWrapper_32 ( // @[package.scala 93:22:@44518.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_33 ( // @[package.scala 93:22:@44530.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_34 ( // @[package.scala 93:22:@44551.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper RetimeWrapper_35 ( // @[package.scala 93:22:@44565.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_36 ( // @[package.scala 93:22:@44580.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_336 RetimeWrapper_37 ( // @[package.scala 93:22:@44589.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_38 ( // @[package.scala 93:22:@44598.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_39 ( // @[package.scala 93:22:@44610.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_40 ( // @[package.scala 93:22:@44631.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper RetimeWrapper_41 ( // @[package.scala 93:22:@44645.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_336 RetimeWrapper_42 ( // @[package.scala 93:22:@44660.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_43 ( // @[package.scala 93:22:@44669.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_44 ( // @[package.scala 93:22:@44678.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_45 ( // @[package.scala 93:22:@44690.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_46 ( // @[package.scala 93:22:@44711.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper RetimeWrapper_47 ( // @[package.scala 93:22:@44725.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_352 RetimeWrapper_48 ( // @[package.scala 93:22:@44740.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_353 RetimeWrapper_49 ( // @[package.scala 93:22:@44749.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_354 RetimeWrapper_50 ( // @[package.scala 93:22:@44758.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_51 ( // @[package.scala 93:22:@44770.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  x303_sum x385_rdcol_1 ( // @[Math.scala 150:24:@44793.4]
    .clock(x385_rdcol_1_clock),
    .reset(x385_rdcol_1_reset),
    .io_a(x385_rdcol_1_io_a),
    .io_b(x385_rdcol_1_io_b),
    .io_flow(x385_rdcol_1_io_flow),
    .io_result(x385_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_52 ( // @[package.scala 93:22:@44808.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  x339 x389_1 ( // @[Math.scala 366:24:@44827.4]
    .clock(x389_1_clock),
    .io_a(x389_1_io_a),
    .io_flow(x389_1_io_flow),
    .io_result(x389_1_io_result)
  );
  x342_div x390_div_1 ( // @[Math.scala 327:24:@44839.4]
    .clock(x390_div_1_clock),
    .io_a(x390_div_1_io_a),
    .io_flow(x390_div_1_io_flow),
    .io_result(x390_div_1_io_result)
  );
  RetimeWrapper_358 RetimeWrapper_53 ( // @[package.scala 93:22:@44849.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  x303_sum x391_sum_1 ( // @[Math.scala 150:24:@44858.4]
    .clock(x391_sum_1_clock),
    .reset(x391_sum_1_reset),
    .io_a(x391_sum_1_io_a),
    .io_b(x391_sum_1_io_b),
    .io_flow(x391_sum_1_io_flow),
    .io_result(x391_sum_1_io_result)
  );
  RetimeWrapper_360 RetimeWrapper_54 ( // @[package.scala 93:22:@44868.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_55 ( // @[package.scala 93:22:@44877.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_56 ( // @[package.scala 93:22:@44889.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  x303_sum x394_rdcol_1 ( // @[Math.scala 150:24:@44912.4]
    .clock(x394_rdcol_1_clock),
    .reset(x394_rdcol_1_reset),
    .io_a(x394_rdcol_1_io_a),
    .io_b(x394_rdcol_1_io_b),
    .io_flow(x394_rdcol_1_io_flow),
    .io_result(x394_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_57 ( // @[package.scala 93:22:@44927.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  x339 x398_1 ( // @[Math.scala 366:24:@44944.4]
    .clock(x398_1_clock),
    .io_a(x398_1_io_a),
    .io_flow(x398_1_io_flow),
    .io_result(x398_1_io_result)
  );
  x342_div x399_div_1 ( // @[Math.scala 327:24:@44956.4]
    .clock(x399_div_1_clock),
    .io_a(x399_div_1_io_a),
    .io_flow(x399_div_1_io_flow),
    .io_result(x399_div_1_io_result)
  );
  x303_sum x400_sum_1 ( // @[Math.scala 150:24:@44966.4]
    .clock(x400_sum_1_clock),
    .reset(x400_sum_1_reset),
    .io_a(x400_sum_1_io_a),
    .io_b(x400_sum_1_io_b),
    .io_flow(x400_sum_1_io_flow),
    .io_result(x400_sum_1_io_result)
  );
  RetimeWrapper_333 RetimeWrapper_58 ( // @[package.scala 93:22:@44976.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_360 RetimeWrapper_59 ( // @[package.scala 93:22:@44985.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_60 ( // @[package.scala 93:22:@44997.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  x604_sub x403_rdrow_1 ( // @[Math.scala 191:24:@45020.4]
    .clock(x403_rdrow_1_clock),
    .reset(x403_rdrow_1_reset),
    .io_a(x403_rdrow_1_io_a),
    .io_b(x403_rdrow_1_io_b),
    .io_flow(x403_rdrow_1_io_flow),
    .io_result(x403_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_61 ( // @[package.scala 93:22:@45046.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_62 ( // @[package.scala 93:22:@45068.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_63 ( // @[package.scala 93:22:@45094.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  x303_sum x626_sum_1 ( // @[Math.scala 150:24:@45115.4]
    .clock(x626_sum_1_clock),
    .reset(x626_sum_1_reset),
    .io_a(x626_sum_1_io_a),
    .io_b(x626_sum_1_io_b),
    .io_flow(x626_sum_1_io_flow),
    .io_result(x626_sum_1_io_result)
  );
  RetimeWrapper_374 RetimeWrapper_64 ( // @[package.scala 93:22:@45125.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_65 ( // @[package.scala 93:22:@45134.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  x303_sum x411_sum_1 ( // @[Math.scala 150:24:@45143.4]
    .clock(x411_sum_1_clock),
    .reset(x411_sum_1_reset),
    .io_a(x411_sum_1_io_a),
    .io_b(x411_sum_1_io_b),
    .io_flow(x411_sum_1_io_flow),
    .io_result(x411_sum_1_io_result)
  );
  RetimeWrapper_308 RetimeWrapper_66 ( // @[package.scala 93:22:@45153.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_67 ( // @[package.scala 93:22:@45162.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_68 ( // @[package.scala 93:22:@45174.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_69 ( // @[package.scala 93:22:@45201.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  x303_sum x416_sum_1 ( // @[Math.scala 150:24:@45210.4]
    .clock(x416_sum_1_clock),
    .reset(x416_sum_1_reset),
    .io_a(x416_sum_1_io_a),
    .io_b(x416_sum_1_io_b),
    .io_flow(x416_sum_1_io_flow),
    .io_result(x416_sum_1_io_result)
  );
  RetimeWrapper_333 RetimeWrapper_70 ( // @[package.scala 93:22:@45220.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_71 ( // @[package.scala 93:22:@45232.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_72 ( // @[package.scala 93:22:@45259.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  x303_sum x421_sum_1 ( // @[Math.scala 150:24:@45268.4]
    .clock(x421_sum_1_clock),
    .reset(x421_sum_1_reset),
    .io_a(x421_sum_1_io_a),
    .io_b(x421_sum_1_io_b),
    .io_flow(x421_sum_1_io_flow),
    .io_result(x421_sum_1_io_result)
  );
  RetimeWrapper_333 RetimeWrapper_73 ( // @[package.scala 93:22:@45278.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_74 ( // @[package.scala 93:22:@45290.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper RetimeWrapper_75 ( // @[package.scala 93:22:@45311.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_76 ( // @[package.scala 93:22:@45326.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_390 RetimeWrapper_77 ( // @[package.scala 93:22:@45335.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  x303_sum x426_sum_1 ( // @[Math.scala 150:24:@45346.4]
    .clock(x426_sum_1_clock),
    .reset(x426_sum_1_reset),
    .io_a(x426_sum_1_io_a),
    .io_b(x426_sum_1_io_b),
    .io_flow(x426_sum_1_io_flow),
    .io_result(x426_sum_1_io_result)
  );
  RetimeWrapper_333 RetimeWrapper_78 ( // @[package.scala 93:22:@45356.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_79 ( // @[package.scala 93:22:@45365.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_80 ( // @[package.scala 93:22:@45377.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  x303_sum x431_sum_1 ( // @[Math.scala 150:24:@45404.4]
    .clock(x431_sum_1_clock),
    .reset(x431_sum_1_reset),
    .io_a(x431_sum_1_io_a),
    .io_b(x431_sum_1_io_b),
    .io_flow(x431_sum_1_io_flow),
    .io_result(x431_sum_1_io_result)
  );
  RetimeWrapper_333 RetimeWrapper_81 ( // @[package.scala 93:22:@45414.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_82 ( // @[package.scala 93:22:@45426.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  x303_sum x436_sum_1 ( // @[Math.scala 150:24:@45453.4]
    .clock(x436_sum_1_clock),
    .reset(x436_sum_1_reset),
    .io_a(x436_sum_1_io_a),
    .io_b(x436_sum_1_io_b),
    .io_flow(x436_sum_1_io_flow),
    .io_result(x436_sum_1_io_result)
  );
  RetimeWrapper_333 RetimeWrapper_83 ( // @[package.scala 93:22:@45463.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_84 ( // @[package.scala 93:22:@45475.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  x604_sub x439_rdrow_1 ( // @[Math.scala 191:24:@45498.4]
    .clock(x439_rdrow_1_clock),
    .reset(x439_rdrow_1_reset),
    .io_a(x439_rdrow_1_io_a),
    .io_b(x439_rdrow_1_io_b),
    .io_flow(x439_rdrow_1_io_flow),
    .io_result(x439_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_85 ( // @[package.scala 93:22:@45524.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_86 ( // @[package.scala 93:22:@45546.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_87 ( // @[package.scala 93:22:@45572.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  x303_sum x631_sum_1 ( // @[Math.scala 150:24:@45593.4]
    .clock(x631_sum_1_clock),
    .reset(x631_sum_1_reset),
    .io_a(x631_sum_1_io_a),
    .io_b(x631_sum_1_io_b),
    .io_flow(x631_sum_1_io_flow),
    .io_result(x631_sum_1_io_result)
  );
  RetimeWrapper_374 RetimeWrapper_88 ( // @[package.scala 93:22:@45603.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  x303_sum x447_sum_1 ( // @[Math.scala 150:24:@45612.4]
    .clock(x447_sum_1_clock),
    .reset(x447_sum_1_reset),
    .io_a(x447_sum_1_io_a),
    .io_b(x447_sum_1_io_b),
    .io_flow(x447_sum_1_io_flow),
    .io_result(x447_sum_1_io_result)
  );
  RetimeWrapper_308 RetimeWrapper_89 ( // @[package.scala 93:22:@45622.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_90 ( // @[package.scala 93:22:@45631.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_91 ( // @[package.scala 93:22:@45643.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  x303_sum x452_sum_1 ( // @[Math.scala 150:24:@45670.4]
    .clock(x452_sum_1_clock),
    .reset(x452_sum_1_reset),
    .io_a(x452_sum_1_io_a),
    .io_b(x452_sum_1_io_b),
    .io_flow(x452_sum_1_io_flow),
    .io_result(x452_sum_1_io_result)
  );
  RetimeWrapper_333 RetimeWrapper_92 ( // @[package.scala 93:22:@45680.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_93 ( // @[package.scala 93:22:@45692.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  x303_sum x457_sum_1 ( // @[Math.scala 150:24:@45719.4]
    .clock(x457_sum_1_clock),
    .reset(x457_sum_1_reset),
    .io_a(x457_sum_1_io_a),
    .io_b(x457_sum_1_io_b),
    .io_flow(x457_sum_1_io_flow),
    .io_result(x457_sum_1_io_result)
  );
  RetimeWrapper_333 RetimeWrapper_94 ( // @[package.scala 93:22:@45729.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_95 ( // @[package.scala 93:22:@45741.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_390 RetimeWrapper_96 ( // @[package.scala 93:22:@45768.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  x303_sum x462_sum_1 ( // @[Math.scala 150:24:@45779.4]
    .clock(x462_sum_1_clock),
    .reset(x462_sum_1_reset),
    .io_a(x462_sum_1_io_a),
    .io_b(x462_sum_1_io_b),
    .io_flow(x462_sum_1_io_flow),
    .io_result(x462_sum_1_io_result)
  );
  RetimeWrapper_333 RetimeWrapper_97 ( // @[package.scala 93:22:@45789.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_98 ( // @[package.scala 93:22:@45798.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_99 ( // @[package.scala 93:22:@45810.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  x303_sum x467_sum_1 ( // @[Math.scala 150:24:@45837.4]
    .clock(x467_sum_1_clock),
    .reset(x467_sum_1_reset),
    .io_a(x467_sum_1_io_a),
    .io_b(x467_sum_1_io_b),
    .io_flow(x467_sum_1_io_flow),
    .io_result(x467_sum_1_io_result)
  );
  RetimeWrapper_333 RetimeWrapper_100 ( // @[package.scala 93:22:@45847.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_101 ( // @[package.scala 93:22:@45859.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  x303_sum x472_sum_1 ( // @[Math.scala 150:24:@45886.4]
    .clock(x472_sum_1_clock),
    .reset(x472_sum_1_reset),
    .io_a(x472_sum_1_io_a),
    .io_b(x472_sum_1_io_b),
    .io_flow(x472_sum_1_io_flow),
    .io_result(x472_sum_1_io_result)
  );
  RetimeWrapper_333 RetimeWrapper_102 ( // @[package.scala 93:22:@45896.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_334 RetimeWrapper_103 ( // @[package.scala 93:22:@45908.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  x475 x475_1 ( // @[Math.scala 262:24:@45931.4]
    .clock(x475_1_clock),
    .io_a(x475_1_io_a),
    .io_b(x475_1_io_b),
    .io_flow(x475_1_io_flow),
    .io_result(x475_1_io_result)
  );
  x475 x476_1 ( // @[Math.scala 262:24:@45943.4]
    .clock(x476_1_clock),
    .io_a(x476_1_io_a),
    .io_b(x476_1_io_b),
    .io_flow(x476_1_io_flow),
    .io_result(x476_1_io_result)
  );
  x475 x477_1 ( // @[Math.scala 262:24:@45955.4]
    .clock(x477_1_clock),
    .io_a(x477_1_io_a),
    .io_b(x477_1_io_b),
    .io_flow(x477_1_io_flow),
    .io_result(x477_1_io_result)
  );
  x475 x478_1 ( // @[Math.scala 262:24:@45967.4]
    .clock(x478_1_clock),
    .io_a(x478_1_io_a),
    .io_b(x478_1_io_b),
    .io_flow(x478_1_io_flow),
    .io_result(x478_1_io_result)
  );
  x475 x479_1 ( // @[Math.scala 262:24:@45979.4]
    .clock(x479_1_clock),
    .io_a(x479_1_io_a),
    .io_b(x479_1_io_b),
    .io_flow(x479_1_io_flow),
    .io_result(x479_1_io_result)
  );
  x475 x480_1 ( // @[Math.scala 262:24:@45991.4]
    .clock(x480_1_clock),
    .io_a(x480_1_io_a),
    .io_b(x480_1_io_b),
    .io_flow(x480_1_io_flow),
    .io_result(x480_1_io_result)
  );
  x475 x481_1 ( // @[Math.scala 262:24:@46003.4]
    .clock(x481_1_clock),
    .io_a(x481_1_io_a),
    .io_b(x481_1_io_b),
    .io_flow(x481_1_io_flow),
    .io_result(x481_1_io_result)
  );
  x475 x482_1 ( // @[Math.scala 262:24:@46015.4]
    .clock(x482_1_clock),
    .io_a(x482_1_io_a),
    .io_b(x482_1_io_b),
    .io_flow(x482_1_io_flow),
    .io_result(x482_1_io_result)
  );
  x475 x483_1 ( // @[Math.scala 262:24:@46027.4]
    .clock(x483_1_clock),
    .io_a(x483_1_io_a),
    .io_b(x483_1_io_b),
    .io_flow(x483_1_io_flow),
    .io_result(x483_1_io_result)
  );
  x484_x3 x484_x3_1 ( // @[Math.scala 150:24:@46037.4]
    .clock(x484_x3_1_clock),
    .reset(x484_x3_1_reset),
    .io_a(x484_x3_1_io_a),
    .io_b(x484_x3_1_io_b),
    .io_flow(x484_x3_1_io_flow),
    .io_result(x484_x3_1_io_result)
  );
  x484_x3 x485_x4_1 ( // @[Math.scala 150:24:@46047.4]
    .clock(x485_x4_1_clock),
    .reset(x485_x4_1_reset),
    .io_a(x485_x4_1_io_a),
    .io_b(x485_x4_1_io_b),
    .io_flow(x485_x4_1_io_flow),
    .io_result(x485_x4_1_io_result)
  );
  x484_x3 x486_x3_1 ( // @[Math.scala 150:24:@46057.4]
    .clock(x486_x3_1_clock),
    .reset(x486_x3_1_reset),
    .io_a(x486_x3_1_io_a),
    .io_b(x486_x3_1_io_b),
    .io_flow(x486_x3_1_io_flow),
    .io_result(x486_x3_1_io_result)
  );
  x484_x3 x487_x4_1 ( // @[Math.scala 150:24:@46067.4]
    .clock(x487_x4_1_clock),
    .reset(x487_x4_1_reset),
    .io_a(x487_x4_1_io_a),
    .io_b(x487_x4_1_io_b),
    .io_flow(x487_x4_1_io_flow),
    .io_result(x487_x4_1_io_result)
  );
  x484_x3 x488_x3_1 ( // @[Math.scala 150:24:@46077.4]
    .clock(x488_x3_1_clock),
    .reset(x488_x3_1_reset),
    .io_a(x488_x3_1_io_a),
    .io_b(x488_x3_1_io_b),
    .io_flow(x488_x3_1_io_flow),
    .io_result(x488_x3_1_io_result)
  );
  x484_x3 x489_x4_1 ( // @[Math.scala 150:24:@46087.4]
    .clock(x489_x4_1_clock),
    .reset(x489_x4_1_reset),
    .io_a(x489_x4_1_io_a),
    .io_b(x489_x4_1_io_b),
    .io_flow(x489_x4_1_io_flow),
    .io_result(x489_x4_1_io_result)
  );
  x484_x3 x490_x3_1 ( // @[Math.scala 150:24:@46097.4]
    .clock(x490_x3_1_clock),
    .reset(x490_x3_1_reset),
    .io_a(x490_x3_1_io_a),
    .io_b(x490_x3_1_io_b),
    .io_flow(x490_x3_1_io_flow),
    .io_result(x490_x3_1_io_result)
  );
  RetimeWrapper_301 RetimeWrapper_104 ( // @[package.scala 93:22:@46107.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  x484_x3 x491_sum_1 ( // @[Math.scala 150:24:@46116.4]
    .clock(x491_sum_1_clock),
    .reset(x491_sum_1_reset),
    .io_a(x491_sum_1_io_a),
    .io_b(x491_sum_1_io_b),
    .io_flow(x491_sum_1_io_flow),
    .io_result(x491_sum_1_io_result)
  );
  x492 x492_1 ( // @[Math.scala 720:24:@46126.4]
    .io_b(x492_1_io_b),
    .io_result(x492_1_io_result)
  );
  x493_mul x493_mul_1 ( // @[Math.scala 262:24:@46137.4]
    .clock(x493_mul_1_clock),
    .io_a(x493_mul_1_io_a),
    .io_flow(x493_mul_1_io_flow),
    .io_result(x493_mul_1_io_result)
  );
  x494 x494_1 ( // @[Math.scala 720:24:@46147.4]
    .io_b(x494_1_io_b),
    .io_result(x494_1_io_result)
  );
  x475 x495_1 ( // @[Math.scala 262:24:@46158.4]
    .clock(x495_1_clock),
    .io_a(x495_1_io_a),
    .io_b(x495_1_io_b),
    .io_flow(x495_1_io_flow),
    .io_result(x495_1_io_result)
  );
  x475 x496_1 ( // @[Math.scala 262:24:@46170.4]
    .clock(x496_1_clock),
    .io_a(x496_1_io_a),
    .io_b(x496_1_io_b),
    .io_flow(x496_1_io_flow),
    .io_result(x496_1_io_result)
  );
  x475 x497_1 ( // @[Math.scala 262:24:@46182.4]
    .clock(x497_1_clock),
    .io_a(x497_1_io_a),
    .io_b(x497_1_io_b),
    .io_flow(x497_1_io_flow),
    .io_result(x497_1_io_result)
  );
  x475 x498_1 ( // @[Math.scala 262:24:@46194.4]
    .clock(x498_1_clock),
    .io_a(x498_1_io_a),
    .io_b(x498_1_io_b),
    .io_flow(x498_1_io_flow),
    .io_result(x498_1_io_result)
  );
  x475 x499_1 ( // @[Math.scala 262:24:@46206.4]
    .clock(x499_1_clock),
    .io_a(x499_1_io_a),
    .io_b(x499_1_io_b),
    .io_flow(x499_1_io_flow),
    .io_result(x499_1_io_result)
  );
  x475 x500_1 ( // @[Math.scala 262:24:@46218.4]
    .clock(x500_1_clock),
    .io_a(x500_1_io_a),
    .io_b(x500_1_io_b),
    .io_flow(x500_1_io_flow),
    .io_result(x500_1_io_result)
  );
  x475 x501_1 ( // @[Math.scala 262:24:@46232.4]
    .clock(x501_1_clock),
    .io_a(x501_1_io_a),
    .io_b(x501_1_io_b),
    .io_flow(x501_1_io_flow),
    .io_result(x501_1_io_result)
  );
  x475 x502_1 ( // @[Math.scala 262:24:@46244.4]
    .clock(x502_1_clock),
    .io_a(x502_1_io_a),
    .io_b(x502_1_io_b),
    .io_flow(x502_1_io_flow),
    .io_result(x502_1_io_result)
  );
  x475 x503_1 ( // @[Math.scala 262:24:@46256.4]
    .clock(x503_1_clock),
    .io_a(x503_1_io_a),
    .io_b(x503_1_io_b),
    .io_flow(x503_1_io_flow),
    .io_result(x503_1_io_result)
  );
  x484_x3 x504_x3_1 ( // @[Math.scala 150:24:@46266.4]
    .clock(x504_x3_1_clock),
    .reset(x504_x3_1_reset),
    .io_a(x504_x3_1_io_a),
    .io_b(x504_x3_1_io_b),
    .io_flow(x504_x3_1_io_flow),
    .io_result(x504_x3_1_io_result)
  );
  x484_x3 x505_x4_1 ( // @[Math.scala 150:24:@46276.4]
    .clock(x505_x4_1_clock),
    .reset(x505_x4_1_reset),
    .io_a(x505_x4_1_io_a),
    .io_b(x505_x4_1_io_b),
    .io_flow(x505_x4_1_io_flow),
    .io_result(x505_x4_1_io_result)
  );
  x484_x3 x506_x3_1 ( // @[Math.scala 150:24:@46286.4]
    .clock(x506_x3_1_clock),
    .reset(x506_x3_1_reset),
    .io_a(x506_x3_1_io_a),
    .io_b(x506_x3_1_io_b),
    .io_flow(x506_x3_1_io_flow),
    .io_result(x506_x3_1_io_result)
  );
  x484_x3 x507_x4_1 ( // @[Math.scala 150:24:@46296.4]
    .clock(x507_x4_1_clock),
    .reset(x507_x4_1_reset),
    .io_a(x507_x4_1_io_a),
    .io_b(x507_x4_1_io_b),
    .io_flow(x507_x4_1_io_flow),
    .io_result(x507_x4_1_io_result)
  );
  x484_x3 x508_x3_1 ( // @[Math.scala 150:24:@46306.4]
    .clock(x508_x3_1_clock),
    .reset(x508_x3_1_reset),
    .io_a(x508_x3_1_io_a),
    .io_b(x508_x3_1_io_b),
    .io_flow(x508_x3_1_io_flow),
    .io_result(x508_x3_1_io_result)
  );
  x484_x3 x509_x4_1 ( // @[Math.scala 150:24:@46316.4]
    .clock(x509_x4_1_clock),
    .reset(x509_x4_1_reset),
    .io_a(x509_x4_1_io_a),
    .io_b(x509_x4_1_io_b),
    .io_flow(x509_x4_1_io_flow),
    .io_result(x509_x4_1_io_result)
  );
  x484_x3 x510_x3_1 ( // @[Math.scala 150:24:@46326.4]
    .clock(x510_x3_1_clock),
    .reset(x510_x3_1_reset),
    .io_a(x510_x3_1_io_a),
    .io_b(x510_x3_1_io_b),
    .io_flow(x510_x3_1_io_flow),
    .io_result(x510_x3_1_io_result)
  );
  RetimeWrapper_301 RetimeWrapper_105 ( // @[package.scala 93:22:@46336.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  x484_x3 x511_sum_1 ( // @[Math.scala 150:24:@46345.4]
    .clock(x511_sum_1_clock),
    .reset(x511_sum_1_reset),
    .io_a(x511_sum_1_io_a),
    .io_b(x511_sum_1_io_b),
    .io_flow(x511_sum_1_io_flow),
    .io_result(x511_sum_1_io_result)
  );
  x492 x512_1 ( // @[Math.scala 720:24:@46355.4]
    .io_b(x512_1_io_b),
    .io_result(x512_1_io_result)
  );
  x493_mul x513_mul_1 ( // @[Math.scala 262:24:@46366.4]
    .clock(x513_mul_1_clock),
    .io_a(x513_mul_1_io_a),
    .io_flow(x513_mul_1_io_flow),
    .io_result(x513_mul_1_io_result)
  );
  x494 x514_1 ( // @[Math.scala 720:24:@46376.4]
    .io_b(x514_1_io_b),
    .io_result(x514_1_io_result)
  );
  x475 x515_1 ( // @[Math.scala 262:24:@46387.4]
    .clock(x515_1_clock),
    .io_a(x515_1_io_a),
    .io_b(x515_1_io_b),
    .io_flow(x515_1_io_flow),
    .io_result(x515_1_io_result)
  );
  x475 x516_1 ( // @[Math.scala 262:24:@46399.4]
    .clock(x516_1_clock),
    .io_a(x516_1_io_a),
    .io_b(x516_1_io_b),
    .io_flow(x516_1_io_flow),
    .io_result(x516_1_io_result)
  );
  x475 x517_1 ( // @[Math.scala 262:24:@46411.4]
    .clock(x517_1_clock),
    .io_a(x517_1_io_a),
    .io_b(x517_1_io_b),
    .io_flow(x517_1_io_flow),
    .io_result(x517_1_io_result)
  );
  x475 x518_1 ( // @[Math.scala 262:24:@46423.4]
    .clock(x518_1_clock),
    .io_a(x518_1_io_a),
    .io_b(x518_1_io_b),
    .io_flow(x518_1_io_flow),
    .io_result(x518_1_io_result)
  );
  x475 x519_1 ( // @[Math.scala 262:24:@46435.4]
    .clock(x519_1_clock),
    .io_a(x519_1_io_a),
    .io_b(x519_1_io_b),
    .io_flow(x519_1_io_flow),
    .io_result(x519_1_io_result)
  );
  x475 x520_1 ( // @[Math.scala 262:24:@46447.4]
    .clock(x520_1_clock),
    .io_a(x520_1_io_a),
    .io_b(x520_1_io_b),
    .io_flow(x520_1_io_flow),
    .io_result(x520_1_io_result)
  );
  x484_x3 x521_x3_1 ( // @[Math.scala 150:24:@46457.4]
    .clock(x521_x3_1_clock),
    .reset(x521_x3_1_reset),
    .io_a(x521_x3_1_io_a),
    .io_b(x521_x3_1_io_b),
    .io_flow(x521_x3_1_io_flow),
    .io_result(x521_x3_1_io_result)
  );
  x484_x3 x522_x4_1 ( // @[Math.scala 150:24:@46467.4]
    .clock(x522_x4_1_clock),
    .reset(x522_x4_1_reset),
    .io_a(x522_x4_1_io_a),
    .io_b(x522_x4_1_io_b),
    .io_flow(x522_x4_1_io_flow),
    .io_result(x522_x4_1_io_result)
  );
  x484_x3 x523_x3_1 ( // @[Math.scala 150:24:@46477.4]
    .clock(x523_x3_1_clock),
    .reset(x523_x3_1_reset),
    .io_a(x523_x3_1_io_a),
    .io_b(x523_x3_1_io_b),
    .io_flow(x523_x3_1_io_flow),
    .io_result(x523_x3_1_io_result)
  );
  x484_x3 x524_x4_1 ( // @[Math.scala 150:24:@46487.4]
    .clock(x524_x4_1_clock),
    .reset(x524_x4_1_reset),
    .io_a(x524_x4_1_io_a),
    .io_b(x524_x4_1_io_b),
    .io_flow(x524_x4_1_io_flow),
    .io_result(x524_x4_1_io_result)
  );
  x484_x3 x525_x3_1 ( // @[Math.scala 150:24:@46497.4]
    .clock(x525_x3_1_clock),
    .reset(x525_x3_1_reset),
    .io_a(x525_x3_1_io_a),
    .io_b(x525_x3_1_io_b),
    .io_flow(x525_x3_1_io_flow),
    .io_result(x525_x3_1_io_result)
  );
  x484_x3 x526_x4_1 ( // @[Math.scala 150:24:@46507.4]
    .clock(x526_x4_1_clock),
    .reset(x526_x4_1_reset),
    .io_a(x526_x4_1_io_a),
    .io_b(x526_x4_1_io_b),
    .io_flow(x526_x4_1_io_flow),
    .io_result(x526_x4_1_io_result)
  );
  x484_x3 x527_x3_1 ( // @[Math.scala 150:24:@46517.4]
    .clock(x527_x3_1_clock),
    .reset(x527_x3_1_reset),
    .io_a(x527_x3_1_io_a),
    .io_b(x527_x3_1_io_b),
    .io_flow(x527_x3_1_io_flow),
    .io_result(x527_x3_1_io_result)
  );
  RetimeWrapper_301 RetimeWrapper_106 ( // @[package.scala 93:22:@46527.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  x484_x3 x528_sum_1 ( // @[Math.scala 150:24:@46536.4]
    .clock(x528_sum_1_clock),
    .reset(x528_sum_1_reset),
    .io_a(x528_sum_1_io_a),
    .io_b(x528_sum_1_io_b),
    .io_flow(x528_sum_1_io_flow),
    .io_result(x528_sum_1_io_result)
  );
  x492 x529_1 ( // @[Math.scala 720:24:@46546.4]
    .io_b(x529_1_io_b),
    .io_result(x529_1_io_result)
  );
  x493_mul x530_mul_1 ( // @[Math.scala 262:24:@46557.4]
    .clock(x530_mul_1_clock),
    .io_a(x530_mul_1_io_a),
    .io_flow(x530_mul_1_io_flow),
    .io_result(x530_mul_1_io_result)
  );
  x494 x531_1 ( // @[Math.scala 720:24:@46567.4]
    .io_b(x531_1_io_b),
    .io_result(x531_1_io_result)
  );
  x475 x532_1 ( // @[Math.scala 262:24:@46578.4]
    .clock(x532_1_clock),
    .io_a(x532_1_io_a),
    .io_b(x532_1_io_b),
    .io_flow(x532_1_io_flow),
    .io_result(x532_1_io_result)
  );
  x475 x533_1 ( // @[Math.scala 262:24:@46590.4]
    .clock(x533_1_clock),
    .io_a(x533_1_io_a),
    .io_b(x533_1_io_b),
    .io_flow(x533_1_io_flow),
    .io_result(x533_1_io_result)
  );
  x475 x534_1 ( // @[Math.scala 262:24:@46602.4]
    .clock(x534_1_clock),
    .io_a(x534_1_io_a),
    .io_b(x534_1_io_b),
    .io_flow(x534_1_io_flow),
    .io_result(x534_1_io_result)
  );
  x475 x535_1 ( // @[Math.scala 262:24:@46614.4]
    .clock(x535_1_clock),
    .io_a(x535_1_io_a),
    .io_b(x535_1_io_b),
    .io_flow(x535_1_io_flow),
    .io_result(x535_1_io_result)
  );
  x475 x536_1 ( // @[Math.scala 262:24:@46626.4]
    .clock(x536_1_clock),
    .io_a(x536_1_io_a),
    .io_b(x536_1_io_b),
    .io_flow(x536_1_io_flow),
    .io_result(x536_1_io_result)
  );
  x475 x537_1 ( // @[Math.scala 262:24:@46638.4]
    .clock(x537_1_clock),
    .io_a(x537_1_io_a),
    .io_b(x537_1_io_b),
    .io_flow(x537_1_io_flow),
    .io_result(x537_1_io_result)
  );
  x484_x3 x538_x3_1 ( // @[Math.scala 150:24:@46648.4]
    .clock(x538_x3_1_clock),
    .reset(x538_x3_1_reset),
    .io_a(x538_x3_1_io_a),
    .io_b(x538_x3_1_io_b),
    .io_flow(x538_x3_1_io_flow),
    .io_result(x538_x3_1_io_result)
  );
  x484_x3 x539_x4_1 ( // @[Math.scala 150:24:@46658.4]
    .clock(x539_x4_1_clock),
    .reset(x539_x4_1_reset),
    .io_a(x539_x4_1_io_a),
    .io_b(x539_x4_1_io_b),
    .io_flow(x539_x4_1_io_flow),
    .io_result(x539_x4_1_io_result)
  );
  x484_x3 x540_x3_1 ( // @[Math.scala 150:24:@46668.4]
    .clock(x540_x3_1_clock),
    .reset(x540_x3_1_reset),
    .io_a(x540_x3_1_io_a),
    .io_b(x540_x3_1_io_b),
    .io_flow(x540_x3_1_io_flow),
    .io_result(x540_x3_1_io_result)
  );
  x484_x3 x541_x4_1 ( // @[Math.scala 150:24:@46678.4]
    .clock(x541_x4_1_clock),
    .reset(x541_x4_1_reset),
    .io_a(x541_x4_1_io_a),
    .io_b(x541_x4_1_io_b),
    .io_flow(x541_x4_1_io_flow),
    .io_result(x541_x4_1_io_result)
  );
  x484_x3 x542_x3_1 ( // @[Math.scala 150:24:@46688.4]
    .clock(x542_x3_1_clock),
    .reset(x542_x3_1_reset),
    .io_a(x542_x3_1_io_a),
    .io_b(x542_x3_1_io_b),
    .io_flow(x542_x3_1_io_flow),
    .io_result(x542_x3_1_io_result)
  );
  x484_x3 x543_x4_1 ( // @[Math.scala 150:24:@46698.4]
    .clock(x543_x4_1_clock),
    .reset(x543_x4_1_reset),
    .io_a(x543_x4_1_io_a),
    .io_b(x543_x4_1_io_b),
    .io_flow(x543_x4_1_io_flow),
    .io_result(x543_x4_1_io_result)
  );
  x484_x3 x544_x3_1 ( // @[Math.scala 150:24:@46708.4]
    .clock(x544_x3_1_clock),
    .reset(x544_x3_1_reset),
    .io_a(x544_x3_1_io_a),
    .io_b(x544_x3_1_io_b),
    .io_flow(x544_x3_1_io_flow),
    .io_result(x544_x3_1_io_result)
  );
  RetimeWrapper_301 RetimeWrapper_107 ( // @[package.scala 93:22:@46718.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  x484_x3 x545_sum_1 ( // @[Math.scala 150:24:@46727.4]
    .clock(x545_sum_1_clock),
    .reset(x545_sum_1_reset),
    .io_a(x545_sum_1_io_a),
    .io_b(x545_sum_1_io_b),
    .io_flow(x545_sum_1_io_flow),
    .io_result(x545_sum_1_io_result)
  );
  x492 x546_1 ( // @[Math.scala 720:24:@46737.4]
    .io_b(x546_1_io_b),
    .io_result(x546_1_io_result)
  );
  x493_mul x547_mul_1 ( // @[Math.scala 262:24:@46750.4]
    .clock(x547_mul_1_clock),
    .io_a(x547_mul_1_io_a),
    .io_flow(x547_mul_1_io_flow),
    .io_result(x547_mul_1_io_result)
  );
  x494 x548_1 ( // @[Math.scala 720:24:@46760.4]
    .io_b(x548_1_io_b),
    .io_result(x548_1_io_result)
  );
  RetimeWrapper_464 RetimeWrapper_108 ( // @[package.scala 93:22:@46779.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_109 ( // @[package.scala 93:22:@46788.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_110 ( // @[package.scala 93:22:@46797.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_111 ( // @[package.scala 93:22:@46806.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  assign b330 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 62:18:@43744.4]
  assign b331 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 63:18:@43745.4]
  assign _T_205 = b330 & b331; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 67:30:@43747.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 67:37:@43748.4]
  assign _T_210 = io_in_x289_TID == 8'h0; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 69:76:@43753.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 69:62:@43754.4]
  assign _T_213 = io_in_x289_TDEST == 8'h0; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 69:101:@43755.4]
  assign x637_x332_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@43764.4 package.scala 96:25:@43765.4]
  assign b328_number = __io_result; // @[Math.scala 723:22:@43729.4 Math.scala 724:14:@43730.4]
  assign _T_247 = $signed(b328_number); // @[Math.scala 406:49:@43929.4]
  assign _T_249 = $signed(_T_247) & $signed(32'sh3); // @[Math.scala 406:56:@43931.4]
  assign _T_250 = $signed(_T_249); // @[Math.scala 406:56:@43932.4]
  assign x617_number = $unsigned(_T_250); // @[implicits.scala 133:21:@43933.4]
  assign _T_260 = $signed(x617_number); // @[Math.scala 406:49:@43942.4]
  assign _T_262 = $signed(_T_260) & $signed(32'sh3); // @[Math.scala 406:56:@43944.4]
  assign _T_263 = $signed(_T_262); // @[Math.scala 406:56:@43945.4]
  assign _T_274 = x617_number[31]; // @[FixedPoint.scala 50:25:@43963.4]
  assign _T_278 = _T_274 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@43965.4]
  assign _T_279 = x617_number[31:2]; // @[FixedPoint.scala 18:52:@43966.4]
  assign _T_285 = _T_279 == 30'h3fffffff; // @[Math.scala 451:55:@43968.4]
  assign _T_286 = x617_number[1:0]; // @[FixedPoint.scala 18:52:@43969.4]
  assign _T_292 = _T_286 != 2'h0; // @[Math.scala 451:110:@43971.4]
  assign _T_293 = _T_285 & _T_292; // @[Math.scala 451:94:@43972.4]
  assign _T_295 = {_T_278,_T_279}; // @[Cat.scala 30:58:@43974.4]
  assign x340_1_number = _T_293 ? 32'h0 : _T_295; // @[Math.scala 454:20:@43975.4]
  assign _GEN_0 = {{8'd0}, x340_1_number}; // @[Math.scala 461:32:@43980.4]
  assign _T_300 = _GEN_0 << 8; // @[Math.scala 461:32:@43980.4]
  assign _GEN_1 = {{6'd0}, x340_1_number}; // @[Math.scala 461:32:@43985.4]
  assign _T_303 = _GEN_1 << 6; // @[Math.scala 461:32:@43985.4]
  assign _T_339 = ~ io_sigsIn_break; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 117:101:@44083.4]
  assign _T_343 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@44091.4 package.scala 96:25:@44092.4]
  assign _T_345 = io_rr ? _T_343 : 1'h0; // @[implicits.scala 55:10:@44093.4]
  assign _T_346 = _T_339 & _T_345; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 117:118:@44094.4]
  assign _T_348 = _T_346 & _T_339; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 117:207:@44096.4]
  assign _T_349 = _T_348 & io_sigsIn_backpressure; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 117:226:@44097.4]
  assign x642_b330_D24 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@44062.4 package.scala 96:25:@44063.4]
  assign _T_350 = _T_349 & x642_b330_D24; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 117:252:@44098.4]
  assign x643_b331_D24 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@44071.4 package.scala 96:25:@44072.4]
  assign _T_394 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@44198.4 package.scala 96:25:@44199.4]
  assign _T_396 = io_rr ? _T_394 : 1'h0; // @[implicits.scala 55:10:@44200.4]
  assign _T_397 = _T_339 & _T_396; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 140:118:@44201.4]
  assign _T_399 = _T_397 & _T_339; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 140:207:@44203.4]
  assign _T_400 = _T_399 & io_sigsIn_backpressure; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 140:226:@44204.4]
  assign _T_401 = _T_400 & x642_b330_D24; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 140:252:@44205.4]
  assign _T_442 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@44296.4 package.scala 96:25:@44297.4]
  assign _T_444 = io_rr ? _T_442 : 1'h0; // @[implicits.scala 55:10:@44298.4]
  assign _T_445 = _T_339 & _T_444; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 161:118:@44299.4]
  assign _T_447 = _T_445 & _T_339; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 161:207:@44301.4]
  assign _T_448 = _T_447 & io_sigsIn_backpressure; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 161:226:@44302.4]
  assign _T_449 = _T_448 & x642_b330_D24; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 161:252:@44303.4]
  assign _T_490 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@44394.4 package.scala 96:25:@44395.4]
  assign _T_492 = io_rr ? _T_490 : 1'h0; // @[implicits.scala 55:10:@44396.4]
  assign _T_493 = _T_339 & _T_492; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 188:166:@44397.4]
  assign _T_495 = _T_493 & _T_339; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 188:255:@44399.4]
  assign _T_496 = _T_495 & io_sigsIn_backpressure; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 188:274:@44400.4]
  assign _T_497 = _T_496 & x642_b330_D24; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 188:300:@44401.4]
  assign x655_b328_D26_number = RetimeWrapper_22_io_out; // @[package.scala 96:25:@44415.4 package.scala 96:25:@44416.4]
  assign _T_509 = $signed(x655_b328_D26_number); // @[Math.scala 476:37:@44423.4]
  assign x656_x357_rdcol_D26_number = RetimeWrapper_24_io_out; // @[package.scala 96:25:@44440.4 package.scala 96:25:@44441.4]
  assign _T_522 = $signed(x656_x357_rdcol_D26_number); // @[Math.scala 476:37:@44446.4]
  assign x657_x364_D1 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@44463.4 package.scala 96:25:@44464.4]
  assign x365 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@44454.4 package.scala 96:25:@44455.4]
  assign x366 = x657_x364_D1 | x365; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 203:24:@44467.4]
  assign _T_563 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@44535.4 package.scala 96:25:@44536.4]
  assign _T_565 = io_rr ? _T_563 : 1'h0; // @[implicits.scala 55:10:@44537.4]
  assign _T_566 = _T_339 & _T_565; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 222:194:@44538.4]
  assign x660_x367_D20 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@44496.4 package.scala 96:25:@44497.4]
  assign _T_567 = _T_566 & x660_x367_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 222:283:@44539.4]
  assign x661_b330_D48 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@44505.4 package.scala 96:25:@44506.4]
  assign _T_568 = _T_567 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 222:291:@44540.4]
  assign x662_b331_D48 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@44514.4 package.scala 96:25:@44515.4]
  assign x664_x351_rdcol_D26_number = RetimeWrapper_34_io_out; // @[package.scala 96:25:@44556.4 package.scala 96:25:@44557.4]
  assign _T_579 = $signed(x664_x351_rdcol_D26_number); // @[Math.scala 476:37:@44562.4]
  assign x370 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@44570.4 package.scala 96:25:@44571.4]
  assign x371 = x657_x364_D1 | x370; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 230:24:@44574.4]
  assign _T_608 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@44615.4 package.scala 96:25:@44616.4]
  assign _T_610 = io_rr ? _T_608 : 1'h0; // @[implicits.scala 55:10:@44617.4]
  assign _T_611 = _T_339 & _T_610; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 243:194:@44618.4]
  assign x665_x372_D20 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@44585.4 package.scala 96:25:@44586.4]
  assign _T_612 = _T_611 & x665_x372_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 243:283:@44619.4]
  assign _T_613 = _T_612 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 243:291:@44620.4]
  assign x668_x345_rdcol_D26_number = RetimeWrapper_40_io_out; // @[package.scala 96:25:@44636.4 package.scala 96:25:@44637.4]
  assign _T_624 = $signed(x668_x345_rdcol_D26_number); // @[Math.scala 476:37:@44642.4]
  assign x375 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@44650.4 package.scala 96:25:@44651.4]
  assign x376 = x657_x364_D1 | x375; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 251:24:@44654.4]
  assign _T_653 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@44695.4 package.scala 96:25:@44696.4]
  assign _T_655 = io_rr ? _T_653 : 1'h0; // @[implicits.scala 55:10:@44697.4]
  assign _T_656 = _T_339 & _T_655; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 264:194:@44698.4]
  assign x671_x377_D20 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@44683.4 package.scala 96:25:@44684.4]
  assign _T_657 = _T_656 & x671_x377_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 264:283:@44699.4]
  assign _T_658 = _T_657 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 264:291:@44700.4]
  assign x672_b329_D26_number = RetimeWrapper_46_io_out; // @[package.scala 96:25:@44716.4 package.scala 96:25:@44717.4]
  assign _T_669 = $signed(x672_b329_D26_number); // @[Math.scala 476:37:@44722.4]
  assign x364 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@44431.4 package.scala 96:25:@44432.4]
  assign x380 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@44730.4 package.scala 96:25:@44731.4]
  assign x381 = x364 | x380; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 272:24:@44734.4]
  assign _T_698 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@44775.4 package.scala 96:25:@44776.4]
  assign _T_700 = io_rr ? _T_698 : 1'h0; // @[implicits.scala 55:10:@44777.4]
  assign _T_701 = _T_339 & _T_700; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 285:194:@44778.4]
  assign x675_x382_D21 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@44763.4 package.scala 96:25:@44764.4]
  assign _T_702 = _T_701 & x675_x382_D21; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 285:283:@44779.4]
  assign _T_703 = _T_702 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 285:291:@44780.4]
  assign x385_rdcol_number = x385_rdcol_1_io_result; // @[Math.scala 154:22:@44799.4 Math.scala 155:14:@44800.4]
  assign _T_718 = $signed(x385_rdcol_number); // @[Math.scala 476:37:@44805.4]
  assign x386 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@44813.4 package.scala 96:25:@44814.4]
  assign x387 = x657_x364_D1 | x386; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 293:24:@44817.4]
  assign _T_766 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@44894.4 package.scala 96:25:@44895.4]
  assign _T_768 = io_rr ? _T_766 : 1'h0; // @[implicits.scala 55:10:@44896.4]
  assign _T_769 = _T_339 & _T_768; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 320:194:@44897.4]
  assign x678_x388_D20 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@44882.4 package.scala 96:25:@44883.4]
  assign _T_770 = _T_769 & x678_x388_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 320:283:@44898.4]
  assign _T_771 = _T_770 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 320:291:@44899.4]
  assign x394_rdcol_number = x394_rdcol_1_io_result; // @[Math.scala 154:22:@44918.4 Math.scala 155:14:@44919.4]
  assign _T_786 = $signed(x394_rdcol_number); // @[Math.scala 476:37:@44924.4]
  assign x395 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@44932.4 package.scala 96:25:@44933.4]
  assign x396 = x657_x364_D1 | x395; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 328:59:@44936.4]
  assign _T_829 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@45002.4 package.scala 96:25:@45003.4]
  assign _T_831 = io_rr ? _T_829 : 1'h0; // @[implicits.scala 55:10:@45004.4]
  assign _T_832 = _T_339 & _T_831; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 345:194:@45005.4]
  assign x679_x397_D20 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@44981.4 package.scala 96:25:@44982.4]
  assign _T_833 = _T_832 & x679_x397_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 345:283:@45006.4]
  assign _T_834 = _T_833 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 345:291:@45007.4]
  assign x403_rdrow_number = x403_rdrow_1_io_result; // @[Math.scala 195:22:@45026.4 Math.scala 196:14:@45027.4]
  assign _T_851 = $signed(x403_rdrow_number); // @[Math.scala 406:49:@45033.4]
  assign _T_853 = $signed(_T_851) & $signed(32'sh3); // @[Math.scala 406:56:@45035.4]
  assign _T_854 = $signed(_T_853); // @[Math.scala 406:56:@45036.4]
  assign x622_number = $unsigned(_T_854); // @[implicits.scala 133:21:@45037.4]
  assign x405 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@45051.4 package.scala 96:25:@45052.4]
  assign x406 = x405 | x365; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 355:24:@45055.4]
  assign _T_877 = $signed(x622_number); // @[Math.scala 406:49:@45064.4]
  assign _T_879 = $signed(_T_877) & $signed(32'sh3); // @[Math.scala 406:56:@45066.4]
  assign _T_880 = $signed(_T_879); // @[Math.scala 406:56:@45067.4]
  assign _T_884 = $signed(RetimeWrapper_62_io_out); // @[package.scala 96:25:@45075.4]
  assign _T_888 = x622_number[31]; // @[FixedPoint.scala 50:25:@45082.4]
  assign _T_892 = _T_888 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@45084.4]
  assign _T_893 = x622_number[31:2]; // @[FixedPoint.scala 18:52:@45085.4]
  assign _T_899 = _T_893 == 30'h3fffffff; // @[Math.scala 451:55:@45087.4]
  assign _T_900 = x622_number[1:0]; // @[FixedPoint.scala 18:52:@45088.4]
  assign _T_906 = _T_900 != 2'h0; // @[Math.scala 451:110:@45090.4]
  assign _T_907 = _T_899 & _T_906; // @[Math.scala 451:94:@45091.4]
  assign _T_911 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@45099.4 package.scala 96:25:@45100.4]
  assign x409_1_number = _T_907 ? 32'h0 : _T_911; // @[Math.scala 454:20:@45101.4]
  assign _GEN_2 = {{8'd0}, x409_1_number}; // @[Math.scala 461:32:@45106.4]
  assign _T_916 = _GEN_2 << 8; // @[Math.scala 461:32:@45106.4]
  assign _GEN_3 = {{6'd0}, x409_1_number}; // @[Math.scala 461:32:@45111.4]
  assign _T_919 = _GEN_3 << 6; // @[Math.scala 461:32:@45111.4]
  assign _T_949 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@45179.4 package.scala 96:25:@45180.4]
  assign _T_951 = io_rr ? _T_949 : 1'h0; // @[implicits.scala 55:10:@45181.4]
  assign _T_952 = _T_339 & _T_951; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 382:194:@45182.4]
  assign x684_x407_D20 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@45167.4 package.scala 96:25:@45168.4]
  assign _T_953 = _T_952 & x684_x407_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 382:283:@45183.4]
  assign _T_954 = _T_953 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 382:291:@45184.4]
  assign x414 = x405 | x370; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 386:24:@45195.4]
  assign _T_981 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@45237.4 package.scala 96:25:@45238.4]
  assign _T_983 = io_rr ? _T_981 : 1'h0; // @[implicits.scala 55:10:@45239.4]
  assign _T_984 = _T_339 & _T_983; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 399:194:@45240.4]
  assign x686_x415_D20 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@45225.4 package.scala 96:25:@45226.4]
  assign _T_985 = _T_984 & x686_x415_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 399:283:@45241.4]
  assign _T_986 = _T_985 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 399:291:@45242.4]
  assign x419 = x405 | x375; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 403:24:@45253.4]
  assign _T_1013 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@45295.4 package.scala 96:25:@45296.4]
  assign _T_1015 = io_rr ? _T_1013 : 1'h0; // @[implicits.scala 55:10:@45297.4]
  assign _T_1016 = _T_339 & _T_1015; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 416:194:@45298.4]
  assign x688_x420_D20 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@45283.4 package.scala 96:25:@45284.4]
  assign _T_1017 = _T_1016 & x688_x420_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 416:283:@45299.4]
  assign _T_1018 = _T_1017 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 416:291:@45300.4]
  assign x689_x380_D1 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@45316.4 package.scala 96:25:@45317.4]
  assign x424 = x405 | x689_x380_D1; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 428:59:@45320.4]
  assign _T_1056 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@45382.4 package.scala 96:25:@45383.4]
  assign _T_1058 = io_rr ? _T_1056 : 1'h0; // @[implicits.scala 55:10:@45384.4]
  assign _T_1059 = _T_339 & _T_1058; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 447:194:@45385.4]
  assign x692_x425_D20 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@45361.4 package.scala 96:25:@45362.4]
  assign _T_1060 = _T_1059 & x692_x425_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 447:283:@45386.4]
  assign _T_1061 = _T_1060 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 447:291:@45387.4]
  assign x429 = x405 | x386; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 451:59:@45398.4]
  assign _T_1085 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@45431.4 package.scala 96:25:@45432.4]
  assign _T_1087 = io_rr ? _T_1085 : 1'h0; // @[implicits.scala 55:10:@45433.4]
  assign _T_1088 = _T_339 & _T_1087; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 462:194:@45434.4]
  assign x694_x430_D20 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@45419.4 package.scala 96:25:@45420.4]
  assign _T_1089 = _T_1088 & x694_x430_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 462:283:@45435.4]
  assign _T_1090 = _T_1089 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 462:291:@45436.4]
  assign x434 = x405 | x395; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 466:59:@45447.4]
  assign _T_1114 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@45480.4 package.scala 96:25:@45481.4]
  assign _T_1116 = io_rr ? _T_1114 : 1'h0; // @[implicits.scala 55:10:@45482.4]
  assign _T_1117 = _T_339 & _T_1116; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 477:194:@45483.4]
  assign x695_x435_D20 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@45468.4 package.scala 96:25:@45469.4]
  assign _T_1118 = _T_1117 & x695_x435_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 477:283:@45484.4]
  assign _T_1119 = _T_1118 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 477:291:@45485.4]
  assign x439_rdrow_number = x439_rdrow_1_io_result; // @[Math.scala 195:22:@45504.4 Math.scala 196:14:@45505.4]
  assign _T_1136 = $signed(x439_rdrow_number); // @[Math.scala 406:49:@45511.4]
  assign _T_1138 = $signed(_T_1136) & $signed(32'sh3); // @[Math.scala 406:56:@45513.4]
  assign _T_1139 = $signed(_T_1138); // @[Math.scala 406:56:@45514.4]
  assign x627_number = $unsigned(_T_1139); // @[implicits.scala 133:21:@45515.4]
  assign x441 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@45529.4 package.scala 96:25:@45530.4]
  assign x442 = x441 | x365; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 487:24:@45533.4]
  assign _T_1162 = $signed(x627_number); // @[Math.scala 406:49:@45542.4]
  assign _T_1164 = $signed(_T_1162) & $signed(32'sh3); // @[Math.scala 406:56:@45544.4]
  assign _T_1165 = $signed(_T_1164); // @[Math.scala 406:56:@45545.4]
  assign _T_1169 = $signed(RetimeWrapper_86_io_out); // @[package.scala 96:25:@45553.4]
  assign _T_1173 = x627_number[31]; // @[FixedPoint.scala 50:25:@45560.4]
  assign _T_1177 = _T_1173 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@45562.4]
  assign _T_1178 = x627_number[31:2]; // @[FixedPoint.scala 18:52:@45563.4]
  assign _T_1184 = _T_1178 == 30'h3fffffff; // @[Math.scala 451:55:@45565.4]
  assign _T_1185 = x627_number[1:0]; // @[FixedPoint.scala 18:52:@45566.4]
  assign _T_1191 = _T_1185 != 2'h0; // @[Math.scala 451:110:@45568.4]
  assign _T_1192 = _T_1184 & _T_1191; // @[Math.scala 451:94:@45569.4]
  assign _T_1196 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@45577.4 package.scala 96:25:@45578.4]
  assign x445_1_number = _T_1192 ? 32'h0 : _T_1196; // @[Math.scala 454:20:@45579.4]
  assign _GEN_4 = {{8'd0}, x445_1_number}; // @[Math.scala 461:32:@45584.4]
  assign _T_1201 = _GEN_4 << 8; // @[Math.scala 461:32:@45584.4]
  assign _GEN_5 = {{6'd0}, x445_1_number}; // @[Math.scala 461:32:@45589.4]
  assign _T_1204 = _GEN_5 << 6; // @[Math.scala 461:32:@45589.4]
  assign _T_1231 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@45648.4 package.scala 96:25:@45649.4]
  assign _T_1233 = io_rr ? _T_1231 : 1'h0; // @[implicits.scala 55:10:@45650.4]
  assign _T_1234 = _T_339 & _T_1233; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 512:194:@45651.4]
  assign x698_x443_D20 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@45636.4 package.scala 96:25:@45637.4]
  assign _T_1235 = _T_1234 & x698_x443_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 512:283:@45652.4]
  assign _T_1236 = _T_1235 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 512:291:@45653.4]
  assign x450 = x441 | x370; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 516:24:@45664.4]
  assign _T_1260 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@45697.4 package.scala 96:25:@45698.4]
  assign _T_1262 = io_rr ? _T_1260 : 1'h0; // @[implicits.scala 55:10:@45699.4]
  assign _T_1263 = _T_339 & _T_1262; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 527:194:@45700.4]
  assign x699_x451_D20 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@45685.4 package.scala 96:25:@45686.4]
  assign _T_1264 = _T_1263 & x699_x451_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 527:283:@45701.4]
  assign _T_1265 = _T_1264 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 527:291:@45702.4]
  assign x455 = x441 | x375; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 531:24:@45713.4]
  assign _T_1289 = RetimeWrapper_95_io_out; // @[package.scala 96:25:@45746.4 package.scala 96:25:@45747.4]
  assign _T_1291 = io_rr ? _T_1289 : 1'h0; // @[implicits.scala 55:10:@45748.4]
  assign _T_1292 = _T_339 & _T_1291; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 548:194:@45749.4]
  assign x700_x456_D20 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@45734.4 package.scala 96:25:@45735.4]
  assign _T_1293 = _T_1292 & x700_x456_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 548:283:@45750.4]
  assign _T_1294 = _T_1293 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 548:326:@45751.4]
  assign x460 = x441 | x689_x380_D1; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 552:59:@45762.4]
  assign _T_1326 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@45815.4 package.scala 96:25:@45816.4]
  assign _T_1328 = io_rr ? _T_1326 : 1'h0; // @[implicits.scala 55:10:@45817.4]
  assign _T_1329 = _T_339 & _T_1328; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 569:194:@45818.4]
  assign x702_x461_D20 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@45794.4 package.scala 96:25:@45795.4]
  assign _T_1330 = _T_1329 & x702_x461_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 569:283:@45819.4]
  assign _T_1331 = _T_1330 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 569:291:@45820.4]
  assign x465 = x441 | x386; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 573:59:@45831.4]
  assign _T_1355 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@45864.4 package.scala 96:25:@45865.4]
  assign _T_1357 = io_rr ? _T_1355 : 1'h0; // @[implicits.scala 55:10:@45866.4]
  assign _T_1358 = _T_339 & _T_1357; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 584:194:@45867.4]
  assign x704_x466_D20 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@45852.4 package.scala 96:25:@45853.4]
  assign _T_1359 = _T_1358 & x704_x466_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 584:283:@45868.4]
  assign _T_1360 = _T_1359 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 584:291:@45869.4]
  assign x470 = x441 | x395; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 588:59:@45880.4]
  assign _T_1384 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@45913.4 package.scala 96:25:@45914.4]
  assign _T_1386 = io_rr ? _T_1384 : 1'h0; // @[implicits.scala 55:10:@45915.4]
  assign _T_1387 = _T_339 & _T_1386; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 599:194:@45916.4]
  assign x705_x471_D20 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@45901.4 package.scala 96:25:@45902.4]
  assign _T_1388 = _T_1387 & x705_x471_D20; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 599:283:@45917.4]
  assign _T_1389 = _T_1388 & x661_b330_D48; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 599:291:@45918.4]
  assign x531_number = x531_1_io_result; // @[Math.scala 723:22:@46572.4 Math.scala 724:14:@46573.4]
  assign x548_number = x548_1_io_result; // @[Math.scala 723:22:@46765.4 Math.scala 724:14:@46766.4]
  assign _T_1777 = {x531_number,x548_number}; // @[Cat.scala 30:58:@46774.4]
  assign x494_number = x494_1_io_result; // @[Math.scala 723:22:@46152.4 Math.scala 724:14:@46153.4]
  assign x514_number = x514_1_io_result; // @[Math.scala 723:22:@46381.4 Math.scala 724:14:@46382.4]
  assign _T_1778 = {x494_number,x514_number}; // @[Cat.scala 30:58:@46775.4]
  assign _T_1791 = RetimeWrapper_111_io_out; // @[package.scala 96:25:@46811.4 package.scala 96:25:@46812.4]
  assign _T_1793 = io_rr ? _T_1791 : 1'h0; // @[implicits.scala 55:10:@46813.4]
  assign x711_b330_D69 = RetimeWrapper_110_io_out; // @[package.scala 96:25:@46802.4 package.scala 96:25:@46803.4]
  assign _T_1794 = _T_1793 & x711_b330_D69; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 783:117:@46814.4]
  assign x710_b331_D69 = RetimeWrapper_109_io_out; // @[package.scala 96:25:@46793.4 package.scala 96:25:@46794.4]
  assign _T_1795 = _T_1794 & x710_b331_D69; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 783:123:@46815.4]
  assign x639_x339_D8_number = RetimeWrapper_2_io_out; // @[package.scala 96:25:@44035.4 package.scala 96:25:@44036.4]
  assign x640_x343_sum_D3_number = RetimeWrapper_3_io_out; // @[package.scala 96:25:@44044.4 package.scala 96:25:@44045.4]
  assign x641_x618_D24_number = RetimeWrapper_4_io_out; // @[package.scala 96:25:@44053.4 package.scala 96:25:@44054.4]
  assign x646_x347_D7_number = RetimeWrapper_10_io_out; // @[package.scala 96:25:@44169.4 package.scala 96:25:@44170.4]
  assign x647_x349_sum_D2_number = RetimeWrapper_11_io_out; // @[package.scala 96:25:@44178.4 package.scala 96:25:@44179.4]
  assign x650_x353_D7_number = RetimeWrapper_15_io_out; // @[package.scala 96:25:@44276.4 package.scala 96:25:@44277.4]
  assign x651_x355_sum_D2_number = RetimeWrapper_16_io_out; // @[package.scala 96:25:@44285.4 package.scala 96:25:@44286.4]
  assign x652_x361_sum_D2_number = RetimeWrapper_18_io_out; // @[package.scala 96:25:@44365.4 package.scala 96:25:@44366.4]
  assign x653_x359_D7_number = RetimeWrapper_19_io_out; // @[package.scala 96:25:@44374.4 package.scala 96:25:@44375.4]
  assign x658_x361_sum_D26_number = RetimeWrapper_27_io_out; // @[package.scala 96:25:@44478.4 package.scala 96:25:@44479.4]
  assign x659_x618_D48_number = RetimeWrapper_28_io_out; // @[package.scala 96:25:@44487.4 package.scala 96:25:@44488.4]
  assign x663_x359_D31_number = RetimeWrapper_32_io_out; // @[package.scala 96:25:@44523.4 package.scala 96:25:@44524.4]
  assign x666_x353_D31_number = RetimeWrapper_37_io_out; // @[package.scala 96:25:@44594.4 package.scala 96:25:@44595.4]
  assign x667_x355_sum_D26_number = RetimeWrapper_38_io_out; // @[package.scala 96:25:@44603.4 package.scala 96:25:@44604.4]
  assign x669_x347_D31_number = RetimeWrapper_42_io_out; // @[package.scala 96:25:@44665.4 package.scala 96:25:@44666.4]
  assign x670_x349_sum_D26_number = RetimeWrapper_43_io_out; // @[package.scala 96:25:@44674.4 package.scala 96:25:@44675.4]
  assign x673_x339_D32_number = RetimeWrapper_48_io_out; // @[package.scala 96:25:@44745.4 package.scala 96:25:@44746.4]
  assign x674_x343_sum_D27_number = RetimeWrapper_49_io_out; // @[package.scala 96:25:@44754.4 package.scala 96:25:@44755.4]
  assign x391_sum_number = x391_sum_1_io_result; // @[Math.scala 154:22:@44864.4 Math.scala 155:14:@44865.4]
  assign x677_x389_D5_number = RetimeWrapper_54_io_out; // @[package.scala 96:25:@44873.4 package.scala 96:25:@44874.4]
  assign x400_sum_number = x400_sum_1_io_result; // @[Math.scala 154:22:@44972.4 Math.scala 155:14:@44973.4]
  assign x680_x398_D5_number = RetimeWrapper_59_io_out; // @[package.scala 96:25:@44990.4 package.scala 96:25:@44991.4]
  assign x411_sum_number = x411_sum_1_io_result; // @[Math.scala 154:22:@45149.4 Math.scala 155:14:@45150.4]
  assign x683_x623_D20_number = RetimeWrapper_66_io_out; // @[package.scala 96:25:@45158.4 package.scala 96:25:@45159.4]
  assign x416_sum_number = x416_sum_1_io_result; // @[Math.scala 154:22:@45216.4 Math.scala 155:14:@45217.4]
  assign x421_sum_number = x421_sum_1_io_result; // @[Math.scala 154:22:@45274.4 Math.scala 155:14:@45275.4]
  assign x693_x426_sum_D1_number = RetimeWrapper_79_io_out; // @[package.scala 96:25:@45370.4 package.scala 96:25:@45371.4]
  assign x431_sum_number = x431_sum_1_io_result; // @[Math.scala 154:22:@45410.4 Math.scala 155:14:@45411.4]
  assign x436_sum_number = x436_sum_1_io_result; // @[Math.scala 154:22:@45459.4 Math.scala 155:14:@45460.4]
  assign x447_sum_number = x447_sum_1_io_result; // @[Math.scala 154:22:@45618.4 Math.scala 155:14:@45619.4]
  assign x697_x628_D20_number = RetimeWrapper_89_io_out; // @[package.scala 96:25:@45627.4 package.scala 96:25:@45628.4]
  assign x452_sum_number = x452_sum_1_io_result; // @[Math.scala 154:22:@45676.4 Math.scala 155:14:@45677.4]
  assign x457_sum_number = x457_sum_1_io_result; // @[Math.scala 154:22:@45725.4 Math.scala 155:14:@45726.4]
  assign x703_x462_sum_D1_number = RetimeWrapper_98_io_out; // @[package.scala 96:25:@45803.4 package.scala 96:25:@45804.4]
  assign x467_sum_number = x467_sum_1_io_result; // @[Math.scala 154:22:@45843.4 Math.scala 155:14:@45844.4]
  assign x472_sum_number = x472_sum_1_io_result; // @[Math.scala 154:22:@45892.4 Math.scala 155:14:@45893.4]
  assign io_in_x289_TREADY = _T_211 & _T_213; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 67:22:@43749.4 sm_x553_inr_Foreach_SAMPLER_BOX.scala 69:22:@43757.4]
  assign io_in_x290_TVALID = _T_1795 & io_sigsIn_backpressure; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 783:22:@46817.4]
  assign io_in_x290_TDATA = {{128'd0}, RetimeWrapper_108_io_out}; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 784:24:@46818.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@43727.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@43739.4]
  assign RetimeWrapper_clock = clock; // @[:@43760.4]
  assign RetimeWrapper_reset = reset; // @[:@43761.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@43763.4]
  assign RetimeWrapper_io_in = io_in_x289_TDATA[127:0]; // @[package.scala 94:16:@43762.4]
  assign x334_lb_0_clock = clock; // @[:@43770.4]
  assign x334_lb_0_reset = reset; // @[:@43771.4]
  assign x334_lb_0_io_rPort_17_banks_1 = x673_x339_D32_number[2:0]; // @[MemInterfaceType.scala 106:58:@45390.4]
  assign x334_lb_0_io_rPort_17_banks_0 = x683_x623_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@45389.4]
  assign x334_lb_0_io_rPort_17_ofs_0 = x693_x426_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@45391.4]
  assign x334_lb_0_io_rPort_17_en_0 = _T_1061 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@45393.4]
  assign x334_lb_0_io_rPort_17_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45392.4]
  assign x334_lb_0_io_rPort_16_banks_1 = x680_x398_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@45488.4]
  assign x334_lb_0_io_rPort_16_banks_0 = x683_x623_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@45487.4]
  assign x334_lb_0_io_rPort_16_ofs_0 = x436_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@45489.4]
  assign x334_lb_0_io_rPort_16_en_0 = _T_1119 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@45491.4]
  assign x334_lb_0_io_rPort_16_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45490.4]
  assign x334_lb_0_io_rPort_15_banks_1 = x666_x353_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@44623.4]
  assign x334_lb_0_io_rPort_15_banks_0 = x659_x618_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@44622.4]
  assign x334_lb_0_io_rPort_15_ofs_0 = x667_x355_sum_D26_number[8:0]; // @[MemInterfaceType.scala 107:54:@44624.4]
  assign x334_lb_0_io_rPort_15_en_0 = _T_613 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@44626.4]
  assign x334_lb_0_io_rPort_15_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@44625.4]
  assign x334_lb_0_io_rPort_14_banks_1 = x669_x347_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@45303.4]
  assign x334_lb_0_io_rPort_14_banks_0 = x683_x623_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@45302.4]
  assign x334_lb_0_io_rPort_14_ofs_0 = x421_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@45304.4]
  assign x334_lb_0_io_rPort_14_en_0 = _T_1018 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@45306.4]
  assign x334_lb_0_io_rPort_14_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45305.4]
  assign x334_lb_0_io_rPort_13_banks_1 = x677_x389_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@45439.4]
  assign x334_lb_0_io_rPort_13_banks_0 = x683_x623_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@45438.4]
  assign x334_lb_0_io_rPort_13_ofs_0 = x431_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@45440.4]
  assign x334_lb_0_io_rPort_13_en_0 = _T_1090 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@45442.4]
  assign x334_lb_0_io_rPort_13_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45441.4]
  assign x334_lb_0_io_rPort_12_banks_1 = x673_x339_D32_number[2:0]; // @[MemInterfaceType.scala 106:58:@44783.4]
  assign x334_lb_0_io_rPort_12_banks_0 = x659_x618_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@44782.4]
  assign x334_lb_0_io_rPort_12_ofs_0 = x674_x343_sum_D27_number[8:0]; // @[MemInterfaceType.scala 107:54:@44784.4]
  assign x334_lb_0_io_rPort_12_en_0 = _T_703 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@44786.4]
  assign x334_lb_0_io_rPort_12_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@44785.4]
  assign x334_lb_0_io_rPort_11_banks_1 = x669_x347_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@44703.4]
  assign x334_lb_0_io_rPort_11_banks_0 = x659_x618_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@44702.4]
  assign x334_lb_0_io_rPort_11_ofs_0 = x670_x349_sum_D26_number[8:0]; // @[MemInterfaceType.scala 107:54:@44704.4]
  assign x334_lb_0_io_rPort_11_en_0 = _T_658 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@44706.4]
  assign x334_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@44705.4]
  assign x334_lb_0_io_rPort_10_banks_1 = x680_x398_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@45010.4]
  assign x334_lb_0_io_rPort_10_banks_0 = x659_x618_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@45009.4]
  assign x334_lb_0_io_rPort_10_ofs_0 = x400_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@45011.4]
  assign x334_lb_0_io_rPort_10_en_0 = _T_834 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@45013.4]
  assign x334_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45012.4]
  assign x334_lb_0_io_rPort_9_banks_1 = x663_x359_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@44543.4]
  assign x334_lb_0_io_rPort_9_banks_0 = x659_x618_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@44542.4]
  assign x334_lb_0_io_rPort_9_ofs_0 = x658_x361_sum_D26_number[8:0]; // @[MemInterfaceType.scala 107:54:@44544.4]
  assign x334_lb_0_io_rPort_9_en_0 = _T_568 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@44546.4]
  assign x334_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@44545.4]
  assign x334_lb_0_io_rPort_8_banks_1 = x673_x339_D32_number[2:0]; // @[MemInterfaceType.scala 106:58:@45823.4]
  assign x334_lb_0_io_rPort_8_banks_0 = x697_x628_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@45822.4]
  assign x334_lb_0_io_rPort_8_ofs_0 = x703_x462_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@45824.4]
  assign x334_lb_0_io_rPort_8_en_0 = _T_1331 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@45826.4]
  assign x334_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45825.4]
  assign x334_lb_0_io_rPort_7_banks_1 = x669_x347_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@45754.4]
  assign x334_lb_0_io_rPort_7_banks_0 = x697_x628_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@45753.4]
  assign x334_lb_0_io_rPort_7_ofs_0 = x457_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@45755.4]
  assign x334_lb_0_io_rPort_7_en_0 = _T_1294 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@45757.4]
  assign x334_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45756.4]
  assign x334_lb_0_io_rPort_6_banks_1 = x680_x398_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@45921.4]
  assign x334_lb_0_io_rPort_6_banks_0 = x697_x628_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@45920.4]
  assign x334_lb_0_io_rPort_6_ofs_0 = x472_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@45922.4]
  assign x334_lb_0_io_rPort_6_en_0 = _T_1389 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@45924.4]
  assign x334_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45923.4]
  assign x334_lb_0_io_rPort_5_banks_1 = x663_x359_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@45187.4]
  assign x334_lb_0_io_rPort_5_banks_0 = x683_x623_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@45186.4]
  assign x334_lb_0_io_rPort_5_ofs_0 = x411_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@45188.4]
  assign x334_lb_0_io_rPort_5_en_0 = _T_954 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@45190.4]
  assign x334_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45189.4]
  assign x334_lb_0_io_rPort_4_banks_1 = x677_x389_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@44902.4]
  assign x334_lb_0_io_rPort_4_banks_0 = x659_x618_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@44901.4]
  assign x334_lb_0_io_rPort_4_ofs_0 = x391_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@44903.4]
  assign x334_lb_0_io_rPort_4_en_0 = _T_771 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@44905.4]
  assign x334_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@44904.4]
  assign x334_lb_0_io_rPort_3_banks_1 = x666_x353_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@45705.4]
  assign x334_lb_0_io_rPort_3_banks_0 = x697_x628_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@45704.4]
  assign x334_lb_0_io_rPort_3_ofs_0 = x452_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@45706.4]
  assign x334_lb_0_io_rPort_3_en_0 = _T_1265 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@45708.4]
  assign x334_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45707.4]
  assign x334_lb_0_io_rPort_2_banks_1 = x663_x359_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@45656.4]
  assign x334_lb_0_io_rPort_2_banks_0 = x697_x628_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@45655.4]
  assign x334_lb_0_io_rPort_2_ofs_0 = x447_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@45657.4]
  assign x334_lb_0_io_rPort_2_en_0 = _T_1236 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@45659.4]
  assign x334_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45658.4]
  assign x334_lb_0_io_rPort_1_banks_1 = x666_x353_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@45245.4]
  assign x334_lb_0_io_rPort_1_banks_0 = x683_x623_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@45244.4]
  assign x334_lb_0_io_rPort_1_ofs_0 = x416_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@45246.4]
  assign x334_lb_0_io_rPort_1_en_0 = _T_986 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@45248.4]
  assign x334_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45247.4]
  assign x334_lb_0_io_rPort_0_banks_1 = x677_x389_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@45872.4]
  assign x334_lb_0_io_rPort_0_banks_0 = x697_x628_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@45871.4]
  assign x334_lb_0_io_rPort_0_ofs_0 = x467_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@45873.4]
  assign x334_lb_0_io_rPort_0_en_0 = _T_1360 & x662_b331_D48; // @[MemInterfaceType.scala 110:79:@45875.4]
  assign x334_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@45874.4]
  assign x334_lb_0_io_wPort_3_banks_1 = x653_x359_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@44404.4]
  assign x334_lb_0_io_wPort_3_banks_0 = x641_x618_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@44403.4]
  assign x334_lb_0_io_wPort_3_ofs_0 = x652_x361_sum_D2_number[8:0]; // @[MemInterfaceType.scala 89:54:@44405.4]
  assign x334_lb_0_io_wPort_3_data_0 = RetimeWrapper_20_io_out; // @[MemInterfaceType.scala 90:56:@44406.4]
  assign x334_lb_0_io_wPort_3_en_0 = _T_497 & x643_b331_D24; // @[MemInterfaceType.scala 93:57:@44408.4]
  assign x334_lb_0_io_wPort_2_banks_1 = x650_x353_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@44306.4]
  assign x334_lb_0_io_wPort_2_banks_0 = x641_x618_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@44305.4]
  assign x334_lb_0_io_wPort_2_ofs_0 = x651_x355_sum_D2_number[8:0]; // @[MemInterfaceType.scala 89:54:@44307.4]
  assign x334_lb_0_io_wPort_2_data_0 = RetimeWrapper_14_io_out; // @[MemInterfaceType.scala 90:56:@44308.4]
  assign x334_lb_0_io_wPort_2_en_0 = _T_449 & x643_b331_D24; // @[MemInterfaceType.scala 93:57:@44310.4]
  assign x334_lb_0_io_wPort_1_banks_1 = x646_x347_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@44208.4]
  assign x334_lb_0_io_wPort_1_banks_0 = x641_x618_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@44207.4]
  assign x334_lb_0_io_wPort_1_ofs_0 = x647_x349_sum_D2_number[8:0]; // @[MemInterfaceType.scala 89:54:@44209.4]
  assign x334_lb_0_io_wPort_1_data_0 = RetimeWrapper_12_io_out; // @[MemInterfaceType.scala 90:56:@44210.4]
  assign x334_lb_0_io_wPort_1_en_0 = _T_401 & x643_b331_D24; // @[MemInterfaceType.scala 93:57:@44212.4]
  assign x334_lb_0_io_wPort_0_banks_1 = x639_x339_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@44101.4]
  assign x334_lb_0_io_wPort_0_banks_0 = x641_x618_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@44100.4]
  assign x334_lb_0_io_wPort_0_ofs_0 = x640_x343_sum_D3_number[8:0]; // @[MemInterfaceType.scala 89:54:@44102.4]
  assign x334_lb_0_io_wPort_0_data_0 = RetimeWrapper_7_io_out; // @[MemInterfaceType.scala 90:56:@44103.4]
  assign x334_lb_0_io_wPort_0_en_0 = _T_350 & x643_b331_D24; // @[MemInterfaceType.scala 93:57:@44105.4]
  assign x339_1_clock = clock; // @[:@43953.4]
  assign x339_1_io_a = __1_io_result; // @[Math.scala 367:17:@43955.4]
  assign x339_1_io_flow = io_in_x290_TREADY; // @[Math.scala 369:20:@43957.4]
  assign x621_sum_1_clock = clock; // @[:@43990.4]
  assign x621_sum_1_reset = reset; // @[:@43991.4]
  assign x621_sum_1_io_a = _T_300[31:0]; // @[Math.scala 151:17:@43992.4]
  assign x621_sum_1_io_b = _T_303[31:0]; // @[Math.scala 152:17:@43993.4]
  assign x621_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@43994.4]
  assign x342_div_1_clock = clock; // @[:@44002.4]
  assign x342_div_1_io_a = __1_io_result; // @[Math.scala 328:17:@44004.4]
  assign x342_div_1_io_flow = io_in_x290_TREADY; // @[Math.scala 330:20:@44006.4]
  assign RetimeWrapper_1_clock = clock; // @[:@44012.4]
  assign RetimeWrapper_1_reset = reset; // @[:@44013.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44015.4]
  assign RetimeWrapper_1_io_in = x621_sum_1_io_result; // @[package.scala 94:16:@44014.4]
  assign x343_sum_1_clock = clock; // @[:@44021.4]
  assign x343_sum_1_reset = reset; // @[:@44022.4]
  assign x343_sum_1_io_a = RetimeWrapper_1_io_out; // @[Math.scala 151:17:@44023.4]
  assign x343_sum_1_io_b = x342_div_1_io_result; // @[Math.scala 152:17:@44024.4]
  assign x343_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@44025.4]
  assign RetimeWrapper_2_clock = clock; // @[:@44031.4]
  assign RetimeWrapper_2_reset = reset; // @[:@44032.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44034.4]
  assign RetimeWrapper_2_io_in = x339_1_io_result; // @[package.scala 94:16:@44033.4]
  assign RetimeWrapper_3_clock = clock; // @[:@44040.4]
  assign RetimeWrapper_3_reset = reset; // @[:@44041.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44043.4]
  assign RetimeWrapper_3_io_in = x343_sum_1_io_result; // @[package.scala 94:16:@44042.4]
  assign RetimeWrapper_4_clock = clock; // @[:@44049.4]
  assign RetimeWrapper_4_reset = reset; // @[:@44050.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44052.4]
  assign RetimeWrapper_4_io_in = $unsigned(_T_263); // @[package.scala 94:16:@44051.4]
  assign RetimeWrapper_5_clock = clock; // @[:@44058.4]
  assign RetimeWrapper_5_reset = reset; // @[:@44059.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44061.4]
  assign RetimeWrapper_5_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@44060.4]
  assign RetimeWrapper_6_clock = clock; // @[:@44067.4]
  assign RetimeWrapper_6_reset = reset; // @[:@44068.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44070.4]
  assign RetimeWrapper_6_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@44069.4]
  assign RetimeWrapper_7_clock = clock; // @[:@44076.4]
  assign RetimeWrapper_7_reset = reset; // @[:@44077.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44079.4]
  assign RetimeWrapper_7_io_in = x637_x332_D1_0_number[31:0]; // @[package.scala 94:16:@44078.4]
  assign RetimeWrapper_8_clock = clock; // @[:@44087.4]
  assign RetimeWrapper_8_reset = reset; // @[:@44088.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44090.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44089.4]
  assign x345_rdcol_1_clock = clock; // @[:@44110.4]
  assign x345_rdcol_1_reset = reset; // @[:@44111.4]
  assign x345_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@44112.4]
  assign x345_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@44113.4]
  assign x345_rdcol_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@44114.4]
  assign x347_1_clock = clock; // @[:@44124.4]
  assign x347_1_io_a = x345_rdcol_1_io_result; // @[Math.scala 367:17:@44126.4]
  assign x347_1_io_flow = io_in_x290_TREADY; // @[Math.scala 369:20:@44128.4]
  assign x348_div_1_clock = clock; // @[:@44136.4]
  assign x348_div_1_io_a = x345_rdcol_1_io_result; // @[Math.scala 328:17:@44138.4]
  assign x348_div_1_io_flow = io_in_x290_TREADY; // @[Math.scala 330:20:@44140.4]
  assign RetimeWrapper_9_clock = clock; // @[:@44146.4]
  assign RetimeWrapper_9_reset = reset; // @[:@44147.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44149.4]
  assign RetimeWrapper_9_io_in = x621_sum_1_io_result; // @[package.scala 94:16:@44148.4]
  assign x349_sum_1_clock = clock; // @[:@44155.4]
  assign x349_sum_1_reset = reset; // @[:@44156.4]
  assign x349_sum_1_io_a = RetimeWrapper_9_io_out; // @[Math.scala 151:17:@44157.4]
  assign x349_sum_1_io_b = x348_div_1_io_result; // @[Math.scala 152:17:@44158.4]
  assign x349_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@44159.4]
  assign RetimeWrapper_10_clock = clock; // @[:@44165.4]
  assign RetimeWrapper_10_reset = reset; // @[:@44166.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44168.4]
  assign RetimeWrapper_10_io_in = x347_1_io_result; // @[package.scala 94:16:@44167.4]
  assign RetimeWrapper_11_clock = clock; // @[:@44174.4]
  assign RetimeWrapper_11_reset = reset; // @[:@44175.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44177.4]
  assign RetimeWrapper_11_io_in = x349_sum_1_io_result; // @[package.scala 94:16:@44176.4]
  assign RetimeWrapper_12_clock = clock; // @[:@44183.4]
  assign RetimeWrapper_12_reset = reset; // @[:@44184.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44186.4]
  assign RetimeWrapper_12_io_in = x637_x332_D1_0_number[63:32]; // @[package.scala 94:16:@44185.4]
  assign RetimeWrapper_13_clock = clock; // @[:@44194.4]
  assign RetimeWrapper_13_reset = reset; // @[:@44195.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44197.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44196.4]
  assign x351_rdcol_1_clock = clock; // @[:@44217.4]
  assign x351_rdcol_1_reset = reset; // @[:@44218.4]
  assign x351_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@44219.4]
  assign x351_rdcol_1_io_b = 32'h2; // @[Math.scala 152:17:@44220.4]
  assign x351_rdcol_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@44221.4]
  assign x353_1_clock = clock; // @[:@44231.4]
  assign x353_1_io_a = x351_rdcol_1_io_result; // @[Math.scala 367:17:@44233.4]
  assign x353_1_io_flow = io_in_x290_TREADY; // @[Math.scala 369:20:@44235.4]
  assign x354_div_1_clock = clock; // @[:@44243.4]
  assign x354_div_1_io_a = x351_rdcol_1_io_result; // @[Math.scala 328:17:@44245.4]
  assign x354_div_1_io_flow = io_in_x290_TREADY; // @[Math.scala 330:20:@44247.4]
  assign x355_sum_1_clock = clock; // @[:@44253.4]
  assign x355_sum_1_reset = reset; // @[:@44254.4]
  assign x355_sum_1_io_a = RetimeWrapper_9_io_out; // @[Math.scala 151:17:@44255.4]
  assign x355_sum_1_io_b = x354_div_1_io_result; // @[Math.scala 152:17:@44256.4]
  assign x355_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@44257.4]
  assign RetimeWrapper_14_clock = clock; // @[:@44263.4]
  assign RetimeWrapper_14_reset = reset; // @[:@44264.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44266.4]
  assign RetimeWrapper_14_io_in = x637_x332_D1_0_number[95:64]; // @[package.scala 94:16:@44265.4]
  assign RetimeWrapper_15_clock = clock; // @[:@44272.4]
  assign RetimeWrapper_15_reset = reset; // @[:@44273.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44275.4]
  assign RetimeWrapper_15_io_in = x353_1_io_result; // @[package.scala 94:16:@44274.4]
  assign RetimeWrapper_16_clock = clock; // @[:@44281.4]
  assign RetimeWrapper_16_reset = reset; // @[:@44282.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44284.4]
  assign RetimeWrapper_16_io_in = x355_sum_1_io_result; // @[package.scala 94:16:@44283.4]
  assign RetimeWrapper_17_clock = clock; // @[:@44292.4]
  assign RetimeWrapper_17_reset = reset; // @[:@44293.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44295.4]
  assign RetimeWrapper_17_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44294.4]
  assign x357_rdcol_1_clock = clock; // @[:@44315.4]
  assign x357_rdcol_1_reset = reset; // @[:@44316.4]
  assign x357_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@44317.4]
  assign x357_rdcol_1_io_b = 32'h3; // @[Math.scala 152:17:@44318.4]
  assign x357_rdcol_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@44319.4]
  assign x359_1_clock = clock; // @[:@44329.4]
  assign x359_1_io_a = x357_rdcol_1_io_result; // @[Math.scala 367:17:@44331.4]
  assign x359_1_io_flow = io_in_x290_TREADY; // @[Math.scala 369:20:@44333.4]
  assign x360_div_1_clock = clock; // @[:@44341.4]
  assign x360_div_1_io_a = x357_rdcol_1_io_result; // @[Math.scala 328:17:@44343.4]
  assign x360_div_1_io_flow = io_in_x290_TREADY; // @[Math.scala 330:20:@44345.4]
  assign x361_sum_1_clock = clock; // @[:@44351.4]
  assign x361_sum_1_reset = reset; // @[:@44352.4]
  assign x361_sum_1_io_a = RetimeWrapper_9_io_out; // @[Math.scala 151:17:@44353.4]
  assign x361_sum_1_io_b = x360_div_1_io_result; // @[Math.scala 152:17:@44354.4]
  assign x361_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@44355.4]
  assign RetimeWrapper_18_clock = clock; // @[:@44361.4]
  assign RetimeWrapper_18_reset = reset; // @[:@44362.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44364.4]
  assign RetimeWrapper_18_io_in = x361_sum_1_io_result; // @[package.scala 94:16:@44363.4]
  assign RetimeWrapper_19_clock = clock; // @[:@44370.4]
  assign RetimeWrapper_19_reset = reset; // @[:@44371.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44373.4]
  assign RetimeWrapper_19_io_in = x359_1_io_result; // @[package.scala 94:16:@44372.4]
  assign RetimeWrapper_20_clock = clock; // @[:@44379.4]
  assign RetimeWrapper_20_reset = reset; // @[:@44380.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44382.4]
  assign RetimeWrapper_20_io_in = x637_x332_D1_0_number[127:96]; // @[package.scala 94:16:@44381.4]
  assign RetimeWrapper_21_clock = clock; // @[:@44390.4]
  assign RetimeWrapper_21_reset = reset; // @[:@44391.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44393.4]
  assign RetimeWrapper_21_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44392.4]
  assign RetimeWrapper_22_clock = clock; // @[:@44411.4]
  assign RetimeWrapper_22_reset = reset; // @[:@44412.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44414.4]
  assign RetimeWrapper_22_io_in = __io_result; // @[package.scala 94:16:@44413.4]
  assign RetimeWrapper_23_clock = clock; // @[:@44427.4]
  assign RetimeWrapper_23_reset = reset; // @[:@44428.4]
  assign RetimeWrapper_23_io_flow = io_in_x290_TREADY; // @[package.scala 95:18:@44430.4]
  assign RetimeWrapper_23_io_in = $signed(_T_509) < $signed(32'sh0); // @[package.scala 94:16:@44429.4]
  assign RetimeWrapper_24_clock = clock; // @[:@44436.4]
  assign RetimeWrapper_24_reset = reset; // @[:@44437.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44439.4]
  assign RetimeWrapper_24_io_in = x357_rdcol_1_io_result; // @[package.scala 94:16:@44438.4]
  assign RetimeWrapper_25_clock = clock; // @[:@44450.4]
  assign RetimeWrapper_25_reset = reset; // @[:@44451.4]
  assign RetimeWrapper_25_io_flow = io_in_x290_TREADY; // @[package.scala 95:18:@44453.4]
  assign RetimeWrapper_25_io_in = $signed(_T_522) < $signed(32'sh0); // @[package.scala 94:16:@44452.4]
  assign RetimeWrapper_26_clock = clock; // @[:@44459.4]
  assign RetimeWrapper_26_reset = reset; // @[:@44460.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44462.4]
  assign RetimeWrapper_26_io_in = RetimeWrapper_23_io_out; // @[package.scala 94:16:@44461.4]
  assign RetimeWrapper_27_clock = clock; // @[:@44474.4]
  assign RetimeWrapper_27_reset = reset; // @[:@44475.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44477.4]
  assign RetimeWrapper_27_io_in = x361_sum_1_io_result; // @[package.scala 94:16:@44476.4]
  assign RetimeWrapper_28_clock = clock; // @[:@44483.4]
  assign RetimeWrapper_28_reset = reset; // @[:@44484.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44486.4]
  assign RetimeWrapper_28_io_in = $unsigned(_T_263); // @[package.scala 94:16:@44485.4]
  assign RetimeWrapper_29_clock = clock; // @[:@44492.4]
  assign RetimeWrapper_29_reset = reset; // @[:@44493.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44495.4]
  assign RetimeWrapper_29_io_in = ~ x366; // @[package.scala 94:16:@44494.4]
  assign RetimeWrapper_30_clock = clock; // @[:@44501.4]
  assign RetimeWrapper_30_reset = reset; // @[:@44502.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44504.4]
  assign RetimeWrapper_30_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@44503.4]
  assign RetimeWrapper_31_clock = clock; // @[:@44510.4]
  assign RetimeWrapper_31_reset = reset; // @[:@44511.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44513.4]
  assign RetimeWrapper_31_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@44512.4]
  assign RetimeWrapper_32_clock = clock; // @[:@44519.4]
  assign RetimeWrapper_32_reset = reset; // @[:@44520.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44522.4]
  assign RetimeWrapper_32_io_in = x359_1_io_result; // @[package.scala 94:16:@44521.4]
  assign RetimeWrapper_33_clock = clock; // @[:@44531.4]
  assign RetimeWrapper_33_reset = reset; // @[:@44532.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44534.4]
  assign RetimeWrapper_33_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44533.4]
  assign RetimeWrapper_34_clock = clock; // @[:@44552.4]
  assign RetimeWrapper_34_reset = reset; // @[:@44553.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44555.4]
  assign RetimeWrapper_34_io_in = x351_rdcol_1_io_result; // @[package.scala 94:16:@44554.4]
  assign RetimeWrapper_35_clock = clock; // @[:@44566.4]
  assign RetimeWrapper_35_reset = reset; // @[:@44567.4]
  assign RetimeWrapper_35_io_flow = io_in_x290_TREADY; // @[package.scala 95:18:@44569.4]
  assign RetimeWrapper_35_io_in = $signed(_T_579) < $signed(32'sh0); // @[package.scala 94:16:@44568.4]
  assign RetimeWrapper_36_clock = clock; // @[:@44581.4]
  assign RetimeWrapper_36_reset = reset; // @[:@44582.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44584.4]
  assign RetimeWrapper_36_io_in = ~ x371; // @[package.scala 94:16:@44583.4]
  assign RetimeWrapper_37_clock = clock; // @[:@44590.4]
  assign RetimeWrapper_37_reset = reset; // @[:@44591.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44593.4]
  assign RetimeWrapper_37_io_in = x353_1_io_result; // @[package.scala 94:16:@44592.4]
  assign RetimeWrapper_38_clock = clock; // @[:@44599.4]
  assign RetimeWrapper_38_reset = reset; // @[:@44600.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44602.4]
  assign RetimeWrapper_38_io_in = x355_sum_1_io_result; // @[package.scala 94:16:@44601.4]
  assign RetimeWrapper_39_clock = clock; // @[:@44611.4]
  assign RetimeWrapper_39_reset = reset; // @[:@44612.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44614.4]
  assign RetimeWrapper_39_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44613.4]
  assign RetimeWrapper_40_clock = clock; // @[:@44632.4]
  assign RetimeWrapper_40_reset = reset; // @[:@44633.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44635.4]
  assign RetimeWrapper_40_io_in = x345_rdcol_1_io_result; // @[package.scala 94:16:@44634.4]
  assign RetimeWrapper_41_clock = clock; // @[:@44646.4]
  assign RetimeWrapper_41_reset = reset; // @[:@44647.4]
  assign RetimeWrapper_41_io_flow = io_in_x290_TREADY; // @[package.scala 95:18:@44649.4]
  assign RetimeWrapper_41_io_in = $signed(_T_624) < $signed(32'sh0); // @[package.scala 94:16:@44648.4]
  assign RetimeWrapper_42_clock = clock; // @[:@44661.4]
  assign RetimeWrapper_42_reset = reset; // @[:@44662.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44664.4]
  assign RetimeWrapper_42_io_in = x347_1_io_result; // @[package.scala 94:16:@44663.4]
  assign RetimeWrapper_43_clock = clock; // @[:@44670.4]
  assign RetimeWrapper_43_reset = reset; // @[:@44671.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44673.4]
  assign RetimeWrapper_43_io_in = x349_sum_1_io_result; // @[package.scala 94:16:@44672.4]
  assign RetimeWrapper_44_clock = clock; // @[:@44679.4]
  assign RetimeWrapper_44_reset = reset; // @[:@44680.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44682.4]
  assign RetimeWrapper_44_io_in = ~ x376; // @[package.scala 94:16:@44681.4]
  assign RetimeWrapper_45_clock = clock; // @[:@44691.4]
  assign RetimeWrapper_45_reset = reset; // @[:@44692.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44694.4]
  assign RetimeWrapper_45_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44693.4]
  assign RetimeWrapper_46_clock = clock; // @[:@44712.4]
  assign RetimeWrapper_46_reset = reset; // @[:@44713.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44715.4]
  assign RetimeWrapper_46_io_in = __1_io_result; // @[package.scala 94:16:@44714.4]
  assign RetimeWrapper_47_clock = clock; // @[:@44726.4]
  assign RetimeWrapper_47_reset = reset; // @[:@44727.4]
  assign RetimeWrapper_47_io_flow = io_in_x290_TREADY; // @[package.scala 95:18:@44729.4]
  assign RetimeWrapper_47_io_in = $signed(_T_669) < $signed(32'sh0); // @[package.scala 94:16:@44728.4]
  assign RetimeWrapper_48_clock = clock; // @[:@44741.4]
  assign RetimeWrapper_48_reset = reset; // @[:@44742.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44744.4]
  assign RetimeWrapper_48_io_in = x339_1_io_result; // @[package.scala 94:16:@44743.4]
  assign RetimeWrapper_49_clock = clock; // @[:@44750.4]
  assign RetimeWrapper_49_reset = reset; // @[:@44751.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44753.4]
  assign RetimeWrapper_49_io_in = x343_sum_1_io_result; // @[package.scala 94:16:@44752.4]
  assign RetimeWrapper_50_clock = clock; // @[:@44759.4]
  assign RetimeWrapper_50_reset = reset; // @[:@44760.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44762.4]
  assign RetimeWrapper_50_io_in = ~ x381; // @[package.scala 94:16:@44761.4]
  assign RetimeWrapper_51_clock = clock; // @[:@44771.4]
  assign RetimeWrapper_51_reset = reset; // @[:@44772.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44774.4]
  assign RetimeWrapper_51_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44773.4]
  assign x385_rdcol_1_clock = clock; // @[:@44794.4]
  assign x385_rdcol_1_reset = reset; // @[:@44795.4]
  assign x385_rdcol_1_io_a = RetimeWrapper_46_io_out; // @[Math.scala 151:17:@44796.4]
  assign x385_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@44797.4]
  assign x385_rdcol_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@44798.4]
  assign RetimeWrapper_52_clock = clock; // @[:@44809.4]
  assign RetimeWrapper_52_reset = reset; // @[:@44810.4]
  assign RetimeWrapper_52_io_flow = io_in_x290_TREADY; // @[package.scala 95:18:@44812.4]
  assign RetimeWrapper_52_io_in = $signed(_T_718) < $signed(32'sh0); // @[package.scala 94:16:@44811.4]
  assign x389_1_clock = clock; // @[:@44828.4]
  assign x389_1_io_a = x385_rdcol_1_io_result; // @[Math.scala 367:17:@44830.4]
  assign x389_1_io_flow = io_in_x290_TREADY; // @[Math.scala 369:20:@44832.4]
  assign x390_div_1_clock = clock; // @[:@44840.4]
  assign x390_div_1_io_a = x385_rdcol_1_io_result; // @[Math.scala 328:17:@44842.4]
  assign x390_div_1_io_flow = io_in_x290_TREADY; // @[Math.scala 330:20:@44844.4]
  assign RetimeWrapper_53_clock = clock; // @[:@44850.4]
  assign RetimeWrapper_53_reset = reset; // @[:@44851.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44853.4]
  assign RetimeWrapper_53_io_in = x621_sum_1_io_result; // @[package.scala 94:16:@44852.4]
  assign x391_sum_1_clock = clock; // @[:@44859.4]
  assign x391_sum_1_reset = reset; // @[:@44860.4]
  assign x391_sum_1_io_a = RetimeWrapper_53_io_out; // @[Math.scala 151:17:@44861.4]
  assign x391_sum_1_io_b = x390_div_1_io_result; // @[Math.scala 152:17:@44862.4]
  assign x391_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@44863.4]
  assign RetimeWrapper_54_clock = clock; // @[:@44869.4]
  assign RetimeWrapper_54_reset = reset; // @[:@44870.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44872.4]
  assign RetimeWrapper_54_io_in = x389_1_io_result; // @[package.scala 94:16:@44871.4]
  assign RetimeWrapper_55_clock = clock; // @[:@44878.4]
  assign RetimeWrapper_55_reset = reset; // @[:@44879.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44881.4]
  assign RetimeWrapper_55_io_in = ~ x387; // @[package.scala 94:16:@44880.4]
  assign RetimeWrapper_56_clock = clock; // @[:@44890.4]
  assign RetimeWrapper_56_reset = reset; // @[:@44891.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44893.4]
  assign RetimeWrapper_56_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44892.4]
  assign x394_rdcol_1_clock = clock; // @[:@44913.4]
  assign x394_rdcol_1_reset = reset; // @[:@44914.4]
  assign x394_rdcol_1_io_a = RetimeWrapper_46_io_out; // @[Math.scala 151:17:@44915.4]
  assign x394_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@44916.4]
  assign x394_rdcol_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@44917.4]
  assign RetimeWrapper_57_clock = clock; // @[:@44928.4]
  assign RetimeWrapper_57_reset = reset; // @[:@44929.4]
  assign RetimeWrapper_57_io_flow = io_in_x290_TREADY; // @[package.scala 95:18:@44931.4]
  assign RetimeWrapper_57_io_in = $signed(_T_786) < $signed(32'sh0); // @[package.scala 94:16:@44930.4]
  assign x398_1_clock = clock; // @[:@44945.4]
  assign x398_1_io_a = x394_rdcol_1_io_result; // @[Math.scala 367:17:@44947.4]
  assign x398_1_io_flow = io_in_x290_TREADY; // @[Math.scala 369:20:@44949.4]
  assign x399_div_1_clock = clock; // @[:@44957.4]
  assign x399_div_1_io_a = x394_rdcol_1_io_result; // @[Math.scala 328:17:@44959.4]
  assign x399_div_1_io_flow = io_in_x290_TREADY; // @[Math.scala 330:20:@44961.4]
  assign x400_sum_1_clock = clock; // @[:@44967.4]
  assign x400_sum_1_reset = reset; // @[:@44968.4]
  assign x400_sum_1_io_a = RetimeWrapper_53_io_out; // @[Math.scala 151:17:@44969.4]
  assign x400_sum_1_io_b = x399_div_1_io_result; // @[Math.scala 152:17:@44970.4]
  assign x400_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@44971.4]
  assign RetimeWrapper_58_clock = clock; // @[:@44977.4]
  assign RetimeWrapper_58_reset = reset; // @[:@44978.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44980.4]
  assign RetimeWrapper_58_io_in = ~ x396; // @[package.scala 94:16:@44979.4]
  assign RetimeWrapper_59_clock = clock; // @[:@44986.4]
  assign RetimeWrapper_59_reset = reset; // @[:@44987.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@44989.4]
  assign RetimeWrapper_59_io_in = x398_1_io_result; // @[package.scala 94:16:@44988.4]
  assign RetimeWrapper_60_clock = clock; // @[:@44998.4]
  assign RetimeWrapper_60_reset = reset; // @[:@44999.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45001.4]
  assign RetimeWrapper_60_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45000.4]
  assign x403_rdrow_1_clock = clock; // @[:@45021.4]
  assign x403_rdrow_1_reset = reset; // @[:@45022.4]
  assign x403_rdrow_1_io_a = RetimeWrapper_22_io_out; // @[Math.scala 192:17:@45023.4]
  assign x403_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@45024.4]
  assign x403_rdrow_1_io_flow = io_in_x290_TREADY; // @[Math.scala 194:20:@45025.4]
  assign RetimeWrapper_61_clock = clock; // @[:@45047.4]
  assign RetimeWrapper_61_reset = reset; // @[:@45048.4]
  assign RetimeWrapper_61_io_flow = io_in_x290_TREADY; // @[package.scala 95:18:@45050.4]
  assign RetimeWrapper_61_io_in = $signed(_T_851) < $signed(32'sh0); // @[package.scala 94:16:@45049.4]
  assign RetimeWrapper_62_clock = clock; // @[:@45069.4]
  assign RetimeWrapper_62_reset = reset; // @[:@45070.4]
  assign RetimeWrapper_62_io_flow = io_in_x290_TREADY; // @[package.scala 95:18:@45073.4]
  assign RetimeWrapper_62_io_in = $unsigned(_T_880); // @[package.scala 94:16:@45072.4]
  assign RetimeWrapper_63_clock = clock; // @[:@45095.4]
  assign RetimeWrapper_63_reset = reset; // @[:@45096.4]
  assign RetimeWrapper_63_io_flow = io_in_x290_TREADY; // @[package.scala 95:18:@45098.4]
  assign RetimeWrapper_63_io_in = {_T_892,_T_893}; // @[package.scala 94:16:@45097.4]
  assign x626_sum_1_clock = clock; // @[:@45116.4]
  assign x626_sum_1_reset = reset; // @[:@45117.4]
  assign x626_sum_1_io_a = _T_916[31:0]; // @[Math.scala 151:17:@45118.4]
  assign x626_sum_1_io_b = _T_919[31:0]; // @[Math.scala 152:17:@45119.4]
  assign x626_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@45120.4]
  assign RetimeWrapper_64_clock = clock; // @[:@45126.4]
  assign RetimeWrapper_64_reset = reset; // @[:@45127.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45129.4]
  assign RetimeWrapper_64_io_in = x626_sum_1_io_result; // @[package.scala 94:16:@45128.4]
  assign RetimeWrapper_65_clock = clock; // @[:@45135.4]
  assign RetimeWrapper_65_reset = reset; // @[:@45136.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45138.4]
  assign RetimeWrapper_65_io_in = x360_div_1_io_result; // @[package.scala 94:16:@45137.4]
  assign x411_sum_1_clock = clock; // @[:@45144.4]
  assign x411_sum_1_reset = reset; // @[:@45145.4]
  assign x411_sum_1_io_a = RetimeWrapper_64_io_out; // @[Math.scala 151:17:@45146.4]
  assign x411_sum_1_io_b = RetimeWrapper_65_io_out; // @[Math.scala 152:17:@45147.4]
  assign x411_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@45148.4]
  assign RetimeWrapper_66_clock = clock; // @[:@45154.4]
  assign RetimeWrapper_66_reset = reset; // @[:@45155.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45157.4]
  assign RetimeWrapper_66_io_in = $unsigned(_T_884); // @[package.scala 94:16:@45156.4]
  assign RetimeWrapper_67_clock = clock; // @[:@45163.4]
  assign RetimeWrapper_67_reset = reset; // @[:@45164.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45166.4]
  assign RetimeWrapper_67_io_in = ~ x406; // @[package.scala 94:16:@45165.4]
  assign RetimeWrapper_68_clock = clock; // @[:@45175.4]
  assign RetimeWrapper_68_reset = reset; // @[:@45176.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45178.4]
  assign RetimeWrapper_68_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45177.4]
  assign RetimeWrapper_69_clock = clock; // @[:@45202.4]
  assign RetimeWrapper_69_reset = reset; // @[:@45203.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45205.4]
  assign RetimeWrapper_69_io_in = x354_div_1_io_result; // @[package.scala 94:16:@45204.4]
  assign x416_sum_1_clock = clock; // @[:@45211.4]
  assign x416_sum_1_reset = reset; // @[:@45212.4]
  assign x416_sum_1_io_a = RetimeWrapper_64_io_out; // @[Math.scala 151:17:@45213.4]
  assign x416_sum_1_io_b = RetimeWrapper_69_io_out; // @[Math.scala 152:17:@45214.4]
  assign x416_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@45215.4]
  assign RetimeWrapper_70_clock = clock; // @[:@45221.4]
  assign RetimeWrapper_70_reset = reset; // @[:@45222.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45224.4]
  assign RetimeWrapper_70_io_in = ~ x414; // @[package.scala 94:16:@45223.4]
  assign RetimeWrapper_71_clock = clock; // @[:@45233.4]
  assign RetimeWrapper_71_reset = reset; // @[:@45234.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45236.4]
  assign RetimeWrapper_71_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45235.4]
  assign RetimeWrapper_72_clock = clock; // @[:@45260.4]
  assign RetimeWrapper_72_reset = reset; // @[:@45261.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45263.4]
  assign RetimeWrapper_72_io_in = x348_div_1_io_result; // @[package.scala 94:16:@45262.4]
  assign x421_sum_1_clock = clock; // @[:@45269.4]
  assign x421_sum_1_reset = reset; // @[:@45270.4]
  assign x421_sum_1_io_a = RetimeWrapper_64_io_out; // @[Math.scala 151:17:@45271.4]
  assign x421_sum_1_io_b = RetimeWrapper_72_io_out; // @[Math.scala 152:17:@45272.4]
  assign x421_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@45273.4]
  assign RetimeWrapper_73_clock = clock; // @[:@45279.4]
  assign RetimeWrapper_73_reset = reset; // @[:@45280.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45282.4]
  assign RetimeWrapper_73_io_in = ~ x419; // @[package.scala 94:16:@45281.4]
  assign RetimeWrapper_74_clock = clock; // @[:@45291.4]
  assign RetimeWrapper_74_reset = reset; // @[:@45292.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45294.4]
  assign RetimeWrapper_74_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45293.4]
  assign RetimeWrapper_75_clock = clock; // @[:@45312.4]
  assign RetimeWrapper_75_reset = reset; // @[:@45313.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45315.4]
  assign RetimeWrapper_75_io_in = RetimeWrapper_47_io_out; // @[package.scala 94:16:@45314.4]
  assign RetimeWrapper_76_clock = clock; // @[:@45327.4]
  assign RetimeWrapper_76_reset = reset; // @[:@45328.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45330.4]
  assign RetimeWrapper_76_io_in = x342_div_1_io_result; // @[package.scala 94:16:@45329.4]
  assign RetimeWrapper_77_clock = clock; // @[:@45336.4]
  assign RetimeWrapper_77_reset = reset; // @[:@45337.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45339.4]
  assign RetimeWrapper_77_io_in = x626_sum_1_io_result; // @[package.scala 94:16:@45338.4]
  assign x426_sum_1_clock = clock; // @[:@45347.4]
  assign x426_sum_1_reset = reset; // @[:@45348.4]
  assign x426_sum_1_io_a = RetimeWrapper_77_io_out; // @[Math.scala 151:17:@45349.4]
  assign x426_sum_1_io_b = RetimeWrapper_76_io_out; // @[Math.scala 152:17:@45350.4]
  assign x426_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@45351.4]
  assign RetimeWrapper_78_clock = clock; // @[:@45357.4]
  assign RetimeWrapper_78_reset = reset; // @[:@45358.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45360.4]
  assign RetimeWrapper_78_io_in = ~ x424; // @[package.scala 94:16:@45359.4]
  assign RetimeWrapper_79_clock = clock; // @[:@45366.4]
  assign RetimeWrapper_79_reset = reset; // @[:@45367.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45369.4]
  assign RetimeWrapper_79_io_in = x426_sum_1_io_result; // @[package.scala 94:16:@45368.4]
  assign RetimeWrapper_80_clock = clock; // @[:@45378.4]
  assign RetimeWrapper_80_reset = reset; // @[:@45379.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45381.4]
  assign RetimeWrapper_80_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45380.4]
  assign x431_sum_1_clock = clock; // @[:@45405.4]
  assign x431_sum_1_reset = reset; // @[:@45406.4]
  assign x431_sum_1_io_a = RetimeWrapper_64_io_out; // @[Math.scala 151:17:@45407.4]
  assign x431_sum_1_io_b = x390_div_1_io_result; // @[Math.scala 152:17:@45408.4]
  assign x431_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@45409.4]
  assign RetimeWrapper_81_clock = clock; // @[:@45415.4]
  assign RetimeWrapper_81_reset = reset; // @[:@45416.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45418.4]
  assign RetimeWrapper_81_io_in = ~ x429; // @[package.scala 94:16:@45417.4]
  assign RetimeWrapper_82_clock = clock; // @[:@45427.4]
  assign RetimeWrapper_82_reset = reset; // @[:@45428.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45430.4]
  assign RetimeWrapper_82_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45429.4]
  assign x436_sum_1_clock = clock; // @[:@45454.4]
  assign x436_sum_1_reset = reset; // @[:@45455.4]
  assign x436_sum_1_io_a = RetimeWrapper_64_io_out; // @[Math.scala 151:17:@45456.4]
  assign x436_sum_1_io_b = x399_div_1_io_result; // @[Math.scala 152:17:@45457.4]
  assign x436_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@45458.4]
  assign RetimeWrapper_83_clock = clock; // @[:@45464.4]
  assign RetimeWrapper_83_reset = reset; // @[:@45465.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45467.4]
  assign RetimeWrapper_83_io_in = ~ x434; // @[package.scala 94:16:@45466.4]
  assign RetimeWrapper_84_clock = clock; // @[:@45476.4]
  assign RetimeWrapper_84_reset = reset; // @[:@45477.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45479.4]
  assign RetimeWrapper_84_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45478.4]
  assign x439_rdrow_1_clock = clock; // @[:@45499.4]
  assign x439_rdrow_1_reset = reset; // @[:@45500.4]
  assign x439_rdrow_1_io_a = RetimeWrapper_22_io_out; // @[Math.scala 192:17:@45501.4]
  assign x439_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@45502.4]
  assign x439_rdrow_1_io_flow = io_in_x290_TREADY; // @[Math.scala 194:20:@45503.4]
  assign RetimeWrapper_85_clock = clock; // @[:@45525.4]
  assign RetimeWrapper_85_reset = reset; // @[:@45526.4]
  assign RetimeWrapper_85_io_flow = io_in_x290_TREADY; // @[package.scala 95:18:@45528.4]
  assign RetimeWrapper_85_io_in = $signed(_T_1136) < $signed(32'sh0); // @[package.scala 94:16:@45527.4]
  assign RetimeWrapper_86_clock = clock; // @[:@45547.4]
  assign RetimeWrapper_86_reset = reset; // @[:@45548.4]
  assign RetimeWrapper_86_io_flow = io_in_x290_TREADY; // @[package.scala 95:18:@45551.4]
  assign RetimeWrapper_86_io_in = $unsigned(_T_1165); // @[package.scala 94:16:@45550.4]
  assign RetimeWrapper_87_clock = clock; // @[:@45573.4]
  assign RetimeWrapper_87_reset = reset; // @[:@45574.4]
  assign RetimeWrapper_87_io_flow = io_in_x290_TREADY; // @[package.scala 95:18:@45576.4]
  assign RetimeWrapper_87_io_in = {_T_1177,_T_1178}; // @[package.scala 94:16:@45575.4]
  assign x631_sum_1_clock = clock; // @[:@45594.4]
  assign x631_sum_1_reset = reset; // @[:@45595.4]
  assign x631_sum_1_io_a = _T_1201[31:0]; // @[Math.scala 151:17:@45596.4]
  assign x631_sum_1_io_b = _T_1204[31:0]; // @[Math.scala 152:17:@45597.4]
  assign x631_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@45598.4]
  assign RetimeWrapper_88_clock = clock; // @[:@45604.4]
  assign RetimeWrapper_88_reset = reset; // @[:@45605.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45607.4]
  assign RetimeWrapper_88_io_in = x631_sum_1_io_result; // @[package.scala 94:16:@45606.4]
  assign x447_sum_1_clock = clock; // @[:@45613.4]
  assign x447_sum_1_reset = reset; // @[:@45614.4]
  assign x447_sum_1_io_a = RetimeWrapper_88_io_out; // @[Math.scala 151:17:@45615.4]
  assign x447_sum_1_io_b = RetimeWrapper_65_io_out; // @[Math.scala 152:17:@45616.4]
  assign x447_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@45617.4]
  assign RetimeWrapper_89_clock = clock; // @[:@45623.4]
  assign RetimeWrapper_89_reset = reset; // @[:@45624.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45626.4]
  assign RetimeWrapper_89_io_in = $unsigned(_T_1169); // @[package.scala 94:16:@45625.4]
  assign RetimeWrapper_90_clock = clock; // @[:@45632.4]
  assign RetimeWrapper_90_reset = reset; // @[:@45633.4]
  assign RetimeWrapper_90_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45635.4]
  assign RetimeWrapper_90_io_in = ~ x442; // @[package.scala 94:16:@45634.4]
  assign RetimeWrapper_91_clock = clock; // @[:@45644.4]
  assign RetimeWrapper_91_reset = reset; // @[:@45645.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45647.4]
  assign RetimeWrapper_91_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45646.4]
  assign x452_sum_1_clock = clock; // @[:@45671.4]
  assign x452_sum_1_reset = reset; // @[:@45672.4]
  assign x452_sum_1_io_a = RetimeWrapper_88_io_out; // @[Math.scala 151:17:@45673.4]
  assign x452_sum_1_io_b = RetimeWrapper_69_io_out; // @[Math.scala 152:17:@45674.4]
  assign x452_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@45675.4]
  assign RetimeWrapper_92_clock = clock; // @[:@45681.4]
  assign RetimeWrapper_92_reset = reset; // @[:@45682.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45684.4]
  assign RetimeWrapper_92_io_in = ~ x450; // @[package.scala 94:16:@45683.4]
  assign RetimeWrapper_93_clock = clock; // @[:@45693.4]
  assign RetimeWrapper_93_reset = reset; // @[:@45694.4]
  assign RetimeWrapper_93_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45696.4]
  assign RetimeWrapper_93_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45695.4]
  assign x457_sum_1_clock = clock; // @[:@45720.4]
  assign x457_sum_1_reset = reset; // @[:@45721.4]
  assign x457_sum_1_io_a = RetimeWrapper_88_io_out; // @[Math.scala 151:17:@45722.4]
  assign x457_sum_1_io_b = RetimeWrapper_72_io_out; // @[Math.scala 152:17:@45723.4]
  assign x457_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@45724.4]
  assign RetimeWrapper_94_clock = clock; // @[:@45730.4]
  assign RetimeWrapper_94_reset = reset; // @[:@45731.4]
  assign RetimeWrapper_94_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45733.4]
  assign RetimeWrapper_94_io_in = ~ x455; // @[package.scala 94:16:@45732.4]
  assign RetimeWrapper_95_clock = clock; // @[:@45742.4]
  assign RetimeWrapper_95_reset = reset; // @[:@45743.4]
  assign RetimeWrapper_95_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45745.4]
  assign RetimeWrapper_95_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45744.4]
  assign RetimeWrapper_96_clock = clock; // @[:@45769.4]
  assign RetimeWrapper_96_reset = reset; // @[:@45770.4]
  assign RetimeWrapper_96_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45772.4]
  assign RetimeWrapper_96_io_in = x631_sum_1_io_result; // @[package.scala 94:16:@45771.4]
  assign x462_sum_1_clock = clock; // @[:@45780.4]
  assign x462_sum_1_reset = reset; // @[:@45781.4]
  assign x462_sum_1_io_a = RetimeWrapper_96_io_out; // @[Math.scala 151:17:@45782.4]
  assign x462_sum_1_io_b = RetimeWrapper_76_io_out; // @[Math.scala 152:17:@45783.4]
  assign x462_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@45784.4]
  assign RetimeWrapper_97_clock = clock; // @[:@45790.4]
  assign RetimeWrapper_97_reset = reset; // @[:@45791.4]
  assign RetimeWrapper_97_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45793.4]
  assign RetimeWrapper_97_io_in = ~ x460; // @[package.scala 94:16:@45792.4]
  assign RetimeWrapper_98_clock = clock; // @[:@45799.4]
  assign RetimeWrapper_98_reset = reset; // @[:@45800.4]
  assign RetimeWrapper_98_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45802.4]
  assign RetimeWrapper_98_io_in = x462_sum_1_io_result; // @[package.scala 94:16:@45801.4]
  assign RetimeWrapper_99_clock = clock; // @[:@45811.4]
  assign RetimeWrapper_99_reset = reset; // @[:@45812.4]
  assign RetimeWrapper_99_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45814.4]
  assign RetimeWrapper_99_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45813.4]
  assign x467_sum_1_clock = clock; // @[:@45838.4]
  assign x467_sum_1_reset = reset; // @[:@45839.4]
  assign x467_sum_1_io_a = RetimeWrapper_88_io_out; // @[Math.scala 151:17:@45840.4]
  assign x467_sum_1_io_b = x390_div_1_io_result; // @[Math.scala 152:17:@45841.4]
  assign x467_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@45842.4]
  assign RetimeWrapper_100_clock = clock; // @[:@45848.4]
  assign RetimeWrapper_100_reset = reset; // @[:@45849.4]
  assign RetimeWrapper_100_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45851.4]
  assign RetimeWrapper_100_io_in = ~ x465; // @[package.scala 94:16:@45850.4]
  assign RetimeWrapper_101_clock = clock; // @[:@45860.4]
  assign RetimeWrapper_101_reset = reset; // @[:@45861.4]
  assign RetimeWrapper_101_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45863.4]
  assign RetimeWrapper_101_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45862.4]
  assign x472_sum_1_clock = clock; // @[:@45887.4]
  assign x472_sum_1_reset = reset; // @[:@45888.4]
  assign x472_sum_1_io_a = RetimeWrapper_88_io_out; // @[Math.scala 151:17:@45889.4]
  assign x472_sum_1_io_b = x399_div_1_io_result; // @[Math.scala 152:17:@45890.4]
  assign x472_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@45891.4]
  assign RetimeWrapper_102_clock = clock; // @[:@45897.4]
  assign RetimeWrapper_102_reset = reset; // @[:@45898.4]
  assign RetimeWrapper_102_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45900.4]
  assign RetimeWrapper_102_io_in = ~ x470; // @[package.scala 94:16:@45899.4]
  assign RetimeWrapper_103_clock = clock; // @[:@45909.4]
  assign RetimeWrapper_103_reset = reset; // @[:@45910.4]
  assign RetimeWrapper_103_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45912.4]
  assign RetimeWrapper_103_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45911.4]
  assign x475_1_clock = clock; // @[:@45932.4]
  assign x475_1_io_a = x334_lb_0_io_rPort_9_output_0; // @[Math.scala 263:17:@45934.4]
  assign x475_1_io_b = 32'h1; // @[Math.scala 264:17:@45935.4]
  assign x475_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@45936.4]
  assign x476_1_clock = clock; // @[:@45944.4]
  assign x476_1_io_a = x334_lb_0_io_rPort_15_output_0; // @[Math.scala 263:17:@45946.4]
  assign x476_1_io_b = 32'h2; // @[Math.scala 264:17:@45947.4]
  assign x476_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@45948.4]
  assign x477_1_clock = clock; // @[:@45956.4]
  assign x477_1_io_a = x334_lb_0_io_rPort_11_output_0; // @[Math.scala 263:17:@45958.4]
  assign x477_1_io_b = 32'h1; // @[Math.scala 264:17:@45959.4]
  assign x477_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@45960.4]
  assign x478_1_clock = clock; // @[:@45968.4]
  assign x478_1_io_a = x334_lb_0_io_rPort_5_output_0; // @[Math.scala 263:17:@45970.4]
  assign x478_1_io_b = 32'h2; // @[Math.scala 264:17:@45971.4]
  assign x478_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@45972.4]
  assign x479_1_clock = clock; // @[:@45980.4]
  assign x479_1_io_a = x334_lb_0_io_rPort_1_output_0; // @[Math.scala 263:17:@45982.4]
  assign x479_1_io_b = 32'h4; // @[Math.scala 264:17:@45983.4]
  assign x479_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@45984.4]
  assign x480_1_clock = clock; // @[:@45992.4]
  assign x480_1_io_a = x334_lb_0_io_rPort_14_output_0; // @[Math.scala 263:17:@45994.4]
  assign x480_1_io_b = 32'h2; // @[Math.scala 264:17:@45995.4]
  assign x480_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@45996.4]
  assign x481_1_clock = clock; // @[:@46004.4]
  assign x481_1_io_a = x334_lb_0_io_rPort_2_output_0; // @[Math.scala 263:17:@46006.4]
  assign x481_1_io_b = 32'h1; // @[Math.scala 264:17:@46007.4]
  assign x481_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46008.4]
  assign x482_1_clock = clock; // @[:@46016.4]
  assign x482_1_io_a = x334_lb_0_io_rPort_3_output_0; // @[Math.scala 263:17:@46018.4]
  assign x482_1_io_b = 32'h2; // @[Math.scala 264:17:@46019.4]
  assign x482_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46020.4]
  assign x483_1_clock = clock; // @[:@46028.4]
  assign x483_1_io_a = x334_lb_0_io_rPort_7_output_0; // @[Math.scala 263:17:@46030.4]
  assign x483_1_io_b = 32'h1; // @[Math.scala 264:17:@46031.4]
  assign x483_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46032.4]
  assign x484_x3_1_clock = clock; // @[:@46038.4]
  assign x484_x3_1_reset = reset; // @[:@46039.4]
  assign x484_x3_1_io_a = x475_1_io_result; // @[Math.scala 151:17:@46040.4]
  assign x484_x3_1_io_b = x476_1_io_result; // @[Math.scala 152:17:@46041.4]
  assign x484_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46042.4]
  assign x485_x4_1_clock = clock; // @[:@46048.4]
  assign x485_x4_1_reset = reset; // @[:@46049.4]
  assign x485_x4_1_io_a = x477_1_io_result; // @[Math.scala 151:17:@46050.4]
  assign x485_x4_1_io_b = x478_1_io_result; // @[Math.scala 152:17:@46051.4]
  assign x485_x4_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46052.4]
  assign x486_x3_1_clock = clock; // @[:@46058.4]
  assign x486_x3_1_reset = reset; // @[:@46059.4]
  assign x486_x3_1_io_a = x479_1_io_result; // @[Math.scala 151:17:@46060.4]
  assign x486_x3_1_io_b = x480_1_io_result; // @[Math.scala 152:17:@46061.4]
  assign x486_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46062.4]
  assign x487_x4_1_clock = clock; // @[:@46068.4]
  assign x487_x4_1_reset = reset; // @[:@46069.4]
  assign x487_x4_1_io_a = x481_1_io_result; // @[Math.scala 151:17:@46070.4]
  assign x487_x4_1_io_b = x482_1_io_result; // @[Math.scala 152:17:@46071.4]
  assign x487_x4_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46072.4]
  assign x488_x3_1_clock = clock; // @[:@46078.4]
  assign x488_x3_1_reset = reset; // @[:@46079.4]
  assign x488_x3_1_io_a = x484_x3_1_io_result; // @[Math.scala 151:17:@46080.4]
  assign x488_x3_1_io_b = x485_x4_1_io_result; // @[Math.scala 152:17:@46081.4]
  assign x488_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46082.4]
  assign x489_x4_1_clock = clock; // @[:@46088.4]
  assign x489_x4_1_reset = reset; // @[:@46089.4]
  assign x489_x4_1_io_a = x486_x3_1_io_result; // @[Math.scala 151:17:@46090.4]
  assign x489_x4_1_io_b = x487_x4_1_io_result; // @[Math.scala 152:17:@46091.4]
  assign x489_x4_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46092.4]
  assign x490_x3_1_clock = clock; // @[:@46098.4]
  assign x490_x3_1_reset = reset; // @[:@46099.4]
  assign x490_x3_1_io_a = x488_x3_1_io_result; // @[Math.scala 151:17:@46100.4]
  assign x490_x3_1_io_b = x489_x4_1_io_result; // @[Math.scala 152:17:@46101.4]
  assign x490_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46102.4]
  assign RetimeWrapper_104_clock = clock; // @[:@46108.4]
  assign RetimeWrapper_104_reset = reset; // @[:@46109.4]
  assign RetimeWrapper_104_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46111.4]
  assign RetimeWrapper_104_io_in = x483_1_io_result; // @[package.scala 94:16:@46110.4]
  assign x491_sum_1_clock = clock; // @[:@46117.4]
  assign x491_sum_1_reset = reset; // @[:@46118.4]
  assign x491_sum_1_io_a = x490_x3_1_io_result; // @[Math.scala 151:17:@46119.4]
  assign x491_sum_1_io_b = RetimeWrapper_104_io_out; // @[Math.scala 152:17:@46120.4]
  assign x491_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46121.4]
  assign x492_1_io_b = x491_sum_1_io_result; // @[Math.scala 721:17:@46129.4]
  assign x493_mul_1_clock = clock; // @[:@46138.4]
  assign x493_mul_1_io_a = x492_1_io_result; // @[Math.scala 263:17:@46140.4]
  assign x493_mul_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46142.4]
  assign x494_1_io_b = x493_mul_1_io_result; // @[Math.scala 721:17:@46150.4]
  assign x495_1_clock = clock; // @[:@46159.4]
  assign x495_1_io_a = x334_lb_0_io_rPort_15_output_0; // @[Math.scala 263:17:@46161.4]
  assign x495_1_io_b = 32'h1; // @[Math.scala 264:17:@46162.4]
  assign x495_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46163.4]
  assign x496_1_clock = clock; // @[:@46171.4]
  assign x496_1_io_a = x334_lb_0_io_rPort_11_output_0; // @[Math.scala 263:17:@46173.4]
  assign x496_1_io_b = 32'h2; // @[Math.scala 264:17:@46174.4]
  assign x496_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46175.4]
  assign x497_1_clock = clock; // @[:@46183.4]
  assign x497_1_io_a = x334_lb_0_io_rPort_12_output_0; // @[Math.scala 263:17:@46185.4]
  assign x497_1_io_b = 32'h1; // @[Math.scala 264:17:@46186.4]
  assign x497_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46187.4]
  assign x498_1_clock = clock; // @[:@46195.4]
  assign x498_1_io_a = x334_lb_0_io_rPort_1_output_0; // @[Math.scala 263:17:@46197.4]
  assign x498_1_io_b = 32'h2; // @[Math.scala 264:17:@46198.4]
  assign x498_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46199.4]
  assign x499_1_clock = clock; // @[:@46207.4]
  assign x499_1_io_a = x334_lb_0_io_rPort_14_output_0; // @[Math.scala 263:17:@46209.4]
  assign x499_1_io_b = 32'h4; // @[Math.scala 264:17:@46210.4]
  assign x499_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46211.4]
  assign x500_1_clock = clock; // @[:@46219.4]
  assign x500_1_io_a = x334_lb_0_io_rPort_17_output_0; // @[Math.scala 263:17:@46221.4]
  assign x500_1_io_b = 32'h2; // @[Math.scala 264:17:@46222.4]
  assign x500_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46223.4]
  assign x501_1_clock = clock; // @[:@46233.4]
  assign x501_1_io_a = x334_lb_0_io_rPort_3_output_0; // @[Math.scala 263:17:@46235.4]
  assign x501_1_io_b = 32'h1; // @[Math.scala 264:17:@46236.4]
  assign x501_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46237.4]
  assign x502_1_clock = clock; // @[:@46245.4]
  assign x502_1_io_a = x334_lb_0_io_rPort_7_output_0; // @[Math.scala 263:17:@46247.4]
  assign x502_1_io_b = 32'h2; // @[Math.scala 264:17:@46248.4]
  assign x502_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46249.4]
  assign x503_1_clock = clock; // @[:@46257.4]
  assign x503_1_io_a = x334_lb_0_io_rPort_8_output_0; // @[Math.scala 263:17:@46259.4]
  assign x503_1_io_b = 32'h1; // @[Math.scala 264:17:@46260.4]
  assign x503_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46261.4]
  assign x504_x3_1_clock = clock; // @[:@46267.4]
  assign x504_x3_1_reset = reset; // @[:@46268.4]
  assign x504_x3_1_io_a = x495_1_io_result; // @[Math.scala 151:17:@46269.4]
  assign x504_x3_1_io_b = x496_1_io_result; // @[Math.scala 152:17:@46270.4]
  assign x504_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46271.4]
  assign x505_x4_1_clock = clock; // @[:@46277.4]
  assign x505_x4_1_reset = reset; // @[:@46278.4]
  assign x505_x4_1_io_a = x497_1_io_result; // @[Math.scala 151:17:@46279.4]
  assign x505_x4_1_io_b = x498_1_io_result; // @[Math.scala 152:17:@46280.4]
  assign x505_x4_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46281.4]
  assign x506_x3_1_clock = clock; // @[:@46287.4]
  assign x506_x3_1_reset = reset; // @[:@46288.4]
  assign x506_x3_1_io_a = x499_1_io_result; // @[Math.scala 151:17:@46289.4]
  assign x506_x3_1_io_b = x500_1_io_result; // @[Math.scala 152:17:@46290.4]
  assign x506_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46291.4]
  assign x507_x4_1_clock = clock; // @[:@46297.4]
  assign x507_x4_1_reset = reset; // @[:@46298.4]
  assign x507_x4_1_io_a = x501_1_io_result; // @[Math.scala 151:17:@46299.4]
  assign x507_x4_1_io_b = x502_1_io_result; // @[Math.scala 152:17:@46300.4]
  assign x507_x4_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46301.4]
  assign x508_x3_1_clock = clock; // @[:@46307.4]
  assign x508_x3_1_reset = reset; // @[:@46308.4]
  assign x508_x3_1_io_a = x504_x3_1_io_result; // @[Math.scala 151:17:@46309.4]
  assign x508_x3_1_io_b = x505_x4_1_io_result; // @[Math.scala 152:17:@46310.4]
  assign x508_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46311.4]
  assign x509_x4_1_clock = clock; // @[:@46317.4]
  assign x509_x4_1_reset = reset; // @[:@46318.4]
  assign x509_x4_1_io_a = x506_x3_1_io_result; // @[Math.scala 151:17:@46319.4]
  assign x509_x4_1_io_b = x507_x4_1_io_result; // @[Math.scala 152:17:@46320.4]
  assign x509_x4_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46321.4]
  assign x510_x3_1_clock = clock; // @[:@46327.4]
  assign x510_x3_1_reset = reset; // @[:@46328.4]
  assign x510_x3_1_io_a = x508_x3_1_io_result; // @[Math.scala 151:17:@46329.4]
  assign x510_x3_1_io_b = x509_x4_1_io_result; // @[Math.scala 152:17:@46330.4]
  assign x510_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46331.4]
  assign RetimeWrapper_105_clock = clock; // @[:@46337.4]
  assign RetimeWrapper_105_reset = reset; // @[:@46338.4]
  assign RetimeWrapper_105_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46340.4]
  assign RetimeWrapper_105_io_in = x503_1_io_result; // @[package.scala 94:16:@46339.4]
  assign x511_sum_1_clock = clock; // @[:@46346.4]
  assign x511_sum_1_reset = reset; // @[:@46347.4]
  assign x511_sum_1_io_a = x510_x3_1_io_result; // @[Math.scala 151:17:@46348.4]
  assign x511_sum_1_io_b = RetimeWrapper_105_io_out; // @[Math.scala 152:17:@46349.4]
  assign x511_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46350.4]
  assign x512_1_io_b = x511_sum_1_io_result; // @[Math.scala 721:17:@46358.4]
  assign x513_mul_1_clock = clock; // @[:@46367.4]
  assign x513_mul_1_io_a = x512_1_io_result; // @[Math.scala 263:17:@46369.4]
  assign x513_mul_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46371.4]
  assign x514_1_io_b = x513_mul_1_io_result; // @[Math.scala 721:17:@46379.4]
  assign x515_1_clock = clock; // @[:@46388.4]
  assign x515_1_io_a = x334_lb_0_io_rPort_12_output_0; // @[Math.scala 263:17:@46390.4]
  assign x515_1_io_b = 32'h2; // @[Math.scala 264:17:@46391.4]
  assign x515_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46392.4]
  assign x516_1_clock = clock; // @[:@46400.4]
  assign x516_1_io_a = x334_lb_0_io_rPort_4_output_0; // @[Math.scala 263:17:@46402.4]
  assign x516_1_io_b = 32'h1; // @[Math.scala 264:17:@46403.4]
  assign x516_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46404.4]
  assign x517_1_clock = clock; // @[:@46412.4]
  assign x517_1_io_a = x334_lb_0_io_rPort_17_output_0; // @[Math.scala 263:17:@46414.4]
  assign x517_1_io_b = 32'h4; // @[Math.scala 264:17:@46415.4]
  assign x517_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46416.4]
  assign x518_1_clock = clock; // @[:@46424.4]
  assign x518_1_io_a = x334_lb_0_io_rPort_13_output_0; // @[Math.scala 263:17:@46426.4]
  assign x518_1_io_b = 32'h2; // @[Math.scala 264:17:@46427.4]
  assign x518_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46428.4]
  assign x519_1_clock = clock; // @[:@46436.4]
  assign x519_1_io_a = x334_lb_0_io_rPort_8_output_0; // @[Math.scala 263:17:@46438.4]
  assign x519_1_io_b = 32'h2; // @[Math.scala 264:17:@46439.4]
  assign x519_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46440.4]
  assign x520_1_clock = clock; // @[:@46448.4]
  assign x520_1_io_a = x334_lb_0_io_rPort_0_output_0; // @[Math.scala 263:17:@46450.4]
  assign x520_1_io_b = 32'h1; // @[Math.scala 264:17:@46451.4]
  assign x520_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46452.4]
  assign x521_x3_1_clock = clock; // @[:@46458.4]
  assign x521_x3_1_reset = reset; // @[:@46459.4]
  assign x521_x3_1_io_a = x477_1_io_result; // @[Math.scala 151:17:@46460.4]
  assign x521_x3_1_io_b = x515_1_io_result; // @[Math.scala 152:17:@46461.4]
  assign x521_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46462.4]
  assign x522_x4_1_clock = clock; // @[:@46468.4]
  assign x522_x4_1_reset = reset; // @[:@46469.4]
  assign x522_x4_1_io_a = x516_1_io_result; // @[Math.scala 151:17:@46470.4]
  assign x522_x4_1_io_b = x480_1_io_result; // @[Math.scala 152:17:@46471.4]
  assign x522_x4_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46472.4]
  assign x523_x3_1_clock = clock; // @[:@46478.4]
  assign x523_x3_1_reset = reset; // @[:@46479.4]
  assign x523_x3_1_io_a = x517_1_io_result; // @[Math.scala 151:17:@46480.4]
  assign x523_x3_1_io_b = x518_1_io_result; // @[Math.scala 152:17:@46481.4]
  assign x523_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46482.4]
  assign x524_x4_1_clock = clock; // @[:@46488.4]
  assign x524_x4_1_reset = reset; // @[:@46489.4]
  assign x524_x4_1_io_a = x483_1_io_result; // @[Math.scala 151:17:@46490.4]
  assign x524_x4_1_io_b = x519_1_io_result; // @[Math.scala 152:17:@46491.4]
  assign x524_x4_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46492.4]
  assign x525_x3_1_clock = clock; // @[:@46498.4]
  assign x525_x3_1_reset = reset; // @[:@46499.4]
  assign x525_x3_1_io_a = x521_x3_1_io_result; // @[Math.scala 151:17:@46500.4]
  assign x525_x3_1_io_b = x522_x4_1_io_result; // @[Math.scala 152:17:@46501.4]
  assign x525_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46502.4]
  assign x526_x4_1_clock = clock; // @[:@46508.4]
  assign x526_x4_1_reset = reset; // @[:@46509.4]
  assign x526_x4_1_io_a = x523_x3_1_io_result; // @[Math.scala 151:17:@46510.4]
  assign x526_x4_1_io_b = x524_x4_1_io_result; // @[Math.scala 152:17:@46511.4]
  assign x526_x4_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46512.4]
  assign x527_x3_1_clock = clock; // @[:@46518.4]
  assign x527_x3_1_reset = reset; // @[:@46519.4]
  assign x527_x3_1_io_a = x525_x3_1_io_result; // @[Math.scala 151:17:@46520.4]
  assign x527_x3_1_io_b = x526_x4_1_io_result; // @[Math.scala 152:17:@46521.4]
  assign x527_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46522.4]
  assign RetimeWrapper_106_clock = clock; // @[:@46528.4]
  assign RetimeWrapper_106_reset = reset; // @[:@46529.4]
  assign RetimeWrapper_106_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46531.4]
  assign RetimeWrapper_106_io_in = x520_1_io_result; // @[package.scala 94:16:@46530.4]
  assign x528_sum_1_clock = clock; // @[:@46537.4]
  assign x528_sum_1_reset = reset; // @[:@46538.4]
  assign x528_sum_1_io_a = x527_x3_1_io_result; // @[Math.scala 151:17:@46539.4]
  assign x528_sum_1_io_b = RetimeWrapper_106_io_out; // @[Math.scala 152:17:@46540.4]
  assign x528_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46541.4]
  assign x529_1_io_b = x528_sum_1_io_result; // @[Math.scala 721:17:@46549.4]
  assign x530_mul_1_clock = clock; // @[:@46558.4]
  assign x530_mul_1_io_a = x529_1_io_result; // @[Math.scala 263:17:@46560.4]
  assign x530_mul_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46562.4]
  assign x531_1_io_b = x530_mul_1_io_result; // @[Math.scala 721:17:@46570.4]
  assign x532_1_clock = clock; // @[:@46579.4]
  assign x532_1_io_a = x334_lb_0_io_rPort_4_output_0; // @[Math.scala 263:17:@46581.4]
  assign x532_1_io_b = 32'h2; // @[Math.scala 264:17:@46582.4]
  assign x532_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46583.4]
  assign x533_1_clock = clock; // @[:@46591.4]
  assign x533_1_io_a = x334_lb_0_io_rPort_10_output_0; // @[Math.scala 263:17:@46593.4]
  assign x533_1_io_b = 32'h1; // @[Math.scala 264:17:@46594.4]
  assign x533_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46595.4]
  assign x534_1_clock = clock; // @[:@46603.4]
  assign x534_1_io_a = x334_lb_0_io_rPort_13_output_0; // @[Math.scala 263:17:@46605.4]
  assign x534_1_io_b = 32'h4; // @[Math.scala 264:17:@46606.4]
  assign x534_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46607.4]
  assign x535_1_clock = clock; // @[:@46615.4]
  assign x535_1_io_a = x334_lb_0_io_rPort_16_output_0; // @[Math.scala 263:17:@46617.4]
  assign x535_1_io_b = 32'h2; // @[Math.scala 264:17:@46618.4]
  assign x535_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46619.4]
  assign x536_1_clock = clock; // @[:@46627.4]
  assign x536_1_io_a = x334_lb_0_io_rPort_0_output_0; // @[Math.scala 263:17:@46629.4]
  assign x536_1_io_b = 32'h2; // @[Math.scala 264:17:@46630.4]
  assign x536_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46631.4]
  assign x537_1_clock = clock; // @[:@46639.4]
  assign x537_1_io_a = x334_lb_0_io_rPort_6_output_0; // @[Math.scala 263:17:@46641.4]
  assign x537_1_io_b = 32'h1; // @[Math.scala 264:17:@46642.4]
  assign x537_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46643.4]
  assign x538_x3_1_clock = clock; // @[:@46649.4]
  assign x538_x3_1_reset = reset; // @[:@46650.4]
  assign x538_x3_1_io_a = x497_1_io_result; // @[Math.scala 151:17:@46651.4]
  assign x538_x3_1_io_b = x532_1_io_result; // @[Math.scala 152:17:@46652.4]
  assign x538_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46653.4]
  assign x539_x4_1_clock = clock; // @[:@46659.4]
  assign x539_x4_1_reset = reset; // @[:@46660.4]
  assign x539_x4_1_io_a = x533_1_io_result; // @[Math.scala 151:17:@46661.4]
  assign x539_x4_1_io_b = x500_1_io_result; // @[Math.scala 152:17:@46662.4]
  assign x539_x4_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46663.4]
  assign x540_x3_1_clock = clock; // @[:@46669.4]
  assign x540_x3_1_reset = reset; // @[:@46670.4]
  assign x540_x3_1_io_a = x534_1_io_result; // @[Math.scala 151:17:@46671.4]
  assign x540_x3_1_io_b = x535_1_io_result; // @[Math.scala 152:17:@46672.4]
  assign x540_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46673.4]
  assign x541_x4_1_clock = clock; // @[:@46679.4]
  assign x541_x4_1_reset = reset; // @[:@46680.4]
  assign x541_x4_1_io_a = x503_1_io_result; // @[Math.scala 151:17:@46681.4]
  assign x541_x4_1_io_b = x536_1_io_result; // @[Math.scala 152:17:@46682.4]
  assign x541_x4_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46683.4]
  assign x542_x3_1_clock = clock; // @[:@46689.4]
  assign x542_x3_1_reset = reset; // @[:@46690.4]
  assign x542_x3_1_io_a = x538_x3_1_io_result; // @[Math.scala 151:17:@46691.4]
  assign x542_x3_1_io_b = x539_x4_1_io_result; // @[Math.scala 152:17:@46692.4]
  assign x542_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46693.4]
  assign x543_x4_1_clock = clock; // @[:@46699.4]
  assign x543_x4_1_reset = reset; // @[:@46700.4]
  assign x543_x4_1_io_a = x540_x3_1_io_result; // @[Math.scala 151:17:@46701.4]
  assign x543_x4_1_io_b = x541_x4_1_io_result; // @[Math.scala 152:17:@46702.4]
  assign x543_x4_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46703.4]
  assign x544_x3_1_clock = clock; // @[:@46709.4]
  assign x544_x3_1_reset = reset; // @[:@46710.4]
  assign x544_x3_1_io_a = x542_x3_1_io_result; // @[Math.scala 151:17:@46711.4]
  assign x544_x3_1_io_b = x543_x4_1_io_result; // @[Math.scala 152:17:@46712.4]
  assign x544_x3_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46713.4]
  assign RetimeWrapper_107_clock = clock; // @[:@46719.4]
  assign RetimeWrapper_107_reset = reset; // @[:@46720.4]
  assign RetimeWrapper_107_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46722.4]
  assign RetimeWrapper_107_io_in = x537_1_io_result; // @[package.scala 94:16:@46721.4]
  assign x545_sum_1_clock = clock; // @[:@46728.4]
  assign x545_sum_1_reset = reset; // @[:@46729.4]
  assign x545_sum_1_io_a = x544_x3_1_io_result; // @[Math.scala 151:17:@46730.4]
  assign x545_sum_1_io_b = RetimeWrapper_107_io_out; // @[Math.scala 152:17:@46731.4]
  assign x545_sum_1_io_flow = io_in_x290_TREADY; // @[Math.scala 153:20:@46732.4]
  assign x546_1_io_b = x545_sum_1_io_result; // @[Math.scala 721:17:@46740.4]
  assign x547_mul_1_clock = clock; // @[:@46751.4]
  assign x547_mul_1_io_a = x546_1_io_result; // @[Math.scala 263:17:@46753.4]
  assign x547_mul_1_io_flow = io_in_x290_TREADY; // @[Math.scala 265:20:@46755.4]
  assign x548_1_io_b = x547_mul_1_io_result; // @[Math.scala 721:17:@46763.4]
  assign RetimeWrapper_108_clock = clock; // @[:@46780.4]
  assign RetimeWrapper_108_reset = reset; // @[:@46781.4]
  assign RetimeWrapper_108_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46783.4]
  assign RetimeWrapper_108_io_in = {_T_1778,_T_1777}; // @[package.scala 94:16:@46782.4]
  assign RetimeWrapper_109_clock = clock; // @[:@46789.4]
  assign RetimeWrapper_109_reset = reset; // @[:@46790.4]
  assign RetimeWrapper_109_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46792.4]
  assign RetimeWrapper_109_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@46791.4]
  assign RetimeWrapper_110_clock = clock; // @[:@46798.4]
  assign RetimeWrapper_110_reset = reset; // @[:@46799.4]
  assign RetimeWrapper_110_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46801.4]
  assign RetimeWrapper_110_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@46800.4]
  assign RetimeWrapper_111_clock = clock; // @[:@46807.4]
  assign RetimeWrapper_111_reset = reset; // @[:@46808.4]
  assign RetimeWrapper_111_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46810.4]
  assign RetimeWrapper_111_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46809.4]
endmodule
module x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1( // @[:@46828.2]
  input          clock, // @[:@46829.4]
  input          reset, // @[:@46830.4]
  input          io_in_x289_TVALID, // @[:@46831.4]
  output         io_in_x289_TREADY, // @[:@46831.4]
  input  [255:0] io_in_x289_TDATA, // @[:@46831.4]
  input  [7:0]   io_in_x289_TID, // @[:@46831.4]
  input  [7:0]   io_in_x289_TDEST, // @[:@46831.4]
  output         io_in_x290_TVALID, // @[:@46831.4]
  input          io_in_x290_TREADY, // @[:@46831.4]
  output [255:0] io_in_x290_TDATA, // @[:@46831.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@46831.4]
  input          io_sigsIn_smChildAcks_0, // @[:@46831.4]
  output         io_sigsOut_smDoneIn_0, // @[:@46831.4]
  input          io_rr // @[:@46831.4]
);
  wire  x327_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@46865.4]
  wire  x327_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@46865.4]
  wire  x327_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@46865.4]
  wire  x327_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@46865.4]
  wire [12:0] x327_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@46865.4]
  wire [12:0] x327_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@46865.4]
  wire  x327_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@46865.4]
  wire  x327_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@46865.4]
  wire  x327_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@46865.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 32:18:@46925.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 32:18:@46925.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 32:18:@46925.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 32:18:@46925.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 32:18:@46925.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 32:18:@46925.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 32:18:@46925.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 32:18:@46925.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 32:18:@46925.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 32:18:@46925.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 32:18:@46925.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 32:18:@46925.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@46953.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@46953.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@46953.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@46953.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@46953.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@46995.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@46995.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@46995.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@46995.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@46995.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@47003.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@47003.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@47003.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@47003.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@47003.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x289_TREADY; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire [255:0] x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x289_TDATA; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire [7:0] x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x289_TID; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire [7:0] x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x289_TDEST; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x290_TVALID; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x290_TREADY; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire [255:0] x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x290_TDATA; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire [31:0] x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire [31:0] x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
  wire  _T_240; // @[package.scala 96:25:@46958.4 package.scala 96:25:@46959.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x554_outr_UnitPipe.scala 69:66:@46964.4]
  wire  _T_253; // @[package.scala 96:25:@47000.4 package.scala 96:25:@47001.4]
  wire  _T_259; // @[package.scala 96:25:@47008.4 package.scala 96:25:@47009.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@47011.4]
  wire  x553_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@47012.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@47020.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@47021.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@47033.4]
  x297_ctrchain x327_ctrchain ( // @[SpatialBlocks.scala 37:22:@46865.4]
    .clock(x327_ctrchain_clock),
    .reset(x327_ctrchain_reset),
    .io_input_reset(x327_ctrchain_io_input_reset),
    .io_input_enable(x327_ctrchain_io_input_enable),
    .io_output_counts_1(x327_ctrchain_io_output_counts_1),
    .io_output_counts_0(x327_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x327_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x327_ctrchain_io_output_oobs_1),
    .io_output_done(x327_ctrchain_io_output_done)
  );
  x553_inr_Foreach_SAMPLER_BOX_sm x553_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 32:18:@46925.4]
    .clock(x553_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x553_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x553_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x553_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x553_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x553_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x553_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x553_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x553_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x553_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x553_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x553_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@46953.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@46995.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@47003.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1 x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 796:24:@47037.4]
    .clock(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x289_TREADY(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x289_TREADY),
    .io_in_x289_TDATA(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x289_TDATA),
    .io_in_x289_TID(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x289_TID),
    .io_in_x289_TDEST(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x289_TDEST),
    .io_in_x290_TVALID(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x290_TVALID),
    .io_in_x290_TREADY(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x290_TREADY),
    .io_in_x290_TDATA(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x290_TDATA),
    .io_sigsIn_backpressure(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@46958.4 package.scala 96:25:@46959.4]
  assign x553_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x289_TVALID | x553_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x554_outr_UnitPipe.scala 69:66:@46964.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@47000.4 package.scala 96:25:@47001.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@47008.4 package.scala 96:25:@47009.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@47011.4]
  assign x553_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@47012.4]
  assign _T_264 = x553_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@47020.4]
  assign _T_265 = ~ x553_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@47021.4]
  assign _T_272 = x553_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@47033.4]
  assign io_in_x289_TREADY = x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x289_TREADY; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 48:23:@47095.4]
  assign io_in_x290_TVALID = x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x290_TVALID; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 49:23:@47105.4]
  assign io_in_x290_TDATA = x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x290_TDATA; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 49:23:@47103.4]
  assign io_sigsOut_smDoneIn_0 = x553_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@47018.4]
  assign x327_ctrchain_clock = clock; // @[:@46866.4]
  assign x327_ctrchain_reset = reset; // @[:@46867.4]
  assign x327_ctrchain_io_input_reset = x553_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@47036.4]
  assign x327_ctrchain_io_input_enable = _T_272 & x553_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@46988.4 SpatialBlocks.scala 159:42:@47035.4]
  assign x553_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@46926.4]
  assign x553_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@46927.4]
  assign x553_inr_Foreach_SAMPLER_BOX_sm_io_enable = x553_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x553_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@47015.4]
  assign x553_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x554_outr_UnitPipe.scala 67:50:@46961.4]
  assign x553_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@47017.4]
  assign x553_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x290_TREADY | x553_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@46989.4]
  assign x553_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x554_outr_UnitPipe.scala 71:48:@46967.4]
  assign RetimeWrapper_clock = clock; // @[:@46954.4]
  assign RetimeWrapper_reset = reset; // @[:@46955.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@46957.4]
  assign RetimeWrapper_io_in = x327_ctrchain_io_output_done; // @[package.scala 94:16:@46956.4]
  assign RetimeWrapper_1_clock = clock; // @[:@46996.4]
  assign RetimeWrapper_1_reset = reset; // @[:@46997.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@46999.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@46998.4]
  assign RetimeWrapper_2_clock = clock; // @[:@47004.4]
  assign RetimeWrapper_2_reset = reset; // @[:@47005.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@47007.4]
  assign RetimeWrapper_2_io_in = x553_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@47006.4]
  assign x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@47038.4]
  assign x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@47039.4]
  assign x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x289_TDATA = io_in_x289_TDATA; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 48:23:@47094.4]
  assign x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x289_TID = io_in_x289_TID; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 48:23:@47090.4]
  assign x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x289_TDEST = io_in_x289_TDEST; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 48:23:@47089.4]
  assign x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x290_TREADY = io_in_x290_TREADY; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 49:23:@47104.4]
  assign x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x290_TREADY | x553_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 801:22:@47122.4]
  assign x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 801:22:@47120.4]
  assign x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x553_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 801:22:@47118.4]
  assign x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x327_ctrchain_io_output_counts_1[12]}},x327_ctrchain_io_output_counts_1}; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 801:22:@47113.4]
  assign x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x327_ctrchain_io_output_counts_0[12]}},x327_ctrchain_io_output_counts_0}; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 801:22:@47112.4]
  assign x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x327_ctrchain_io_output_oobs_0; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 801:22:@47110.4]
  assign x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x327_ctrchain_io_output_oobs_1; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 801:22:@47111.4]
  assign x553_inr_Foreach_SAMPLER_BOX_kernelx553_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x553_inr_Foreach_SAMPLER_BOX.scala 800:18:@47106.4]
endmodule
module x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1( // @[:@47136.2]
  input          clock, // @[:@47137.4]
  input          reset, // @[:@47138.4]
  input          io_in_x289_TVALID, // @[:@47139.4]
  output         io_in_x289_TREADY, // @[:@47139.4]
  input  [255:0] io_in_x289_TDATA, // @[:@47139.4]
  input  [7:0]   io_in_x289_TID, // @[:@47139.4]
  input  [7:0]   io_in_x289_TDEST, // @[:@47139.4]
  output         io_in_x290_TVALID, // @[:@47139.4]
  input          io_in_x290_TREADY, // @[:@47139.4]
  output [255:0] io_in_x290_TDATA, // @[:@47139.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@47139.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@47139.4]
  input          io_sigsIn_smChildAcks_0, // @[:@47139.4]
  input          io_sigsIn_smChildAcks_1, // @[:@47139.4]
  output         io_sigsOut_smDoneIn_0, // @[:@47139.4]
  output         io_sigsOut_smDoneIn_1, // @[:@47139.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@47139.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@47139.4]
  input          io_rr // @[:@47139.4]
);
  wire  x292_fifoinraw_0_clock; // @[m_x292_fifoinraw_0.scala 27:17:@47153.4]
  wire  x292_fifoinraw_0_reset; // @[m_x292_fifoinraw_0.scala 27:17:@47153.4]
  wire  x293_fifoinpacked_0_clock; // @[m_x293_fifoinpacked_0.scala 27:17:@47177.4]
  wire  x293_fifoinpacked_0_reset; // @[m_x293_fifoinpacked_0.scala 27:17:@47177.4]
  wire  x293_fifoinpacked_0_io_wPort_0_en_0; // @[m_x293_fifoinpacked_0.scala 27:17:@47177.4]
  wire  x293_fifoinpacked_0_io_full; // @[m_x293_fifoinpacked_0.scala 27:17:@47177.4]
  wire  x293_fifoinpacked_0_io_active_0_in; // @[m_x293_fifoinpacked_0.scala 27:17:@47177.4]
  wire  x293_fifoinpacked_0_io_active_0_out; // @[m_x293_fifoinpacked_0.scala 27:17:@47177.4]
  wire  x294_fifooutraw_0_clock; // @[m_x294_fifooutraw_0.scala 27:17:@47201.4]
  wire  x294_fifooutraw_0_reset; // @[m_x294_fifooutraw_0.scala 27:17:@47201.4]
  wire  x297_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@47225.4]
  wire  x297_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@47225.4]
  wire  x297_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@47225.4]
  wire  x297_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@47225.4]
  wire [12:0] x297_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@47225.4]
  wire [12:0] x297_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@47225.4]
  wire  x297_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@47225.4]
  wire  x297_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@47225.4]
  wire  x297_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@47225.4]
  wire  x323_inr_Foreach_sm_clock; // @[sm_x323_inr_Foreach.scala 32:18:@47285.4]
  wire  x323_inr_Foreach_sm_reset; // @[sm_x323_inr_Foreach.scala 32:18:@47285.4]
  wire  x323_inr_Foreach_sm_io_enable; // @[sm_x323_inr_Foreach.scala 32:18:@47285.4]
  wire  x323_inr_Foreach_sm_io_done; // @[sm_x323_inr_Foreach.scala 32:18:@47285.4]
  wire  x323_inr_Foreach_sm_io_doneLatch; // @[sm_x323_inr_Foreach.scala 32:18:@47285.4]
  wire  x323_inr_Foreach_sm_io_ctrDone; // @[sm_x323_inr_Foreach.scala 32:18:@47285.4]
  wire  x323_inr_Foreach_sm_io_datapathEn; // @[sm_x323_inr_Foreach.scala 32:18:@47285.4]
  wire  x323_inr_Foreach_sm_io_ctrInc; // @[sm_x323_inr_Foreach.scala 32:18:@47285.4]
  wire  x323_inr_Foreach_sm_io_ctrRst; // @[sm_x323_inr_Foreach.scala 32:18:@47285.4]
  wire  x323_inr_Foreach_sm_io_parentAck; // @[sm_x323_inr_Foreach.scala 32:18:@47285.4]
  wire  x323_inr_Foreach_sm_io_backpressure; // @[sm_x323_inr_Foreach.scala 32:18:@47285.4]
  wire  x323_inr_Foreach_sm_io_break; // @[sm_x323_inr_Foreach.scala 32:18:@47285.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@47313.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@47313.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@47313.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@47313.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@47313.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@47359.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@47359.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@47359.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@47359.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@47359.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@47367.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@47367.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@47367.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@47367.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@47367.4]
  wire  x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_clock; // @[sm_x323_inr_Foreach.scala 126:24:@47402.4]
  wire  x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_reset; // @[sm_x323_inr_Foreach.scala 126:24:@47402.4]
  wire  x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_in_x293_fifoinpacked_0_wPort_0_en_0; // @[sm_x323_inr_Foreach.scala 126:24:@47402.4]
  wire  x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_in_x293_fifoinpacked_0_full; // @[sm_x323_inr_Foreach.scala 126:24:@47402.4]
  wire  x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_in_x293_fifoinpacked_0_active_0_in; // @[sm_x323_inr_Foreach.scala 126:24:@47402.4]
  wire  x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_in_x293_fifoinpacked_0_active_0_out; // @[sm_x323_inr_Foreach.scala 126:24:@47402.4]
  wire  x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x323_inr_Foreach.scala 126:24:@47402.4]
  wire  x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x323_inr_Foreach.scala 126:24:@47402.4]
  wire  x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x323_inr_Foreach.scala 126:24:@47402.4]
  wire [31:0] x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x323_inr_Foreach.scala 126:24:@47402.4]
  wire [31:0] x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x323_inr_Foreach.scala 126:24:@47402.4]
  wire  x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x323_inr_Foreach.scala 126:24:@47402.4]
  wire  x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x323_inr_Foreach.scala 126:24:@47402.4]
  wire  x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_rr; // @[sm_x323_inr_Foreach.scala 126:24:@47402.4]
  wire  x554_outr_UnitPipe_sm_clock; // @[sm_x554_outr_UnitPipe.scala 32:18:@47534.4]
  wire  x554_outr_UnitPipe_sm_reset; // @[sm_x554_outr_UnitPipe.scala 32:18:@47534.4]
  wire  x554_outr_UnitPipe_sm_io_enable; // @[sm_x554_outr_UnitPipe.scala 32:18:@47534.4]
  wire  x554_outr_UnitPipe_sm_io_done; // @[sm_x554_outr_UnitPipe.scala 32:18:@47534.4]
  wire  x554_outr_UnitPipe_sm_io_rst; // @[sm_x554_outr_UnitPipe.scala 32:18:@47534.4]
  wire  x554_outr_UnitPipe_sm_io_ctrDone; // @[sm_x554_outr_UnitPipe.scala 32:18:@47534.4]
  wire  x554_outr_UnitPipe_sm_io_ctrInc; // @[sm_x554_outr_UnitPipe.scala 32:18:@47534.4]
  wire  x554_outr_UnitPipe_sm_io_parentAck; // @[sm_x554_outr_UnitPipe.scala 32:18:@47534.4]
  wire  x554_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x554_outr_UnitPipe.scala 32:18:@47534.4]
  wire  x554_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x554_outr_UnitPipe.scala 32:18:@47534.4]
  wire  x554_outr_UnitPipe_sm_io_childAck_0; // @[sm_x554_outr_UnitPipe.scala 32:18:@47534.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@47591.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@47591.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@47591.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@47591.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@47591.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@47599.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@47599.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@47599.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@47599.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@47599.4]
  wire  x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_clock; // @[sm_x554_outr_UnitPipe.scala 76:24:@47629.4]
  wire  x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_reset; // @[sm_x554_outr_UnitPipe.scala 76:24:@47629.4]
  wire  x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x289_TVALID; // @[sm_x554_outr_UnitPipe.scala 76:24:@47629.4]
  wire  x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x289_TREADY; // @[sm_x554_outr_UnitPipe.scala 76:24:@47629.4]
  wire [255:0] x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x289_TDATA; // @[sm_x554_outr_UnitPipe.scala 76:24:@47629.4]
  wire [7:0] x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x289_TID; // @[sm_x554_outr_UnitPipe.scala 76:24:@47629.4]
  wire [7:0] x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x289_TDEST; // @[sm_x554_outr_UnitPipe.scala 76:24:@47629.4]
  wire  x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x290_TVALID; // @[sm_x554_outr_UnitPipe.scala 76:24:@47629.4]
  wire  x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x290_TREADY; // @[sm_x554_outr_UnitPipe.scala 76:24:@47629.4]
  wire [255:0] x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x290_TDATA; // @[sm_x554_outr_UnitPipe.scala 76:24:@47629.4]
  wire  x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x554_outr_UnitPipe.scala 76:24:@47629.4]
  wire  x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x554_outr_UnitPipe.scala 76:24:@47629.4]
  wire  x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x554_outr_UnitPipe.scala 76:24:@47629.4]
  wire  x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_rr; // @[sm_x554_outr_UnitPipe.scala 76:24:@47629.4]
  wire  _T_254; // @[package.scala 96:25:@47318.4 package.scala 96:25:@47319.4]
  wire  _T_260; // @[implicits.scala 47:10:@47322.4]
  wire  _T_261; // @[sm_x555_outr_UnitPipe.scala 70:41:@47323.4]
  wire  _T_262; // @[sm_x555_outr_UnitPipe.scala 70:78:@47324.4]
  wire  _T_263; // @[sm_x555_outr_UnitPipe.scala 70:76:@47325.4]
  wire  _T_275; // @[package.scala 96:25:@47364.4 package.scala 96:25:@47365.4]
  wire  _T_281; // @[package.scala 96:25:@47372.4 package.scala 96:25:@47373.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@47375.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@47384.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@47385.4]
  wire  _T_354; // @[package.scala 100:49:@47562.4]
  reg  _T_357; // @[package.scala 48:56:@47563.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@47596.4 package.scala 96:25:@47597.4]
  wire  _T_377; // @[package.scala 96:25:@47604.4 package.scala 96:25:@47605.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@47607.4]
  x292_fifoinraw_0 x292_fifoinraw_0 ( // @[m_x292_fifoinraw_0.scala 27:17:@47153.4]
    .clock(x292_fifoinraw_0_clock),
    .reset(x292_fifoinraw_0_reset)
  );
  x293_fifoinpacked_0 x293_fifoinpacked_0 ( // @[m_x293_fifoinpacked_0.scala 27:17:@47177.4]
    .clock(x293_fifoinpacked_0_clock),
    .reset(x293_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x293_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x293_fifoinpacked_0_io_full),
    .io_active_0_in(x293_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x293_fifoinpacked_0_io_active_0_out)
  );
  x292_fifoinraw_0 x294_fifooutraw_0 ( // @[m_x294_fifooutraw_0.scala 27:17:@47201.4]
    .clock(x294_fifooutraw_0_clock),
    .reset(x294_fifooutraw_0_reset)
  );
  x297_ctrchain x297_ctrchain ( // @[SpatialBlocks.scala 37:22:@47225.4]
    .clock(x297_ctrchain_clock),
    .reset(x297_ctrchain_reset),
    .io_input_reset(x297_ctrchain_io_input_reset),
    .io_input_enable(x297_ctrchain_io_input_enable),
    .io_output_counts_1(x297_ctrchain_io_output_counts_1),
    .io_output_counts_0(x297_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x297_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x297_ctrchain_io_output_oobs_1),
    .io_output_done(x297_ctrchain_io_output_done)
  );
  x323_inr_Foreach_sm x323_inr_Foreach_sm ( // @[sm_x323_inr_Foreach.scala 32:18:@47285.4]
    .clock(x323_inr_Foreach_sm_clock),
    .reset(x323_inr_Foreach_sm_reset),
    .io_enable(x323_inr_Foreach_sm_io_enable),
    .io_done(x323_inr_Foreach_sm_io_done),
    .io_doneLatch(x323_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x323_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x323_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x323_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x323_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x323_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x323_inr_Foreach_sm_io_backpressure),
    .io_break(x323_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@47313.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@47359.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@47367.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x323_inr_Foreach_kernelx323_inr_Foreach_concrete1 x323_inr_Foreach_kernelx323_inr_Foreach_concrete1 ( // @[sm_x323_inr_Foreach.scala 126:24:@47402.4]
    .clock(x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_clock),
    .reset(x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_reset),
    .io_in_x293_fifoinpacked_0_wPort_0_en_0(x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_in_x293_fifoinpacked_0_wPort_0_en_0),
    .io_in_x293_fifoinpacked_0_full(x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_in_x293_fifoinpacked_0_full),
    .io_in_x293_fifoinpacked_0_active_0_in(x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_in_x293_fifoinpacked_0_active_0_in),
    .io_in_x293_fifoinpacked_0_active_0_out(x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_in_x293_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x554_outr_UnitPipe_sm ( // @[sm_x554_outr_UnitPipe.scala 32:18:@47534.4]
    .clock(x554_outr_UnitPipe_sm_clock),
    .reset(x554_outr_UnitPipe_sm_reset),
    .io_enable(x554_outr_UnitPipe_sm_io_enable),
    .io_done(x554_outr_UnitPipe_sm_io_done),
    .io_rst(x554_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x554_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x554_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x554_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x554_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x554_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x554_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@47591.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@47599.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1 x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1 ( // @[sm_x554_outr_UnitPipe.scala 76:24:@47629.4]
    .clock(x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_clock),
    .reset(x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_reset),
    .io_in_x289_TVALID(x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x289_TVALID),
    .io_in_x289_TREADY(x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x289_TREADY),
    .io_in_x289_TDATA(x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x289_TDATA),
    .io_in_x289_TID(x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x289_TID),
    .io_in_x289_TDEST(x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x289_TDEST),
    .io_in_x290_TVALID(x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x290_TVALID),
    .io_in_x290_TREADY(x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x290_TREADY),
    .io_in_x290_TDATA(x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x290_TDATA),
    .io_sigsIn_smEnableOuts_0(x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@47318.4 package.scala 96:25:@47319.4]
  assign _T_260 = x293_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@47322.4]
  assign _T_261 = ~ _T_260; // @[sm_x555_outr_UnitPipe.scala 70:41:@47323.4]
  assign _T_262 = ~ x293_fifoinpacked_0_io_active_0_out; // @[sm_x555_outr_UnitPipe.scala 70:78:@47324.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x555_outr_UnitPipe.scala 70:76:@47325.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@47364.4 package.scala 96:25:@47365.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@47372.4 package.scala 96:25:@47373.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@47375.4]
  assign _T_286 = x323_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@47384.4]
  assign _T_287 = ~ x323_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@47385.4]
  assign _T_354 = x554_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@47562.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@47596.4 package.scala 96:25:@47597.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@47604.4 package.scala 96:25:@47605.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@47607.4]
  assign io_in_x289_TREADY = x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x289_TREADY; // @[sm_x554_outr_UnitPipe.scala 48:23:@47685.4]
  assign io_in_x290_TVALID = x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x290_TVALID; // @[sm_x554_outr_UnitPipe.scala 49:23:@47695.4]
  assign io_in_x290_TDATA = x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x290_TDATA; // @[sm_x554_outr_UnitPipe.scala 49:23:@47693.4]
  assign io_sigsOut_smDoneIn_0 = x323_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@47382.4]
  assign io_sigsOut_smDoneIn_1 = x554_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@47614.4]
  assign io_sigsOut_smCtrCopyDone_0 = x323_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@47401.4]
  assign io_sigsOut_smCtrCopyDone_1 = x554_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@47628.4]
  assign x292_fifoinraw_0_clock = clock; // @[:@47154.4]
  assign x292_fifoinraw_0_reset = reset; // @[:@47155.4]
  assign x293_fifoinpacked_0_clock = clock; // @[:@47178.4]
  assign x293_fifoinpacked_0_reset = reset; // @[:@47179.4]
  assign x293_fifoinpacked_0_io_wPort_0_en_0 = x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_in_x293_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@47462.4]
  assign x293_fifoinpacked_0_io_active_0_in = x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_in_x293_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@47461.4]
  assign x294_fifooutraw_0_clock = clock; // @[:@47202.4]
  assign x294_fifooutraw_0_reset = reset; // @[:@47203.4]
  assign x297_ctrchain_clock = clock; // @[:@47226.4]
  assign x297_ctrchain_reset = reset; // @[:@47227.4]
  assign x297_ctrchain_io_input_reset = x323_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@47400.4]
  assign x297_ctrchain_io_input_enable = x323_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@47352.4 SpatialBlocks.scala 159:42:@47399.4]
  assign x323_inr_Foreach_sm_clock = clock; // @[:@47286.4]
  assign x323_inr_Foreach_sm_reset = reset; // @[:@47287.4]
  assign x323_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@47379.4]
  assign x323_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x555_outr_UnitPipe.scala 69:38:@47321.4]
  assign x323_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@47381.4]
  assign x323_inr_Foreach_sm_io_backpressure = _T_263 | x323_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@47353.4]
  assign x323_inr_Foreach_sm_io_break = 1'h0; // @[sm_x555_outr_UnitPipe.scala 73:36:@47331.4]
  assign RetimeWrapper_clock = clock; // @[:@47314.4]
  assign RetimeWrapper_reset = reset; // @[:@47315.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@47317.4]
  assign RetimeWrapper_io_in = x297_ctrchain_io_output_done; // @[package.scala 94:16:@47316.4]
  assign RetimeWrapper_1_clock = clock; // @[:@47360.4]
  assign RetimeWrapper_1_reset = reset; // @[:@47361.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@47363.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@47362.4]
  assign RetimeWrapper_2_clock = clock; // @[:@47368.4]
  assign RetimeWrapper_2_reset = reset; // @[:@47369.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@47371.4]
  assign RetimeWrapper_2_io_in = x323_inr_Foreach_sm_io_done; // @[package.scala 94:16:@47370.4]
  assign x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_clock = clock; // @[:@47403.4]
  assign x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_reset = reset; // @[:@47404.4]
  assign x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_in_x293_fifoinpacked_0_full = x293_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@47456.4]
  assign x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_in_x293_fifoinpacked_0_active_0_out = x293_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@47455.4]
  assign x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x323_inr_Foreach_sm_io_doneLatch; // @[sm_x323_inr_Foreach.scala 131:22:@47485.4]
  assign x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x323_inr_Foreach.scala 131:22:@47483.4]
  assign x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_break = x323_inr_Foreach_sm_io_break; // @[sm_x323_inr_Foreach.scala 131:22:@47481.4]
  assign x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x297_ctrchain_io_output_counts_1[12]}},x297_ctrchain_io_output_counts_1}; // @[sm_x323_inr_Foreach.scala 131:22:@47476.4]
  assign x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x297_ctrchain_io_output_counts_0[12]}},x297_ctrchain_io_output_counts_0}; // @[sm_x323_inr_Foreach.scala 131:22:@47475.4]
  assign x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x297_ctrchain_io_output_oobs_0; // @[sm_x323_inr_Foreach.scala 131:22:@47473.4]
  assign x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x297_ctrchain_io_output_oobs_1; // @[sm_x323_inr_Foreach.scala 131:22:@47474.4]
  assign x323_inr_Foreach_kernelx323_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x323_inr_Foreach.scala 130:18:@47469.4]
  assign x554_outr_UnitPipe_sm_clock = clock; // @[:@47535.4]
  assign x554_outr_UnitPipe_sm_reset = reset; // @[:@47536.4]
  assign x554_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@47611.4]
  assign x554_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@47586.4]
  assign x554_outr_UnitPipe_sm_io_ctrDone = x554_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x555_outr_UnitPipe.scala 78:40:@47566.4]
  assign x554_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@47613.4]
  assign x554_outr_UnitPipe_sm_io_doneIn_0 = x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@47583.4]
  assign RetimeWrapper_3_clock = clock; // @[:@47592.4]
  assign RetimeWrapper_3_reset = reset; // @[:@47593.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@47595.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@47594.4]
  assign RetimeWrapper_4_clock = clock; // @[:@47600.4]
  assign RetimeWrapper_4_reset = reset; // @[:@47601.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@47603.4]
  assign RetimeWrapper_4_io_in = x554_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@47602.4]
  assign x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_clock = clock; // @[:@47630.4]
  assign x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_reset = reset; // @[:@47631.4]
  assign x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x289_TVALID = io_in_x289_TVALID; // @[sm_x554_outr_UnitPipe.scala 48:23:@47686.4]
  assign x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x289_TDATA = io_in_x289_TDATA; // @[sm_x554_outr_UnitPipe.scala 48:23:@47684.4]
  assign x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x289_TID = io_in_x289_TID; // @[sm_x554_outr_UnitPipe.scala 48:23:@47680.4]
  assign x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x289_TDEST = io_in_x289_TDEST; // @[sm_x554_outr_UnitPipe.scala 48:23:@47679.4]
  assign x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_in_x290_TREADY = io_in_x290_TREADY; // @[sm_x554_outr_UnitPipe.scala 49:23:@47694.4]
  assign x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x554_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x554_outr_UnitPipe.scala 81:22:@47704.4]
  assign x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x554_outr_UnitPipe_sm_io_childAck_0; // @[sm_x554_outr_UnitPipe.scala 81:22:@47702.4]
  assign x554_outr_UnitPipe_kernelx554_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x554_outr_UnitPipe.scala 80:18:@47696.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x577_outr_UnitPipe_sm( // @[:@48193.2]
  input   clock, // @[:@48194.4]
  input   reset, // @[:@48195.4]
  input   io_enable, // @[:@48196.4]
  output  io_done, // @[:@48196.4]
  input   io_parentAck, // @[:@48196.4]
  input   io_doneIn_0, // @[:@48196.4]
  input   io_doneIn_1, // @[:@48196.4]
  input   io_doneIn_2, // @[:@48196.4]
  output  io_enableOut_0, // @[:@48196.4]
  output  io_enableOut_1, // @[:@48196.4]
  output  io_enableOut_2, // @[:@48196.4]
  output  io_childAck_0, // @[:@48196.4]
  output  io_childAck_1, // @[:@48196.4]
  output  io_childAck_2, // @[:@48196.4]
  input   io_ctrCopyDone_0, // @[:@48196.4]
  input   io_ctrCopyDone_1, // @[:@48196.4]
  input   io_ctrCopyDone_2 // @[:@48196.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@48199.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@48199.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@48199.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@48199.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@48199.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@48199.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@48202.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@48202.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@48202.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@48202.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@48202.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@48202.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@48205.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@48205.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@48205.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@48205.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@48205.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@48205.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@48208.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@48208.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@48208.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@48208.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@48208.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@48208.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@48211.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@48211.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@48211.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@48211.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@48211.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@48211.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@48214.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@48214.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@48214.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@48214.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@48214.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@48214.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@48255.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@48255.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@48255.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@48255.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@48255.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@48255.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@48258.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@48258.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@48258.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@48258.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@48258.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@48258.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@48261.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@48261.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@48261.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@48261.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@48261.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@48261.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@48312.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@48312.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@48312.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@48312.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@48312.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@48326.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@48326.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@48326.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@48326.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@48326.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@48344.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@48344.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@48344.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@48344.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@48344.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@48381.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@48381.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@48381.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@48381.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@48381.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@48395.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@48395.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@48395.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@48395.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@48395.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@48413.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@48413.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@48413.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@48413.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@48413.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@48450.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@48450.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@48450.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@48450.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@48450.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@48464.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@48464.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@48464.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@48464.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@48464.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@48482.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@48482.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@48482.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@48482.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@48482.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@48539.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@48539.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@48539.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@48539.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@48539.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@48556.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@48556.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@48556.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@48556.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@48556.4]
  wire  _T_77; // @[Controllers.scala 80:47:@48217.4]
  wire  allDone; // @[Controllers.scala 80:47:@48218.4]
  wire  _T_151; // @[Controllers.scala 165:35:@48296.4]
  wire  _T_153; // @[Controllers.scala 165:60:@48297.4]
  wire  _T_154; // @[Controllers.scala 165:58:@48298.4]
  wire  _T_156; // @[Controllers.scala 165:76:@48299.4]
  wire  _T_157; // @[Controllers.scala 165:74:@48300.4]
  wire  _T_161; // @[Controllers.scala 165:109:@48303.4]
  wire  _T_164; // @[Controllers.scala 165:141:@48305.4]
  wire  _T_172; // @[package.scala 96:25:@48317.4 package.scala 96:25:@48318.4]
  wire  _T_176; // @[Controllers.scala 167:54:@48320.4]
  wire  _T_177; // @[Controllers.scala 167:52:@48321.4]
  wire  _T_184; // @[package.scala 96:25:@48331.4 package.scala 96:25:@48332.4]
  wire  _T_202; // @[package.scala 96:25:@48349.4 package.scala 96:25:@48350.4]
  wire  _T_206; // @[Controllers.scala 169:67:@48352.4]
  wire  _T_207; // @[Controllers.scala 169:86:@48353.4]
  wire  _T_219; // @[Controllers.scala 165:35:@48365.4]
  wire  _T_221; // @[Controllers.scala 165:60:@48366.4]
  wire  _T_222; // @[Controllers.scala 165:58:@48367.4]
  wire  _T_224; // @[Controllers.scala 165:76:@48368.4]
  wire  _T_225; // @[Controllers.scala 165:74:@48369.4]
  wire  _T_229; // @[Controllers.scala 165:109:@48372.4]
  wire  _T_232; // @[Controllers.scala 165:141:@48374.4]
  wire  _T_240; // @[package.scala 96:25:@48386.4 package.scala 96:25:@48387.4]
  wire  _T_244; // @[Controllers.scala 167:54:@48389.4]
  wire  _T_245; // @[Controllers.scala 167:52:@48390.4]
  wire  _T_252; // @[package.scala 96:25:@48400.4 package.scala 96:25:@48401.4]
  wire  _T_270; // @[package.scala 96:25:@48418.4 package.scala 96:25:@48419.4]
  wire  _T_274; // @[Controllers.scala 169:67:@48421.4]
  wire  _T_275; // @[Controllers.scala 169:86:@48422.4]
  wire  _T_287; // @[Controllers.scala 165:35:@48434.4]
  wire  _T_289; // @[Controllers.scala 165:60:@48435.4]
  wire  _T_290; // @[Controllers.scala 165:58:@48436.4]
  wire  _T_292; // @[Controllers.scala 165:76:@48437.4]
  wire  _T_293; // @[Controllers.scala 165:74:@48438.4]
  wire  _T_297; // @[Controllers.scala 165:109:@48441.4]
  wire  _T_300; // @[Controllers.scala 165:141:@48443.4]
  wire  _T_308; // @[package.scala 96:25:@48455.4 package.scala 96:25:@48456.4]
  wire  _T_312; // @[Controllers.scala 167:54:@48458.4]
  wire  _T_313; // @[Controllers.scala 167:52:@48459.4]
  wire  _T_320; // @[package.scala 96:25:@48469.4 package.scala 96:25:@48470.4]
  wire  _T_338; // @[package.scala 96:25:@48487.4 package.scala 96:25:@48488.4]
  wire  _T_342; // @[Controllers.scala 169:67:@48490.4]
  wire  _T_343; // @[Controllers.scala 169:86:@48491.4]
  wire  _T_358; // @[Controllers.scala 213:68:@48509.4]
  wire  _T_360; // @[Controllers.scala 213:90:@48511.4]
  wire  _T_362; // @[Controllers.scala 213:132:@48513.4]
  wire  _T_366; // @[Controllers.scala 213:68:@48518.4]
  wire  _T_368; // @[Controllers.scala 213:90:@48520.4]
  wire  _T_374; // @[Controllers.scala 213:68:@48526.4]
  wire  _T_376; // @[Controllers.scala 213:90:@48528.4]
  wire  _T_383; // @[package.scala 100:49:@48534.4]
  reg  _T_386; // @[package.scala 48:56:@48535.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@48537.4]
  reg  _T_400; // @[package.scala 48:56:@48553.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@48199.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@48202.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@48205.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@48208.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@48211.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@48214.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@48255.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@48258.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@48261.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@48312.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@48326.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@48344.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@48381.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@48395.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@48413.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@48450.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@48464.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@48482.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@48539.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@48556.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@48217.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@48218.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@48296.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@48297.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@48298.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@48299.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@48300.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@48303.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@48305.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@48317.4 package.scala 96:25:@48318.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@48320.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@48321.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@48331.4 package.scala 96:25:@48332.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@48349.4 package.scala 96:25:@48350.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@48352.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@48353.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@48365.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@48366.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@48367.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@48368.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@48369.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@48372.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@48374.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@48386.4 package.scala 96:25:@48387.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@48389.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@48390.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@48400.4 package.scala 96:25:@48401.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@48418.4 package.scala 96:25:@48419.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@48421.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@48422.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@48434.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@48435.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@48436.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@48437.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@48438.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@48441.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@48443.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@48455.4 package.scala 96:25:@48456.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@48458.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@48459.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@48469.4 package.scala 96:25:@48470.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@48487.4 package.scala 96:25:@48488.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@48490.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@48491.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@48509.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@48511.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@48513.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@48518.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@48520.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@48526.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@48528.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@48534.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@48537.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@48563.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@48517.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@48525.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@48533.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@48504.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@48506.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@48508.4]
  assign active_0_clock = clock; // @[:@48200.4]
  assign active_0_reset = reset; // @[:@48201.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@48307.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@48311.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@48221.4]
  assign active_1_clock = clock; // @[:@48203.4]
  assign active_1_reset = reset; // @[:@48204.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@48376.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@48380.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@48222.4]
  assign active_2_clock = clock; // @[:@48206.4]
  assign active_2_reset = reset; // @[:@48207.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@48445.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@48449.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@48223.4]
  assign done_0_clock = clock; // @[:@48209.4]
  assign done_0_reset = reset; // @[:@48210.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@48357.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@48235.4 Controllers.scala 170:32:@48364.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@48224.4]
  assign done_1_clock = clock; // @[:@48212.4]
  assign done_1_reset = reset; // @[:@48213.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@48426.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@48244.4 Controllers.scala 170:32:@48433.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@48225.4]
  assign done_2_clock = clock; // @[:@48215.4]
  assign done_2_reset = reset; // @[:@48216.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@48495.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@48253.4 Controllers.scala 170:32:@48502.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@48226.4]
  assign iterDone_0_clock = clock; // @[:@48256.4]
  assign iterDone_0_reset = reset; // @[:@48257.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@48325.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@48275.4 Controllers.scala 168:36:@48341.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@48264.4]
  assign iterDone_1_clock = clock; // @[:@48259.4]
  assign iterDone_1_reset = reset; // @[:@48260.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@48394.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@48284.4 Controllers.scala 168:36:@48410.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@48265.4]
  assign iterDone_2_clock = clock; // @[:@48262.4]
  assign iterDone_2_reset = reset; // @[:@48263.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@48463.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@48293.4 Controllers.scala 168:36:@48479.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@48266.4]
  assign RetimeWrapper_clock = clock; // @[:@48313.4]
  assign RetimeWrapper_reset = reset; // @[:@48314.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@48316.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@48315.4]
  assign RetimeWrapper_1_clock = clock; // @[:@48327.4]
  assign RetimeWrapper_1_reset = reset; // @[:@48328.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@48330.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@48329.4]
  assign RetimeWrapper_2_clock = clock; // @[:@48345.4]
  assign RetimeWrapper_2_reset = reset; // @[:@48346.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@48348.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@48347.4]
  assign RetimeWrapper_3_clock = clock; // @[:@48382.4]
  assign RetimeWrapper_3_reset = reset; // @[:@48383.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@48385.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@48384.4]
  assign RetimeWrapper_4_clock = clock; // @[:@48396.4]
  assign RetimeWrapper_4_reset = reset; // @[:@48397.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@48399.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@48398.4]
  assign RetimeWrapper_5_clock = clock; // @[:@48414.4]
  assign RetimeWrapper_5_reset = reset; // @[:@48415.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@48417.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@48416.4]
  assign RetimeWrapper_6_clock = clock; // @[:@48451.4]
  assign RetimeWrapper_6_reset = reset; // @[:@48452.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@48454.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@48453.4]
  assign RetimeWrapper_7_clock = clock; // @[:@48465.4]
  assign RetimeWrapper_7_reset = reset; // @[:@48466.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@48468.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@48467.4]
  assign RetimeWrapper_8_clock = clock; // @[:@48483.4]
  assign RetimeWrapper_8_reset = reset; // @[:@48484.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@48486.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@48485.4]
  assign RetimeWrapper_9_clock = clock; // @[:@48540.4]
  assign RetimeWrapper_9_reset = reset; // @[:@48541.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@48543.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@48542.4]
  assign RetimeWrapper_10_clock = clock; // @[:@48557.4]
  assign RetimeWrapper_10_reset = reset; // @[:@48558.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@48560.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@48559.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x563_inr_UnitPipe_sm( // @[:@48736.2]
  input   clock, // @[:@48737.4]
  input   reset, // @[:@48738.4]
  input   io_enable, // @[:@48739.4]
  output  io_done, // @[:@48739.4]
  output  io_doneLatch, // @[:@48739.4]
  input   io_ctrDone, // @[:@48739.4]
  output  io_datapathEn, // @[:@48739.4]
  output  io_ctrInc, // @[:@48739.4]
  input   io_parentAck, // @[:@48739.4]
  input   io_backpressure // @[:@48739.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@48741.4]
  wire  active_reset; // @[Controllers.scala 261:22:@48741.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@48741.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@48741.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@48741.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@48741.4]
  wire  done_clock; // @[Controllers.scala 262:20:@48744.4]
  wire  done_reset; // @[Controllers.scala 262:20:@48744.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@48744.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@48744.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@48744.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@48744.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@48798.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@48798.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@48798.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@48798.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@48798.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@48806.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@48806.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@48806.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@48806.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@48806.4]
  wire  _T_80; // @[Controllers.scala 264:48:@48749.4]
  wire  _T_81; // @[Controllers.scala 264:46:@48750.4]
  wire  _T_82; // @[Controllers.scala 264:62:@48751.4]
  wire  _T_83; // @[Controllers.scala 264:60:@48752.4]
  wire  _T_100; // @[package.scala 100:49:@48769.4]
  reg  _T_103; // @[package.scala 48:56:@48770.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@48778.4]
  wire  _T_116; // @[Controllers.scala 283:41:@48786.4]
  wire  _T_117; // @[Controllers.scala 283:59:@48787.4]
  wire  _T_119; // @[Controllers.scala 284:37:@48790.4]
  reg  _T_125; // @[package.scala 48:56:@48794.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@48816.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@48819.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@48821.4]
  wire  _T_152; // @[Controllers.scala 292:61:@48822.4]
  wire  _T_153; // @[Controllers.scala 292:24:@48823.4]
  SRFF active ( // @[Controllers.scala 261:22:@48741.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@48744.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@48798.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@48806.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@48749.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@48750.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@48751.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@48752.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@48769.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@48778.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@48786.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@48787.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@48790.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@48821.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@48822.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@48823.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@48797.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@48825.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@48789.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@48792.4]
  assign active_clock = clock; // @[:@48742.4]
  assign active_reset = reset; // @[:@48743.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@48754.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@48758.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@48759.4]
  assign done_clock = clock; // @[:@48745.4]
  assign done_reset = reset; // @[:@48746.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@48774.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@48767.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@48768.4]
  assign RetimeWrapper_clock = clock; // @[:@48799.4]
  assign RetimeWrapper_reset = reset; // @[:@48800.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@48802.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@48801.4]
  assign RetimeWrapper_1_clock = clock; // @[:@48807.4]
  assign RetimeWrapper_1_reset = reset; // @[:@48808.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@48810.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@48809.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1( // @[:@48900.2]
  output        io_in_x556_valid, // @[:@48903.4]
  output [63:0] io_in_x556_bits_addr, // @[:@48903.4]
  output [31:0] io_in_x556_bits_size, // @[:@48903.4]
  input  [63:0] io_in_x287_outdram_number, // @[:@48903.4]
  input         io_sigsIn_backpressure, // @[:@48903.4]
  input         io_sigsIn_datapathEn, // @[:@48903.4]
  input         io_rr // @[:@48903.4]
);
  wire [96:0] x560_tuple; // @[Cat.scala 30:58:@48917.4]
  wire  _T_135; // @[implicits.scala 55:10:@48920.4]
  assign x560_tuple = {33'h7e9000,io_in_x287_outdram_number}; // @[Cat.scala 30:58:@48917.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@48920.4]
  assign io_in_x556_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x563_inr_UnitPipe.scala 65:18:@48923.4]
  assign io_in_x556_bits_addr = x560_tuple[63:0]; // @[sm_x563_inr_UnitPipe.scala 66:22:@48925.4]
  assign io_in_x556_bits_size = x560_tuple[95:64]; // @[sm_x563_inr_UnitPipe.scala 67:22:@48927.4]
endmodule
module FF_13( // @[:@48929.2]
  input         clock, // @[:@48930.4]
  input         reset, // @[:@48931.4]
  output [22:0] io_rPort_0_output_0, // @[:@48932.4]
  input  [22:0] io_wPort_0_data_0, // @[:@48932.4]
  input         io_wPort_0_reset, // @[:@48932.4]
  input         io_wPort_0_en_0 // @[:@48932.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 321:19:@48947.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 325:32:@48949.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 325:12:@48950.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@48949.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 325:12:@48950.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@48952.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@48967.2]
  input         clock, // @[:@48968.4]
  input         reset, // @[:@48969.4]
  input         io_input_reset, // @[:@48970.4]
  input         io_input_enable, // @[:@48970.4]
  output [22:0] io_output_count_0, // @[:@48970.4]
  output        io_output_oobs_0, // @[:@48970.4]
  output        io_output_done // @[:@48970.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@48983.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@48983.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@48983.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@48983.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@48983.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@48983.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@48999.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@48999.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@48999.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@48999.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@48999.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@48999.4]
  wire  _T_36; // @[Counter.scala 264:45:@49002.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@49027.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@49028.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@49029.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@49030.4]
  wire  _T_57; // @[Counter.scala 293:18:@49032.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@49040.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@49043.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@49044.4]
  wire  _T_75; // @[Counter.scala 322:102:@49048.4]
  wire  _T_77; // @[Counter.scala 322:130:@49049.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@48983.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@48999.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@49002.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@49027.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@49028.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@49029.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@49030.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@49032.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@49040.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@49043.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@49044.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@49048.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@49049.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@49047.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@49051.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@49053.4]
  assign bases_0_clock = clock; // @[:@48984.4]
  assign bases_0_reset = reset; // @[:@48985.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@49046.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@49025.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@49026.4]
  assign SRFF_clock = clock; // @[:@49000.4]
  assign SRFF_reset = reset; // @[:@49001.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@49004.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@49006.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@49007.4]
endmodule
module x565_ctrchain( // @[:@49058.2]
  input         clock, // @[:@49059.4]
  input         reset, // @[:@49060.4]
  input         io_input_reset, // @[:@49061.4]
  input         io_input_enable, // @[:@49061.4]
  output [22:0] io_output_counts_0, // @[:@49061.4]
  output        io_output_oobs_0, // @[:@49061.4]
  output        io_output_done // @[:@49061.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@49063.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@49063.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@49063.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@49063.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@49063.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@49063.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@49063.4]
  reg  wasDone; // @[Counter.scala 542:24:@49072.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@49078.4]
  wire  _T_47; // @[Counter.scala 546:80:@49079.4]
  reg  doneLatch; // @[Counter.scala 550:26:@49084.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@49085.4]
  wire  _T_55; // @[Counter.scala 551:19:@49086.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@49063.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@49078.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@49079.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@49085.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@49086.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@49088.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@49090.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@49081.4]
  assign ctrs_0_clock = clock; // @[:@49064.4]
  assign ctrs_0_reset = reset; // @[:@49065.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@49069.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@49070.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x572_inr_Foreach_sm( // @[:@49278.2]
  input   clock, // @[:@49279.4]
  input   reset, // @[:@49280.4]
  input   io_enable, // @[:@49281.4]
  output  io_done, // @[:@49281.4]
  output  io_doneLatch, // @[:@49281.4]
  input   io_ctrDone, // @[:@49281.4]
  output  io_datapathEn, // @[:@49281.4]
  output  io_ctrInc, // @[:@49281.4]
  output  io_ctrRst, // @[:@49281.4]
  input   io_parentAck, // @[:@49281.4]
  input   io_backpressure, // @[:@49281.4]
  input   io_break // @[:@49281.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@49283.4]
  wire  active_reset; // @[Controllers.scala 261:22:@49283.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@49283.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@49283.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@49283.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@49283.4]
  wire  done_clock; // @[Controllers.scala 262:20:@49286.4]
  wire  done_reset; // @[Controllers.scala 262:20:@49286.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@49286.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@49286.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@49286.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@49286.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@49320.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@49320.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@49320.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@49320.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@49320.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@49342.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@49342.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@49342.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@49342.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@49342.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@49354.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@49354.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@49354.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@49354.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@49354.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@49362.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@49362.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@49362.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@49362.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@49362.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@49378.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@49378.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@49378.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@49378.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@49378.4]
  wire  _T_80; // @[Controllers.scala 264:48:@49291.4]
  wire  _T_81; // @[Controllers.scala 264:46:@49292.4]
  wire  _T_82; // @[Controllers.scala 264:62:@49293.4]
  wire  _T_83; // @[Controllers.scala 264:60:@49294.4]
  wire  _T_100; // @[package.scala 100:49:@49311.4]
  reg  _T_103; // @[package.scala 48:56:@49312.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@49325.4 package.scala 96:25:@49326.4]
  wire  _T_110; // @[package.scala 100:49:@49327.4]
  reg  _T_113; // @[package.scala 48:56:@49328.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@49330.4]
  wire  _T_118; // @[Controllers.scala 283:41:@49335.4]
  wire  _T_119; // @[Controllers.scala 283:59:@49336.4]
  wire  _T_121; // @[Controllers.scala 284:37:@49339.4]
  wire  _T_124; // @[package.scala 96:25:@49347.4 package.scala 96:25:@49348.4]
  wire  _T_126; // @[package.scala 100:49:@49349.4]
  reg  _T_129; // @[package.scala 48:56:@49350.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@49372.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@49374.4]
  reg  _T_153; // @[package.scala 48:56:@49375.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@49383.4 package.scala 96:25:@49384.4]
  wire  _T_158; // @[Controllers.scala 292:61:@49385.4]
  wire  _T_159; // @[Controllers.scala 292:24:@49386.4]
  SRFF active ( // @[Controllers.scala 261:22:@49283.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@49286.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@49320.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@49342.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@49354.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@49362.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@49378.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@49291.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@49292.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@49293.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@49294.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@49311.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@49325.4 package.scala 96:25:@49326.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@49327.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@49330.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@49335.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@49336.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@49339.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@49347.4 package.scala 96:25:@49348.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@49349.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@49374.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@49383.4 package.scala 96:25:@49384.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@49385.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@49386.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@49353.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@49388.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@49338.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@49341.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@49333.4]
  assign active_clock = clock; // @[:@49284.4]
  assign active_reset = reset; // @[:@49285.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@49296.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@49300.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@49301.4]
  assign done_clock = clock; // @[:@49287.4]
  assign done_reset = reset; // @[:@49288.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@49316.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@49309.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@49310.4]
  assign RetimeWrapper_clock = clock; // @[:@49321.4]
  assign RetimeWrapper_reset = reset; // @[:@49322.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@49324.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@49323.4]
  assign RetimeWrapper_1_clock = clock; // @[:@49343.4]
  assign RetimeWrapper_1_reset = reset; // @[:@49344.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@49346.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@49345.4]
  assign RetimeWrapper_2_clock = clock; // @[:@49355.4]
  assign RetimeWrapper_2_reset = reset; // @[:@49356.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@49358.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@49357.4]
  assign RetimeWrapper_3_clock = clock; // @[:@49363.4]
  assign RetimeWrapper_3_reset = reset; // @[:@49364.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@49366.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@49365.4]
  assign RetimeWrapper_4_clock = clock; // @[:@49379.4]
  assign RetimeWrapper_4_reset = reset; // @[:@49380.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@49382.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@49381.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x572_inr_Foreach_kernelx572_inr_Foreach_concrete1( // @[:@49595.2]
  input         clock, // @[:@49596.4]
  input         reset, // @[:@49597.4]
  output [20:0] io_in_x291_outbuf_0_rPort_0_ofs_0, // @[:@49598.4]
  output        io_in_x291_outbuf_0_rPort_0_en_0, // @[:@49598.4]
  output        io_in_x291_outbuf_0_rPort_0_backpressure, // @[:@49598.4]
  input  [31:0] io_in_x291_outbuf_0_rPort_0_output_0, // @[:@49598.4]
  output        io_in_x557_valid, // @[:@49598.4]
  output [31:0] io_in_x557_bits_wdata_0, // @[:@49598.4]
  output        io_in_x557_bits_wstrb, // @[:@49598.4]
  input         io_sigsIn_backpressure, // @[:@49598.4]
  input         io_sigsIn_datapathEn, // @[:@49598.4]
  input         io_sigsIn_break, // @[:@49598.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@49598.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@49598.4]
  input         io_rr // @[:@49598.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@49625.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@49625.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@49654.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@49654.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@49654.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@49654.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@49654.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@49663.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@49663.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@49663.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@49663.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@49663.4]
  wire  b567; // @[sm_x572_inr_Foreach.scala 62:18:@49633.4]
  wire  _T_274; // @[sm_x572_inr_Foreach.scala 67:129:@49637.4]
  wire  _T_278; // @[implicits.scala 55:10:@49640.4]
  wire  _T_279; // @[sm_x572_inr_Foreach.scala 67:146:@49641.4]
  wire [32:0] x570_tuple; // @[Cat.scala 30:58:@49651.4]
  wire  _T_290; // @[package.scala 96:25:@49668.4 package.scala 96:25:@49669.4]
  wire  _T_292; // @[implicits.scala 55:10:@49670.4]
  wire  x712_b567_D2; // @[package.scala 96:25:@49659.4 package.scala 96:25:@49660.4]
  wire  _T_293; // @[sm_x572_inr_Foreach.scala 74:112:@49671.4]
  wire [31:0] b566_number; // @[Math.scala 723:22:@49630.4 Math.scala 724:14:@49631.4]
  _ _ ( // @[Math.scala 720:24:@49625.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@49654.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@49663.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b567 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x572_inr_Foreach.scala 62:18:@49633.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x572_inr_Foreach.scala 67:129:@49637.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@49640.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x572_inr_Foreach.scala 67:146:@49641.4]
  assign x570_tuple = {1'h1,io_in_x291_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@49651.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@49668.4 package.scala 96:25:@49669.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@49670.4]
  assign x712_b567_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@49659.4 package.scala 96:25:@49660.4]
  assign _T_293 = _T_292 & x712_b567_D2; // @[sm_x572_inr_Foreach.scala 74:112:@49671.4]
  assign b566_number = __io_result; // @[Math.scala 723:22:@49630.4 Math.scala 724:14:@49631.4]
  assign io_in_x291_outbuf_0_rPort_0_ofs_0 = b566_number[20:0]; // @[MemInterfaceType.scala 107:54:@49644.4]
  assign io_in_x291_outbuf_0_rPort_0_en_0 = _T_279 & b567; // @[MemInterfaceType.scala 110:79:@49646.4]
  assign io_in_x291_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49645.4]
  assign io_in_x557_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x572_inr_Foreach.scala 74:18:@49673.4]
  assign io_in_x557_bits_wdata_0 = x570_tuple[31:0]; // @[sm_x572_inr_Foreach.scala 75:26:@49675.4]
  assign io_in_x557_bits_wstrb = x570_tuple[32]; // @[sm_x572_inr_Foreach.scala 76:23:@49677.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@49628.4]
  assign RetimeWrapper_clock = clock; // @[:@49655.4]
  assign RetimeWrapper_reset = reset; // @[:@49656.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49658.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@49657.4]
  assign RetimeWrapper_1_clock = clock; // @[:@49664.4]
  assign RetimeWrapper_1_reset = reset; // @[:@49665.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49667.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49666.4]
endmodule
module x576_inr_UnitPipe_sm( // @[:@49833.2]
  input   clock, // @[:@49834.4]
  input   reset, // @[:@49835.4]
  input   io_enable, // @[:@49836.4]
  output  io_done, // @[:@49836.4]
  output  io_doneLatch, // @[:@49836.4]
  input   io_ctrDone, // @[:@49836.4]
  output  io_datapathEn, // @[:@49836.4]
  output  io_ctrInc, // @[:@49836.4]
  input   io_parentAck // @[:@49836.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@49838.4]
  wire  active_reset; // @[Controllers.scala 261:22:@49838.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@49838.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@49838.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@49838.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@49838.4]
  wire  done_clock; // @[Controllers.scala 262:20:@49841.4]
  wire  done_reset; // @[Controllers.scala 262:20:@49841.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@49841.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@49841.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@49841.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@49841.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@49875.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@49875.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@49875.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@49875.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@49875.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@49897.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@49897.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@49897.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@49897.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@49897.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@49909.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@49909.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@49909.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@49909.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@49909.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@49917.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@49917.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@49917.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@49917.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@49917.4]
  wire  _T_80; // @[Controllers.scala 264:48:@49846.4]
  wire  _T_81; // @[Controllers.scala 264:46:@49847.4]
  wire  _T_82; // @[Controllers.scala 264:62:@49848.4]
  wire  _T_100; // @[package.scala 100:49:@49866.4]
  reg  _T_103; // @[package.scala 48:56:@49867.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@49890.4]
  wire  _T_124; // @[package.scala 96:25:@49902.4 package.scala 96:25:@49903.4]
  wire  _T_126; // @[package.scala 100:49:@49904.4]
  reg  _T_129; // @[package.scala 48:56:@49905.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@49927.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@49929.4]
  reg  _T_153; // @[package.scala 48:56:@49930.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@49932.4]
  wire  _T_156; // @[Controllers.scala 292:61:@49933.4]
  wire  _T_157; // @[Controllers.scala 292:24:@49934.4]
  SRFF active ( // @[Controllers.scala 261:22:@49838.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@49841.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@49875.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@49897.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@49909.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@49917.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@49846.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@49847.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@49848.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@49866.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@49890.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@49902.4 package.scala 96:25:@49903.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@49904.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@49929.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@49932.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@49933.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@49934.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@49908.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@49936.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@49893.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@49896.4]
  assign active_clock = clock; // @[:@49839.4]
  assign active_reset = reset; // @[:@49840.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@49851.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@49855.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@49856.4]
  assign done_clock = clock; // @[:@49842.4]
  assign done_reset = reset; // @[:@49843.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@49871.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@49864.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@49865.4]
  assign RetimeWrapper_clock = clock; // @[:@49876.4]
  assign RetimeWrapper_reset = reset; // @[:@49877.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@49879.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@49878.4]
  assign RetimeWrapper_1_clock = clock; // @[:@49898.4]
  assign RetimeWrapper_1_reset = reset; // @[:@49899.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@49901.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@49900.4]
  assign RetimeWrapper_2_clock = clock; // @[:@49910.4]
  assign RetimeWrapper_2_reset = reset; // @[:@49911.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@49913.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@49912.4]
  assign RetimeWrapper_3_clock = clock; // @[:@49918.4]
  assign RetimeWrapper_3_reset = reset; // @[:@49919.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@49921.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@49920.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x576_inr_UnitPipe_kernelx576_inr_UnitPipe_concrete1( // @[:@50011.2]
  output  io_in_x558_ready, // @[:@50014.4]
  input   io_sigsIn_datapathEn // @[:@50014.4]
);
  assign io_in_x558_ready = io_sigsIn_datapathEn; // @[sm_x576_inr_UnitPipe.scala 57:18:@50026.4]
endmodule
module x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1( // @[:@50029.2]
  input         clock, // @[:@50030.4]
  input         reset, // @[:@50031.4]
  output        io_in_x558_ready, // @[:@50032.4]
  input         io_in_x558_valid, // @[:@50032.4]
  output [20:0] io_in_x291_outbuf_0_rPort_0_ofs_0, // @[:@50032.4]
  output        io_in_x291_outbuf_0_rPort_0_en_0, // @[:@50032.4]
  output        io_in_x291_outbuf_0_rPort_0_backpressure, // @[:@50032.4]
  input  [31:0] io_in_x291_outbuf_0_rPort_0_output_0, // @[:@50032.4]
  input         io_in_x557_ready, // @[:@50032.4]
  output        io_in_x557_valid, // @[:@50032.4]
  output [31:0] io_in_x557_bits_wdata_0, // @[:@50032.4]
  output        io_in_x557_bits_wstrb, // @[:@50032.4]
  input         io_in_x556_ready, // @[:@50032.4]
  output        io_in_x556_valid, // @[:@50032.4]
  output [63:0] io_in_x556_bits_addr, // @[:@50032.4]
  output [31:0] io_in_x556_bits_size, // @[:@50032.4]
  input  [63:0] io_in_x287_outdram_number, // @[:@50032.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@50032.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@50032.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@50032.4]
  input         io_sigsIn_smChildAcks_0, // @[:@50032.4]
  input         io_sigsIn_smChildAcks_1, // @[:@50032.4]
  input         io_sigsIn_smChildAcks_2, // @[:@50032.4]
  output        io_sigsOut_smDoneIn_0, // @[:@50032.4]
  output        io_sigsOut_smDoneIn_1, // @[:@50032.4]
  output        io_sigsOut_smDoneIn_2, // @[:@50032.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@50032.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@50032.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@50032.4]
  input         io_rr // @[:@50032.4]
);
  wire  x563_inr_UnitPipe_sm_clock; // @[sm_x563_inr_UnitPipe.scala 33:18:@50099.4]
  wire  x563_inr_UnitPipe_sm_reset; // @[sm_x563_inr_UnitPipe.scala 33:18:@50099.4]
  wire  x563_inr_UnitPipe_sm_io_enable; // @[sm_x563_inr_UnitPipe.scala 33:18:@50099.4]
  wire  x563_inr_UnitPipe_sm_io_done; // @[sm_x563_inr_UnitPipe.scala 33:18:@50099.4]
  wire  x563_inr_UnitPipe_sm_io_doneLatch; // @[sm_x563_inr_UnitPipe.scala 33:18:@50099.4]
  wire  x563_inr_UnitPipe_sm_io_ctrDone; // @[sm_x563_inr_UnitPipe.scala 33:18:@50099.4]
  wire  x563_inr_UnitPipe_sm_io_datapathEn; // @[sm_x563_inr_UnitPipe.scala 33:18:@50099.4]
  wire  x563_inr_UnitPipe_sm_io_ctrInc; // @[sm_x563_inr_UnitPipe.scala 33:18:@50099.4]
  wire  x563_inr_UnitPipe_sm_io_parentAck; // @[sm_x563_inr_UnitPipe.scala 33:18:@50099.4]
  wire  x563_inr_UnitPipe_sm_io_backpressure; // @[sm_x563_inr_UnitPipe.scala 33:18:@50099.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@50156.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@50156.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@50156.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@50156.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@50156.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@50164.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@50164.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@50164.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@50164.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@50164.4]
  wire  x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_in_x556_valid; // @[sm_x563_inr_UnitPipe.scala 69:24:@50194.4]
  wire [63:0] x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_in_x556_bits_addr; // @[sm_x563_inr_UnitPipe.scala 69:24:@50194.4]
  wire [31:0] x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_in_x556_bits_size; // @[sm_x563_inr_UnitPipe.scala 69:24:@50194.4]
  wire [63:0] x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_in_x287_outdram_number; // @[sm_x563_inr_UnitPipe.scala 69:24:@50194.4]
  wire  x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x563_inr_UnitPipe.scala 69:24:@50194.4]
  wire  x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x563_inr_UnitPipe.scala 69:24:@50194.4]
  wire  x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_rr; // @[sm_x563_inr_UnitPipe.scala 69:24:@50194.4]
  wire  x565_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@50262.4]
  wire  x565_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@50262.4]
  wire  x565_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@50262.4]
  wire  x565_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@50262.4]
  wire [22:0] x565_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@50262.4]
  wire  x565_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@50262.4]
  wire  x565_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@50262.4]
  wire  x572_inr_Foreach_sm_clock; // @[sm_x572_inr_Foreach.scala 33:18:@50315.4]
  wire  x572_inr_Foreach_sm_reset; // @[sm_x572_inr_Foreach.scala 33:18:@50315.4]
  wire  x572_inr_Foreach_sm_io_enable; // @[sm_x572_inr_Foreach.scala 33:18:@50315.4]
  wire  x572_inr_Foreach_sm_io_done; // @[sm_x572_inr_Foreach.scala 33:18:@50315.4]
  wire  x572_inr_Foreach_sm_io_doneLatch; // @[sm_x572_inr_Foreach.scala 33:18:@50315.4]
  wire  x572_inr_Foreach_sm_io_ctrDone; // @[sm_x572_inr_Foreach.scala 33:18:@50315.4]
  wire  x572_inr_Foreach_sm_io_datapathEn; // @[sm_x572_inr_Foreach.scala 33:18:@50315.4]
  wire  x572_inr_Foreach_sm_io_ctrInc; // @[sm_x572_inr_Foreach.scala 33:18:@50315.4]
  wire  x572_inr_Foreach_sm_io_ctrRst; // @[sm_x572_inr_Foreach.scala 33:18:@50315.4]
  wire  x572_inr_Foreach_sm_io_parentAck; // @[sm_x572_inr_Foreach.scala 33:18:@50315.4]
  wire  x572_inr_Foreach_sm_io_backpressure; // @[sm_x572_inr_Foreach.scala 33:18:@50315.4]
  wire  x572_inr_Foreach_sm_io_break; // @[sm_x572_inr_Foreach.scala 33:18:@50315.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@50343.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@50343.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@50343.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@50343.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@50343.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@50383.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@50383.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@50383.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@50383.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@50383.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@50391.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@50391.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@50391.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@50391.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@50391.4]
  wire  x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_clock; // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
  wire  x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_reset; // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
  wire [20:0] x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x291_outbuf_0_rPort_0_ofs_0; // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
  wire  x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x291_outbuf_0_rPort_0_en_0; // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
  wire  x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x291_outbuf_0_rPort_0_backpressure; // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
  wire [31:0] x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x291_outbuf_0_rPort_0_output_0; // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
  wire  x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x557_valid; // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
  wire [31:0] x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x557_bits_wdata_0; // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
  wire  x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x557_bits_wstrb; // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
  wire  x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
  wire  x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
  wire  x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
  wire [31:0] x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
  wire  x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
  wire  x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_rr; // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
  wire  x576_inr_UnitPipe_sm_clock; // @[sm_x576_inr_UnitPipe.scala 32:18:@50546.4]
  wire  x576_inr_UnitPipe_sm_reset; // @[sm_x576_inr_UnitPipe.scala 32:18:@50546.4]
  wire  x576_inr_UnitPipe_sm_io_enable; // @[sm_x576_inr_UnitPipe.scala 32:18:@50546.4]
  wire  x576_inr_UnitPipe_sm_io_done; // @[sm_x576_inr_UnitPipe.scala 32:18:@50546.4]
  wire  x576_inr_UnitPipe_sm_io_doneLatch; // @[sm_x576_inr_UnitPipe.scala 32:18:@50546.4]
  wire  x576_inr_UnitPipe_sm_io_ctrDone; // @[sm_x576_inr_UnitPipe.scala 32:18:@50546.4]
  wire  x576_inr_UnitPipe_sm_io_datapathEn; // @[sm_x576_inr_UnitPipe.scala 32:18:@50546.4]
  wire  x576_inr_UnitPipe_sm_io_ctrInc; // @[sm_x576_inr_UnitPipe.scala 32:18:@50546.4]
  wire  x576_inr_UnitPipe_sm_io_parentAck; // @[sm_x576_inr_UnitPipe.scala 32:18:@50546.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@50603.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@50603.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@50603.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@50603.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@50603.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@50611.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@50611.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@50611.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@50611.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@50611.4]
  wire  x576_inr_UnitPipe_kernelx576_inr_UnitPipe_concrete1_io_in_x558_ready; // @[sm_x576_inr_UnitPipe.scala 60:24:@50641.4]
  wire  x576_inr_UnitPipe_kernelx576_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x576_inr_UnitPipe.scala 60:24:@50641.4]
  wire  _T_359; // @[package.scala 100:49:@50127.4]
  reg  _T_362; // @[package.scala 48:56:@50128.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@50161.4 package.scala 96:25:@50162.4]
  wire  _T_381; // @[package.scala 96:25:@50169.4 package.scala 96:25:@50170.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@50172.4]
  wire  _T_454; // @[package.scala 96:25:@50348.4 package.scala 96:25:@50349.4]
  wire  _T_468; // @[package.scala 96:25:@50388.4 package.scala 96:25:@50389.4]
  wire  _T_474; // @[package.scala 96:25:@50396.4 package.scala 96:25:@50397.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@50399.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@50408.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@50409.4]
  wire  _T_547; // @[package.scala 100:49:@50574.4]
  reg  _T_550; // @[package.scala 48:56:@50575.4]
  reg [31:0] _RAND_1;
  wire  x576_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x577_outr_UnitPipe.scala 101:55:@50581.4]
  wire  _T_563; // @[package.scala 96:25:@50608.4 package.scala 96:25:@50609.4]
  wire  _T_569; // @[package.scala 96:25:@50616.4 package.scala 96:25:@50617.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@50619.4]
  wire  x576_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@50620.4]
  x563_inr_UnitPipe_sm x563_inr_UnitPipe_sm ( // @[sm_x563_inr_UnitPipe.scala 33:18:@50099.4]
    .clock(x563_inr_UnitPipe_sm_clock),
    .reset(x563_inr_UnitPipe_sm_reset),
    .io_enable(x563_inr_UnitPipe_sm_io_enable),
    .io_done(x563_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x563_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x563_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x563_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x563_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x563_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x563_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@50156.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@50164.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1 x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1 ( // @[sm_x563_inr_UnitPipe.scala 69:24:@50194.4]
    .io_in_x556_valid(x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_in_x556_valid),
    .io_in_x556_bits_addr(x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_in_x556_bits_addr),
    .io_in_x556_bits_size(x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_in_x556_bits_size),
    .io_in_x287_outdram_number(x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_in_x287_outdram_number),
    .io_sigsIn_backpressure(x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_rr)
  );
  x565_ctrchain x565_ctrchain ( // @[SpatialBlocks.scala 37:22:@50262.4]
    .clock(x565_ctrchain_clock),
    .reset(x565_ctrchain_reset),
    .io_input_reset(x565_ctrchain_io_input_reset),
    .io_input_enable(x565_ctrchain_io_input_enable),
    .io_output_counts_0(x565_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x565_ctrchain_io_output_oobs_0),
    .io_output_done(x565_ctrchain_io_output_done)
  );
  x572_inr_Foreach_sm x572_inr_Foreach_sm ( // @[sm_x572_inr_Foreach.scala 33:18:@50315.4]
    .clock(x572_inr_Foreach_sm_clock),
    .reset(x572_inr_Foreach_sm_reset),
    .io_enable(x572_inr_Foreach_sm_io_enable),
    .io_done(x572_inr_Foreach_sm_io_done),
    .io_doneLatch(x572_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x572_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x572_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x572_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x572_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x572_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x572_inr_Foreach_sm_io_backpressure),
    .io_break(x572_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@50343.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@50383.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@50391.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x572_inr_Foreach_kernelx572_inr_Foreach_concrete1 x572_inr_Foreach_kernelx572_inr_Foreach_concrete1 ( // @[sm_x572_inr_Foreach.scala 78:24:@50426.4]
    .clock(x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_clock),
    .reset(x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_reset),
    .io_in_x291_outbuf_0_rPort_0_ofs_0(x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x291_outbuf_0_rPort_0_ofs_0),
    .io_in_x291_outbuf_0_rPort_0_en_0(x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x291_outbuf_0_rPort_0_en_0),
    .io_in_x291_outbuf_0_rPort_0_backpressure(x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x291_outbuf_0_rPort_0_backpressure),
    .io_in_x291_outbuf_0_rPort_0_output_0(x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x291_outbuf_0_rPort_0_output_0),
    .io_in_x557_valid(x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x557_valid),
    .io_in_x557_bits_wdata_0(x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x557_bits_wdata_0),
    .io_in_x557_bits_wstrb(x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x557_bits_wstrb),
    .io_sigsIn_backpressure(x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_rr)
  );
  x576_inr_UnitPipe_sm x576_inr_UnitPipe_sm ( // @[sm_x576_inr_UnitPipe.scala 32:18:@50546.4]
    .clock(x576_inr_UnitPipe_sm_clock),
    .reset(x576_inr_UnitPipe_sm_reset),
    .io_enable(x576_inr_UnitPipe_sm_io_enable),
    .io_done(x576_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x576_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x576_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x576_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x576_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x576_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@50603.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@50611.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x576_inr_UnitPipe_kernelx576_inr_UnitPipe_concrete1 x576_inr_UnitPipe_kernelx576_inr_UnitPipe_concrete1 ( // @[sm_x576_inr_UnitPipe.scala 60:24:@50641.4]
    .io_in_x558_ready(x576_inr_UnitPipe_kernelx576_inr_UnitPipe_concrete1_io_in_x558_ready),
    .io_sigsIn_datapathEn(x576_inr_UnitPipe_kernelx576_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x563_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@50127.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@50161.4 package.scala 96:25:@50162.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@50169.4 package.scala 96:25:@50170.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@50172.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@50348.4 package.scala 96:25:@50349.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@50388.4 package.scala 96:25:@50389.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@50396.4 package.scala 96:25:@50397.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@50399.4]
  assign _T_479 = x572_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@50408.4]
  assign _T_480 = ~ x572_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@50409.4]
  assign _T_547 = x576_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@50574.4]
  assign x576_inr_UnitPipe_sigsIn_forwardpressure = io_in_x558_valid | x576_inr_UnitPipe_sm_io_doneLatch; // @[sm_x577_outr_UnitPipe.scala 101:55:@50581.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@50608.4 package.scala 96:25:@50609.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@50616.4 package.scala 96:25:@50617.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@50619.4]
  assign x576_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@50620.4]
  assign io_in_x558_ready = x576_inr_UnitPipe_kernelx576_inr_UnitPipe_concrete1_io_in_x558_ready; // @[sm_x576_inr_UnitPipe.scala 46:23:@50677.4]
  assign io_in_x291_outbuf_0_rPort_0_ofs_0 = x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x291_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@50477.4]
  assign io_in_x291_outbuf_0_rPort_0_en_0 = x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x291_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@50476.4]
  assign io_in_x291_outbuf_0_rPort_0_backpressure = x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x291_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@50475.4]
  assign io_in_x557_valid = x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x557_valid; // @[sm_x572_inr_Foreach.scala 50:23:@50481.4]
  assign io_in_x557_bits_wdata_0 = x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x557_bits_wdata_0; // @[sm_x572_inr_Foreach.scala 50:23:@50480.4]
  assign io_in_x557_bits_wstrb = x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x557_bits_wstrb; // @[sm_x572_inr_Foreach.scala 50:23:@50479.4]
  assign io_in_x556_valid = x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_in_x556_valid; // @[sm_x563_inr_UnitPipe.scala 49:23:@50232.4]
  assign io_in_x556_bits_addr = x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_in_x556_bits_addr; // @[sm_x563_inr_UnitPipe.scala 49:23:@50231.4]
  assign io_in_x556_bits_size = x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_in_x556_bits_size; // @[sm_x563_inr_UnitPipe.scala 49:23:@50230.4]
  assign io_sigsOut_smDoneIn_0 = x563_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@50179.4]
  assign io_sigsOut_smDoneIn_1 = x572_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@50406.4]
  assign io_sigsOut_smDoneIn_2 = x576_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@50626.4]
  assign io_sigsOut_smCtrCopyDone_0 = x563_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@50193.4]
  assign io_sigsOut_smCtrCopyDone_1 = x572_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@50425.4]
  assign io_sigsOut_smCtrCopyDone_2 = x576_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@50640.4]
  assign x563_inr_UnitPipe_sm_clock = clock; // @[:@50100.4]
  assign x563_inr_UnitPipe_sm_reset = reset; // @[:@50101.4]
  assign x563_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@50176.4]
  assign x563_inr_UnitPipe_sm_io_ctrDone = x563_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x577_outr_UnitPipe.scala 77:39:@50131.4]
  assign x563_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@50178.4]
  assign x563_inr_UnitPipe_sm_io_backpressure = io_in_x556_ready | x563_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@50150.4]
  assign RetimeWrapper_clock = clock; // @[:@50157.4]
  assign RetimeWrapper_reset = reset; // @[:@50158.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@50160.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@50159.4]
  assign RetimeWrapper_1_clock = clock; // @[:@50165.4]
  assign RetimeWrapper_1_reset = reset; // @[:@50166.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@50168.4]
  assign RetimeWrapper_1_io_in = x563_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@50167.4]
  assign x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_in_x287_outdram_number = io_in_x287_outdram_number; // @[sm_x563_inr_UnitPipe.scala 50:31:@50234.4]
  assign x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x556_ready | x563_inr_UnitPipe_sm_io_doneLatch; // @[sm_x563_inr_UnitPipe.scala 74:22:@50249.4]
  assign x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x563_inr_UnitPipe_sm_io_datapathEn; // @[sm_x563_inr_UnitPipe.scala 74:22:@50247.4]
  assign x563_inr_UnitPipe_kernelx563_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x563_inr_UnitPipe.scala 73:18:@50235.4]
  assign x565_ctrchain_clock = clock; // @[:@50263.4]
  assign x565_ctrchain_reset = reset; // @[:@50264.4]
  assign x565_ctrchain_io_input_reset = x572_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@50424.4]
  assign x565_ctrchain_io_input_enable = x572_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@50376.4 SpatialBlocks.scala 159:42:@50423.4]
  assign x572_inr_Foreach_sm_clock = clock; // @[:@50316.4]
  assign x572_inr_Foreach_sm_reset = reset; // @[:@50317.4]
  assign x572_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@50403.4]
  assign x572_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x577_outr_UnitPipe.scala 90:38:@50351.4]
  assign x572_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@50405.4]
  assign x572_inr_Foreach_sm_io_backpressure = io_in_x557_ready | x572_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@50377.4]
  assign x572_inr_Foreach_sm_io_break = 1'h0; // @[sm_x577_outr_UnitPipe.scala 94:36:@50357.4]
  assign RetimeWrapper_2_clock = clock; // @[:@50344.4]
  assign RetimeWrapper_2_reset = reset; // @[:@50345.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@50347.4]
  assign RetimeWrapper_2_io_in = x565_ctrchain_io_output_done; // @[package.scala 94:16:@50346.4]
  assign RetimeWrapper_3_clock = clock; // @[:@50384.4]
  assign RetimeWrapper_3_reset = reset; // @[:@50385.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@50387.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@50386.4]
  assign RetimeWrapper_4_clock = clock; // @[:@50392.4]
  assign RetimeWrapper_4_reset = reset; // @[:@50393.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@50395.4]
  assign RetimeWrapper_4_io_in = x572_inr_Foreach_sm_io_done; // @[package.scala 94:16:@50394.4]
  assign x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_clock = clock; // @[:@50427.4]
  assign x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_reset = reset; // @[:@50428.4]
  assign x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_in_x291_outbuf_0_rPort_0_output_0 = io_in_x291_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@50474.4]
  assign x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x557_ready | x572_inr_Foreach_sm_io_doneLatch; // @[sm_x572_inr_Foreach.scala 83:22:@50497.4]
  assign x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x572_inr_Foreach.scala 83:22:@50495.4]
  assign x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_sigsIn_break = x572_inr_Foreach_sm_io_break; // @[sm_x572_inr_Foreach.scala 83:22:@50493.4]
  assign x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x565_ctrchain_io_output_counts_0[22]}},x565_ctrchain_io_output_counts_0}; // @[sm_x572_inr_Foreach.scala 83:22:@50488.4]
  assign x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x565_ctrchain_io_output_oobs_0; // @[sm_x572_inr_Foreach.scala 83:22:@50487.4]
  assign x572_inr_Foreach_kernelx572_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x572_inr_Foreach.scala 82:18:@50483.4]
  assign x576_inr_UnitPipe_sm_clock = clock; // @[:@50547.4]
  assign x576_inr_UnitPipe_sm_reset = reset; // @[:@50548.4]
  assign x576_inr_UnitPipe_sm_io_enable = x576_inr_UnitPipe_sigsIn_baseEn & x576_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@50623.4]
  assign x576_inr_UnitPipe_sm_io_ctrDone = x576_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x577_outr_UnitPipe.scala 99:39:@50578.4]
  assign x576_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@50625.4]
  assign RetimeWrapper_5_clock = clock; // @[:@50604.4]
  assign RetimeWrapper_5_reset = reset; // @[:@50605.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@50607.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@50606.4]
  assign RetimeWrapper_6_clock = clock; // @[:@50612.4]
  assign RetimeWrapper_6_reset = reset; // @[:@50613.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@50615.4]
  assign RetimeWrapper_6_io_in = x576_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@50614.4]
  assign x576_inr_UnitPipe_kernelx576_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x576_inr_UnitPipe_sm_io_datapathEn; // @[sm_x576_inr_UnitPipe.scala 65:22:@50690.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x632_kernelx632_concrete1( // @[:@50706.2]
  input          clock, // @[:@50707.4]
  input          reset, // @[:@50708.4]
  input          io_in_x289_TVALID, // @[:@50709.4]
  output         io_in_x289_TREADY, // @[:@50709.4]
  input  [255:0] io_in_x289_TDATA, // @[:@50709.4]
  input  [7:0]   io_in_x289_TID, // @[:@50709.4]
  input  [7:0]   io_in_x289_TDEST, // @[:@50709.4]
  output         io_in_x558_ready, // @[:@50709.4]
  input          io_in_x558_valid, // @[:@50709.4]
  output [20:0]  io_in_x291_outbuf_0_rPort_0_ofs_0, // @[:@50709.4]
  output         io_in_x291_outbuf_0_rPort_0_en_0, // @[:@50709.4]
  output         io_in_x291_outbuf_0_rPort_0_backpressure, // @[:@50709.4]
  input  [31:0]  io_in_x291_outbuf_0_rPort_0_output_0, // @[:@50709.4]
  input          io_in_x557_ready, // @[:@50709.4]
  output         io_in_x557_valid, // @[:@50709.4]
  output [31:0]  io_in_x557_bits_wdata_0, // @[:@50709.4]
  output         io_in_x557_bits_wstrb, // @[:@50709.4]
  input          io_in_x556_ready, // @[:@50709.4]
  output         io_in_x556_valid, // @[:@50709.4]
  output [63:0]  io_in_x556_bits_addr, // @[:@50709.4]
  output [31:0]  io_in_x556_bits_size, // @[:@50709.4]
  output         io_in_x290_TVALID, // @[:@50709.4]
  input          io_in_x290_TREADY, // @[:@50709.4]
  output [255:0] io_in_x290_TDATA, // @[:@50709.4]
  input  [63:0]  io_in_x287_outdram_number, // @[:@50709.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@50709.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@50709.4]
  input          io_sigsIn_smChildAcks_0, // @[:@50709.4]
  input          io_sigsIn_smChildAcks_1, // @[:@50709.4]
  output         io_sigsOut_smDoneIn_0, // @[:@50709.4]
  output         io_sigsOut_smDoneIn_1, // @[:@50709.4]
  input          io_rr // @[:@50709.4]
);
  wire  x555_outr_UnitPipe_sm_clock; // @[sm_x555_outr_UnitPipe.scala 32:18:@50782.4]
  wire  x555_outr_UnitPipe_sm_reset; // @[sm_x555_outr_UnitPipe.scala 32:18:@50782.4]
  wire  x555_outr_UnitPipe_sm_io_enable; // @[sm_x555_outr_UnitPipe.scala 32:18:@50782.4]
  wire  x555_outr_UnitPipe_sm_io_done; // @[sm_x555_outr_UnitPipe.scala 32:18:@50782.4]
  wire  x555_outr_UnitPipe_sm_io_parentAck; // @[sm_x555_outr_UnitPipe.scala 32:18:@50782.4]
  wire  x555_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x555_outr_UnitPipe.scala 32:18:@50782.4]
  wire  x555_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x555_outr_UnitPipe.scala 32:18:@50782.4]
  wire  x555_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x555_outr_UnitPipe.scala 32:18:@50782.4]
  wire  x555_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x555_outr_UnitPipe.scala 32:18:@50782.4]
  wire  x555_outr_UnitPipe_sm_io_childAck_0; // @[sm_x555_outr_UnitPipe.scala 32:18:@50782.4]
  wire  x555_outr_UnitPipe_sm_io_childAck_1; // @[sm_x555_outr_UnitPipe.scala 32:18:@50782.4]
  wire  x555_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x555_outr_UnitPipe.scala 32:18:@50782.4]
  wire  x555_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x555_outr_UnitPipe.scala 32:18:@50782.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@50844.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@50844.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@50844.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@50844.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@50844.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@50852.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@50852.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@50852.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@50852.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@50852.4]
  wire  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_clock; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_reset; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x289_TVALID; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x289_TREADY; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire [255:0] x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x289_TDATA; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire [7:0] x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x289_TID; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire [7:0] x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x289_TDEST; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x290_TVALID; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x290_TREADY; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire [255:0] x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x290_TDATA; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_rr; // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
  wire  x577_outr_UnitPipe_sm_clock; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_reset; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_io_enable; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_io_done; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_io_parentAck; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_io_childAck_0; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_io_childAck_1; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_io_childAck_2; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  x577_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@51133.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@51133.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@51133.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@51133.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@51133.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@51141.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@51141.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@51141.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@51141.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@51141.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_clock; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_reset; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x558_ready; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x558_valid; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire [20:0] x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x291_outbuf_0_rPort_0_ofs_0; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x291_outbuf_0_rPort_0_en_0; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x291_outbuf_0_rPort_0_backpressure; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire [31:0] x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x291_outbuf_0_rPort_0_output_0; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x557_ready; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x557_valid; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire [31:0] x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x557_bits_wdata_0; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x557_bits_wstrb; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x556_ready; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x556_valid; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire [63:0] x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x556_bits_addr; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire [31:0] x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x556_bits_size; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire [63:0] x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x287_outdram_number; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_rr; // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
  wire  _T_408; // @[package.scala 96:25:@50849.4 package.scala 96:25:@50850.4]
  wire  _T_414; // @[package.scala 96:25:@50857.4 package.scala 96:25:@50858.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@50860.4]
  wire  _T_508; // @[package.scala 96:25:@51138.4 package.scala 96:25:@51139.4]
  wire  _T_514; // @[package.scala 96:25:@51146.4 package.scala 96:25:@51147.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@51149.4]
  x555_outr_UnitPipe_sm x555_outr_UnitPipe_sm ( // @[sm_x555_outr_UnitPipe.scala 32:18:@50782.4]
    .clock(x555_outr_UnitPipe_sm_clock),
    .reset(x555_outr_UnitPipe_sm_reset),
    .io_enable(x555_outr_UnitPipe_sm_io_enable),
    .io_done(x555_outr_UnitPipe_sm_io_done),
    .io_parentAck(x555_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x555_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x555_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x555_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x555_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x555_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x555_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x555_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x555_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@50844.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@50852.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1 x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1 ( // @[sm_x555_outr_UnitPipe.scala 87:24:@50883.4]
    .clock(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_clock),
    .reset(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_reset),
    .io_in_x289_TVALID(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x289_TVALID),
    .io_in_x289_TREADY(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x289_TREADY),
    .io_in_x289_TDATA(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x289_TDATA),
    .io_in_x289_TID(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x289_TID),
    .io_in_x289_TDEST(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x289_TDEST),
    .io_in_x290_TVALID(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x290_TVALID),
    .io_in_x290_TREADY(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x290_TREADY),
    .io_in_x290_TDATA(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x290_TDATA),
    .io_sigsIn_smEnableOuts_0(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_rr)
  );
  x577_outr_UnitPipe_sm x577_outr_UnitPipe_sm ( // @[sm_x577_outr_UnitPipe.scala 36:18:@51061.4]
    .clock(x577_outr_UnitPipe_sm_clock),
    .reset(x577_outr_UnitPipe_sm_reset),
    .io_enable(x577_outr_UnitPipe_sm_io_enable),
    .io_done(x577_outr_UnitPipe_sm_io_done),
    .io_parentAck(x577_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x577_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x577_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x577_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x577_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x577_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x577_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x577_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x577_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x577_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x577_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x577_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x577_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@51133.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@51141.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1 x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1 ( // @[sm_x577_outr_UnitPipe.scala 108:24:@51173.4]
    .clock(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_clock),
    .reset(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_reset),
    .io_in_x558_ready(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x558_ready),
    .io_in_x558_valid(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x558_valid),
    .io_in_x291_outbuf_0_rPort_0_ofs_0(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x291_outbuf_0_rPort_0_ofs_0),
    .io_in_x291_outbuf_0_rPort_0_en_0(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x291_outbuf_0_rPort_0_en_0),
    .io_in_x291_outbuf_0_rPort_0_backpressure(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x291_outbuf_0_rPort_0_backpressure),
    .io_in_x291_outbuf_0_rPort_0_output_0(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x291_outbuf_0_rPort_0_output_0),
    .io_in_x557_ready(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x557_ready),
    .io_in_x557_valid(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x557_valid),
    .io_in_x557_bits_wdata_0(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x557_bits_wdata_0),
    .io_in_x557_bits_wstrb(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x557_bits_wstrb),
    .io_in_x556_ready(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x556_ready),
    .io_in_x556_valid(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x556_valid),
    .io_in_x556_bits_addr(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x556_bits_addr),
    .io_in_x556_bits_size(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x556_bits_size),
    .io_in_x287_outdram_number(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x287_outdram_number),
    .io_sigsIn_smEnableOuts_0(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@50849.4 package.scala 96:25:@50850.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@50857.4 package.scala 96:25:@50858.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@50860.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@51138.4 package.scala 96:25:@51139.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@51146.4 package.scala 96:25:@51147.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@51149.4]
  assign io_in_x289_TREADY = x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x289_TREADY; // @[sm_x555_outr_UnitPipe.scala 48:23:@50951.4]
  assign io_in_x558_ready = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x558_ready; // @[sm_x577_outr_UnitPipe.scala 58:23:@51255.4]
  assign io_in_x291_outbuf_0_rPort_0_ofs_0 = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x291_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@51259.4]
  assign io_in_x291_outbuf_0_rPort_0_en_0 = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x291_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@51258.4]
  assign io_in_x291_outbuf_0_rPort_0_backpressure = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x291_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@51257.4]
  assign io_in_x557_valid = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x557_valid; // @[sm_x577_outr_UnitPipe.scala 60:23:@51263.4]
  assign io_in_x557_bits_wdata_0 = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x557_bits_wdata_0; // @[sm_x577_outr_UnitPipe.scala 60:23:@51262.4]
  assign io_in_x557_bits_wstrb = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x557_bits_wstrb; // @[sm_x577_outr_UnitPipe.scala 60:23:@51261.4]
  assign io_in_x556_valid = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x556_valid; // @[sm_x577_outr_UnitPipe.scala 61:23:@51267.4]
  assign io_in_x556_bits_addr = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x556_bits_addr; // @[sm_x577_outr_UnitPipe.scala 61:23:@51266.4]
  assign io_in_x556_bits_size = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x556_bits_size; // @[sm_x577_outr_UnitPipe.scala 61:23:@51265.4]
  assign io_in_x290_TVALID = x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x290_TVALID; // @[sm_x555_outr_UnitPipe.scala 49:23:@50961.4]
  assign io_in_x290_TDATA = x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x290_TDATA; // @[sm_x555_outr_UnitPipe.scala 49:23:@50959.4]
  assign io_sigsOut_smDoneIn_0 = x555_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@50867.4]
  assign io_sigsOut_smDoneIn_1 = x577_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@51156.4]
  assign x555_outr_UnitPipe_sm_clock = clock; // @[:@50783.4]
  assign x555_outr_UnitPipe_sm_reset = reset; // @[:@50784.4]
  assign x555_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@50864.4]
  assign x555_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@50866.4]
  assign x555_outr_UnitPipe_sm_io_doneIn_0 = x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@50834.4]
  assign x555_outr_UnitPipe_sm_io_doneIn_1 = x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@50835.4]
  assign x555_outr_UnitPipe_sm_io_ctrCopyDone_0 = x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@50881.4]
  assign x555_outr_UnitPipe_sm_io_ctrCopyDone_1 = x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@50882.4]
  assign RetimeWrapper_clock = clock; // @[:@50845.4]
  assign RetimeWrapper_reset = reset; // @[:@50846.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@50848.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@50847.4]
  assign RetimeWrapper_1_clock = clock; // @[:@50853.4]
  assign RetimeWrapper_1_reset = reset; // @[:@50854.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@50856.4]
  assign RetimeWrapper_1_io_in = x555_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@50855.4]
  assign x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_clock = clock; // @[:@50884.4]
  assign x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_reset = reset; // @[:@50885.4]
  assign x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x289_TVALID = io_in_x289_TVALID; // @[sm_x555_outr_UnitPipe.scala 48:23:@50952.4]
  assign x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x289_TDATA = io_in_x289_TDATA; // @[sm_x555_outr_UnitPipe.scala 48:23:@50950.4]
  assign x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x289_TID = io_in_x289_TID; // @[sm_x555_outr_UnitPipe.scala 48:23:@50946.4]
  assign x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x289_TDEST = io_in_x289_TDEST; // @[sm_x555_outr_UnitPipe.scala 48:23:@50945.4]
  assign x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_in_x290_TREADY = io_in_x290_TREADY; // @[sm_x555_outr_UnitPipe.scala 49:23:@50960.4]
  assign x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x555_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x555_outr_UnitPipe.scala 92:22:@50977.4]
  assign x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x555_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x555_outr_UnitPipe.scala 92:22:@50978.4]
  assign x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x555_outr_UnitPipe_sm_io_childAck_0; // @[sm_x555_outr_UnitPipe.scala 92:22:@50973.4]
  assign x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x555_outr_UnitPipe_sm_io_childAck_1; // @[sm_x555_outr_UnitPipe.scala 92:22:@50974.4]
  assign x555_outr_UnitPipe_kernelx555_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x555_outr_UnitPipe.scala 91:18:@50962.4]
  assign x577_outr_UnitPipe_sm_clock = clock; // @[:@51062.4]
  assign x577_outr_UnitPipe_sm_reset = reset; // @[:@51063.4]
  assign x577_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@51153.4]
  assign x577_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@51155.4]
  assign x577_outr_UnitPipe_sm_io_doneIn_0 = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@51121.4]
  assign x577_outr_UnitPipe_sm_io_doneIn_1 = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@51122.4]
  assign x577_outr_UnitPipe_sm_io_doneIn_2 = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@51123.4]
  assign x577_outr_UnitPipe_sm_io_ctrCopyDone_0 = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@51170.4]
  assign x577_outr_UnitPipe_sm_io_ctrCopyDone_1 = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@51171.4]
  assign x577_outr_UnitPipe_sm_io_ctrCopyDone_2 = x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@51172.4]
  assign RetimeWrapper_2_clock = clock; // @[:@51134.4]
  assign RetimeWrapper_2_reset = reset; // @[:@51135.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@51137.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@51136.4]
  assign RetimeWrapper_3_clock = clock; // @[:@51142.4]
  assign RetimeWrapper_3_reset = reset; // @[:@51143.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@51145.4]
  assign RetimeWrapper_3_io_in = x577_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@51144.4]
  assign x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_clock = clock; // @[:@51174.4]
  assign x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_reset = reset; // @[:@51175.4]
  assign x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x558_valid = io_in_x558_valid; // @[sm_x577_outr_UnitPipe.scala 58:23:@51254.4]
  assign x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x291_outbuf_0_rPort_0_output_0 = io_in_x291_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@51256.4]
  assign x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x557_ready = io_in_x557_ready; // @[sm_x577_outr_UnitPipe.scala 60:23:@51264.4]
  assign x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x556_ready = io_in_x556_ready; // @[sm_x577_outr_UnitPipe.scala 61:23:@51268.4]
  assign x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_in_x287_outdram_number = io_in_x287_outdram_number; // @[sm_x577_outr_UnitPipe.scala 62:31:@51269.4]
  assign x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x577_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x577_outr_UnitPipe.scala 113:22:@51292.4]
  assign x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x577_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x577_outr_UnitPipe.scala 113:22:@51293.4]
  assign x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x577_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x577_outr_UnitPipe.scala 113:22:@51294.4]
  assign x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x577_outr_UnitPipe_sm_io_childAck_0; // @[sm_x577_outr_UnitPipe.scala 113:22:@51286.4]
  assign x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x577_outr_UnitPipe_sm_io_childAck_1; // @[sm_x577_outr_UnitPipe.scala 113:22:@51287.4]
  assign x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x577_outr_UnitPipe_sm_io_childAck_2; // @[sm_x577_outr_UnitPipe.scala 113:22:@51288.4]
  assign x577_outr_UnitPipe_kernelx577_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x577_outr_UnitPipe.scala 112:18:@51270.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@51322.2]
  input          clock, // @[:@51323.4]
  input          reset, // @[:@51324.4]
  input          io_in_x289_TVALID, // @[:@51325.4]
  output         io_in_x289_TREADY, // @[:@51325.4]
  input  [255:0] io_in_x289_TDATA, // @[:@51325.4]
  input  [7:0]   io_in_x289_TID, // @[:@51325.4]
  input  [7:0]   io_in_x289_TDEST, // @[:@51325.4]
  output         io_in_x558_ready, // @[:@51325.4]
  input          io_in_x558_valid, // @[:@51325.4]
  input          io_in_x557_ready, // @[:@51325.4]
  output         io_in_x557_valid, // @[:@51325.4]
  output [31:0]  io_in_x557_bits_wdata_0, // @[:@51325.4]
  output         io_in_x557_bits_wstrb, // @[:@51325.4]
  input          io_in_x556_ready, // @[:@51325.4]
  output         io_in_x556_valid, // @[:@51325.4]
  output [63:0]  io_in_x556_bits_addr, // @[:@51325.4]
  output [31:0]  io_in_x556_bits_size, // @[:@51325.4]
  output         io_in_x290_TVALID, // @[:@51325.4]
  input          io_in_x290_TREADY, // @[:@51325.4]
  output [255:0] io_in_x290_TDATA, // @[:@51325.4]
  input  [63:0]  io_in_x287_outdram_number, // @[:@51325.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@51325.4]
  input          io_sigsIn_smChildAcks_0, // @[:@51325.4]
  output         io_sigsOut_smDoneIn_0, // @[:@51325.4]
  input          io_rr // @[:@51325.4]
);
  wire  x291_outbuf_0_clock; // @[m_x291_outbuf_0.scala 27:17:@51335.4]
  wire  x291_outbuf_0_reset; // @[m_x291_outbuf_0.scala 27:17:@51335.4]
  wire [20:0] x291_outbuf_0_io_rPort_0_ofs_0; // @[m_x291_outbuf_0.scala 27:17:@51335.4]
  wire  x291_outbuf_0_io_rPort_0_en_0; // @[m_x291_outbuf_0.scala 27:17:@51335.4]
  wire  x291_outbuf_0_io_rPort_0_backpressure; // @[m_x291_outbuf_0.scala 27:17:@51335.4]
  wire [31:0] x291_outbuf_0_io_rPort_0_output_0; // @[m_x291_outbuf_0.scala 27:17:@51335.4]
  wire  x632_sm_clock; // @[sm_x632.scala 37:18:@51393.4]
  wire  x632_sm_reset; // @[sm_x632.scala 37:18:@51393.4]
  wire  x632_sm_io_enable; // @[sm_x632.scala 37:18:@51393.4]
  wire  x632_sm_io_done; // @[sm_x632.scala 37:18:@51393.4]
  wire  x632_sm_io_ctrDone; // @[sm_x632.scala 37:18:@51393.4]
  wire  x632_sm_io_ctrInc; // @[sm_x632.scala 37:18:@51393.4]
  wire  x632_sm_io_parentAck; // @[sm_x632.scala 37:18:@51393.4]
  wire  x632_sm_io_doneIn_0; // @[sm_x632.scala 37:18:@51393.4]
  wire  x632_sm_io_doneIn_1; // @[sm_x632.scala 37:18:@51393.4]
  wire  x632_sm_io_enableOut_0; // @[sm_x632.scala 37:18:@51393.4]
  wire  x632_sm_io_enableOut_1; // @[sm_x632.scala 37:18:@51393.4]
  wire  x632_sm_io_childAck_0; // @[sm_x632.scala 37:18:@51393.4]
  wire  x632_sm_io_childAck_1; // @[sm_x632.scala 37:18:@51393.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@51460.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@51460.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@51460.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@51460.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@51460.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@51468.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@51468.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@51468.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@51468.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@51468.4]
  wire  x632_kernelx632_concrete1_clock; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_reset; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_in_x289_TVALID; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_in_x289_TREADY; // @[sm_x632.scala 102:24:@51497.4]
  wire [255:0] x632_kernelx632_concrete1_io_in_x289_TDATA; // @[sm_x632.scala 102:24:@51497.4]
  wire [7:0] x632_kernelx632_concrete1_io_in_x289_TID; // @[sm_x632.scala 102:24:@51497.4]
  wire [7:0] x632_kernelx632_concrete1_io_in_x289_TDEST; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_in_x558_ready; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_in_x558_valid; // @[sm_x632.scala 102:24:@51497.4]
  wire [20:0] x632_kernelx632_concrete1_io_in_x291_outbuf_0_rPort_0_ofs_0; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_in_x291_outbuf_0_rPort_0_en_0; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_in_x291_outbuf_0_rPort_0_backpressure; // @[sm_x632.scala 102:24:@51497.4]
  wire [31:0] x632_kernelx632_concrete1_io_in_x291_outbuf_0_rPort_0_output_0; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_in_x557_ready; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_in_x557_valid; // @[sm_x632.scala 102:24:@51497.4]
  wire [31:0] x632_kernelx632_concrete1_io_in_x557_bits_wdata_0; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_in_x557_bits_wstrb; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_in_x556_ready; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_in_x556_valid; // @[sm_x632.scala 102:24:@51497.4]
  wire [63:0] x632_kernelx632_concrete1_io_in_x556_bits_addr; // @[sm_x632.scala 102:24:@51497.4]
  wire [31:0] x632_kernelx632_concrete1_io_in_x556_bits_size; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_in_x290_TVALID; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_in_x290_TREADY; // @[sm_x632.scala 102:24:@51497.4]
  wire [255:0] x632_kernelx632_concrete1_io_in_x290_TDATA; // @[sm_x632.scala 102:24:@51497.4]
  wire [63:0] x632_kernelx632_concrete1_io_in_x287_outdram_number; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x632.scala 102:24:@51497.4]
  wire  x632_kernelx632_concrete1_io_rr; // @[sm_x632.scala 102:24:@51497.4]
  wire  _T_266; // @[package.scala 100:49:@51426.4]
  reg  _T_269; // @[package.scala 48:56:@51427.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@51465.4 package.scala 96:25:@51466.4]
  wire  _T_289; // @[package.scala 96:25:@51473.4 package.scala 96:25:@51474.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@51476.4]
  x291_outbuf_0 x291_outbuf_0 ( // @[m_x291_outbuf_0.scala 27:17:@51335.4]
    .clock(x291_outbuf_0_clock),
    .reset(x291_outbuf_0_reset),
    .io_rPort_0_ofs_0(x291_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x291_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x291_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x291_outbuf_0_io_rPort_0_output_0)
  );
  x632_sm x632_sm ( // @[sm_x632.scala 37:18:@51393.4]
    .clock(x632_sm_clock),
    .reset(x632_sm_reset),
    .io_enable(x632_sm_io_enable),
    .io_done(x632_sm_io_done),
    .io_ctrDone(x632_sm_io_ctrDone),
    .io_ctrInc(x632_sm_io_ctrInc),
    .io_parentAck(x632_sm_io_parentAck),
    .io_doneIn_0(x632_sm_io_doneIn_0),
    .io_doneIn_1(x632_sm_io_doneIn_1),
    .io_enableOut_0(x632_sm_io_enableOut_0),
    .io_enableOut_1(x632_sm_io_enableOut_1),
    .io_childAck_0(x632_sm_io_childAck_0),
    .io_childAck_1(x632_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@51460.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@51468.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x632_kernelx632_concrete1 x632_kernelx632_concrete1 ( // @[sm_x632.scala 102:24:@51497.4]
    .clock(x632_kernelx632_concrete1_clock),
    .reset(x632_kernelx632_concrete1_reset),
    .io_in_x289_TVALID(x632_kernelx632_concrete1_io_in_x289_TVALID),
    .io_in_x289_TREADY(x632_kernelx632_concrete1_io_in_x289_TREADY),
    .io_in_x289_TDATA(x632_kernelx632_concrete1_io_in_x289_TDATA),
    .io_in_x289_TID(x632_kernelx632_concrete1_io_in_x289_TID),
    .io_in_x289_TDEST(x632_kernelx632_concrete1_io_in_x289_TDEST),
    .io_in_x558_ready(x632_kernelx632_concrete1_io_in_x558_ready),
    .io_in_x558_valid(x632_kernelx632_concrete1_io_in_x558_valid),
    .io_in_x291_outbuf_0_rPort_0_ofs_0(x632_kernelx632_concrete1_io_in_x291_outbuf_0_rPort_0_ofs_0),
    .io_in_x291_outbuf_0_rPort_0_en_0(x632_kernelx632_concrete1_io_in_x291_outbuf_0_rPort_0_en_0),
    .io_in_x291_outbuf_0_rPort_0_backpressure(x632_kernelx632_concrete1_io_in_x291_outbuf_0_rPort_0_backpressure),
    .io_in_x291_outbuf_0_rPort_0_output_0(x632_kernelx632_concrete1_io_in_x291_outbuf_0_rPort_0_output_0),
    .io_in_x557_ready(x632_kernelx632_concrete1_io_in_x557_ready),
    .io_in_x557_valid(x632_kernelx632_concrete1_io_in_x557_valid),
    .io_in_x557_bits_wdata_0(x632_kernelx632_concrete1_io_in_x557_bits_wdata_0),
    .io_in_x557_bits_wstrb(x632_kernelx632_concrete1_io_in_x557_bits_wstrb),
    .io_in_x556_ready(x632_kernelx632_concrete1_io_in_x556_ready),
    .io_in_x556_valid(x632_kernelx632_concrete1_io_in_x556_valid),
    .io_in_x556_bits_addr(x632_kernelx632_concrete1_io_in_x556_bits_addr),
    .io_in_x556_bits_size(x632_kernelx632_concrete1_io_in_x556_bits_size),
    .io_in_x290_TVALID(x632_kernelx632_concrete1_io_in_x290_TVALID),
    .io_in_x290_TREADY(x632_kernelx632_concrete1_io_in_x290_TREADY),
    .io_in_x290_TDATA(x632_kernelx632_concrete1_io_in_x290_TDATA),
    .io_in_x287_outdram_number(x632_kernelx632_concrete1_io_in_x287_outdram_number),
    .io_sigsIn_smEnableOuts_0(x632_kernelx632_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x632_kernelx632_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x632_kernelx632_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x632_kernelx632_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x632_kernelx632_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x632_kernelx632_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x632_kernelx632_concrete1_io_rr)
  );
  assign _T_266 = x632_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@51426.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@51465.4 package.scala 96:25:@51466.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@51473.4 package.scala 96:25:@51474.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@51476.4]
  assign io_in_x289_TREADY = x632_kernelx632_concrete1_io_in_x289_TREADY; // @[sm_x632.scala 63:23:@51583.4]
  assign io_in_x558_ready = x632_kernelx632_concrete1_io_in_x558_ready; // @[sm_x632.scala 64:23:@51587.4]
  assign io_in_x557_valid = x632_kernelx632_concrete1_io_in_x557_valid; // @[sm_x632.scala 66:23:@51595.4]
  assign io_in_x557_bits_wdata_0 = x632_kernelx632_concrete1_io_in_x557_bits_wdata_0; // @[sm_x632.scala 66:23:@51594.4]
  assign io_in_x557_bits_wstrb = x632_kernelx632_concrete1_io_in_x557_bits_wstrb; // @[sm_x632.scala 66:23:@51593.4]
  assign io_in_x556_valid = x632_kernelx632_concrete1_io_in_x556_valid; // @[sm_x632.scala 67:23:@51599.4]
  assign io_in_x556_bits_addr = x632_kernelx632_concrete1_io_in_x556_bits_addr; // @[sm_x632.scala 67:23:@51598.4]
  assign io_in_x556_bits_size = x632_kernelx632_concrete1_io_in_x556_bits_size; // @[sm_x632.scala 67:23:@51597.4]
  assign io_in_x290_TVALID = x632_kernelx632_concrete1_io_in_x290_TVALID; // @[sm_x632.scala 68:23:@51609.4]
  assign io_in_x290_TDATA = x632_kernelx632_concrete1_io_in_x290_TDATA; // @[sm_x632.scala 68:23:@51607.4]
  assign io_sigsOut_smDoneIn_0 = x632_sm_io_done; // @[SpatialBlocks.scala 156:53:@51483.4]
  assign x291_outbuf_0_clock = clock; // @[:@51336.4]
  assign x291_outbuf_0_reset = reset; // @[:@51337.4]
  assign x291_outbuf_0_io_rPort_0_ofs_0 = x632_kernelx632_concrete1_io_in_x291_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@51591.4]
  assign x291_outbuf_0_io_rPort_0_en_0 = x632_kernelx632_concrete1_io_in_x291_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@51590.4]
  assign x291_outbuf_0_io_rPort_0_backpressure = x632_kernelx632_concrete1_io_in_x291_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@51589.4]
  assign x632_sm_clock = clock; // @[:@51394.4]
  assign x632_sm_reset = reset; // @[:@51395.4]
  assign x632_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@51480.4]
  assign x632_sm_io_ctrDone = x632_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:26:@51430.4]
  assign x632_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@51482.4]
  assign x632_sm_io_doneIn_0 = x632_kernelx632_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@51450.4]
  assign x632_sm_io_doneIn_1 = x632_kernelx632_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@51451.4]
  assign RetimeWrapper_clock = clock; // @[:@51461.4]
  assign RetimeWrapper_reset = reset; // @[:@51462.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@51464.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@51463.4]
  assign RetimeWrapper_1_clock = clock; // @[:@51469.4]
  assign RetimeWrapper_1_reset = reset; // @[:@51470.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@51472.4]
  assign RetimeWrapper_1_io_in = x632_sm_io_done; // @[package.scala 94:16:@51471.4]
  assign x632_kernelx632_concrete1_clock = clock; // @[:@51498.4]
  assign x632_kernelx632_concrete1_reset = reset; // @[:@51499.4]
  assign x632_kernelx632_concrete1_io_in_x289_TVALID = io_in_x289_TVALID; // @[sm_x632.scala 63:23:@51584.4]
  assign x632_kernelx632_concrete1_io_in_x289_TDATA = io_in_x289_TDATA; // @[sm_x632.scala 63:23:@51582.4]
  assign x632_kernelx632_concrete1_io_in_x289_TID = io_in_x289_TID; // @[sm_x632.scala 63:23:@51578.4]
  assign x632_kernelx632_concrete1_io_in_x289_TDEST = io_in_x289_TDEST; // @[sm_x632.scala 63:23:@51577.4]
  assign x632_kernelx632_concrete1_io_in_x558_valid = io_in_x558_valid; // @[sm_x632.scala 64:23:@51586.4]
  assign x632_kernelx632_concrete1_io_in_x291_outbuf_0_rPort_0_output_0 = x291_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@51588.4]
  assign x632_kernelx632_concrete1_io_in_x557_ready = io_in_x557_ready; // @[sm_x632.scala 66:23:@51596.4]
  assign x632_kernelx632_concrete1_io_in_x556_ready = io_in_x556_ready; // @[sm_x632.scala 67:23:@51600.4]
  assign x632_kernelx632_concrete1_io_in_x290_TREADY = io_in_x290_TREADY; // @[sm_x632.scala 68:23:@51608.4]
  assign x632_kernelx632_concrete1_io_in_x287_outdram_number = io_in_x287_outdram_number; // @[sm_x632.scala 69:31:@51610.4]
  assign x632_kernelx632_concrete1_io_sigsIn_smEnableOuts_0 = x632_sm_io_enableOut_0; // @[sm_x632.scala 107:22:@51621.4]
  assign x632_kernelx632_concrete1_io_sigsIn_smEnableOuts_1 = x632_sm_io_enableOut_1; // @[sm_x632.scala 107:22:@51622.4]
  assign x632_kernelx632_concrete1_io_sigsIn_smChildAcks_0 = x632_sm_io_childAck_0; // @[sm_x632.scala 107:22:@51617.4]
  assign x632_kernelx632_concrete1_io_sigsIn_smChildAcks_1 = x632_sm_io_childAck_1; // @[sm_x632.scala 107:22:@51618.4]
  assign x632_kernelx632_concrete1_io_rr = io_rr; // @[sm_x632.scala 106:18:@51611.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@51644.2]
  input          clock, // @[:@51645.4]
  input          reset, // @[:@51646.4]
  input          io_enable, // @[:@51647.4]
  output         io_done, // @[:@51647.4]
  input          io_reset, // @[:@51647.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@51647.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@51647.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@51647.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@51647.4]
  output         io_memStreams_loads_0_data_ready, // @[:@51647.4]
  input          io_memStreams_loads_0_data_valid, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@51647.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@51647.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@51647.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@51647.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@51647.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@51647.4]
  input          io_memStreams_stores_0_data_ready, // @[:@51647.4]
  output         io_memStreams_stores_0_data_valid, // @[:@51647.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@51647.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@51647.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@51647.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@51647.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@51647.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@51647.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@51647.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@51647.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@51647.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@51647.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@51647.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@51647.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@51647.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@51647.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@51647.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@51647.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@51647.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@51647.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@51647.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@51647.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@51647.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@51647.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@51647.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@51647.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@51647.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@51647.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@51647.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@51647.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@51647.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@51647.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@51647.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@51647.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@51647.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@51647.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@51647.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@51647.4]
  output         io_heap_0_req_valid, // @[:@51647.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@51647.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@51647.4]
  input          io_heap_0_resp_valid, // @[:@51647.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@51647.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@51647.4]
  input  [63:0]  io_argIns_0, // @[:@51647.4]
  input  [63:0]  io_argIns_1, // @[:@51647.4]
  input          io_argOuts_0_port_ready, // @[:@51647.4]
  output         io_argOuts_0_port_valid, // @[:@51647.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@51647.4]
  input  [63:0]  io_argOuts_0_echo // @[:@51647.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@51795.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@51795.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@51795.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@51795.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@51813.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@51813.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@51813.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@51813.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@51813.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@51822.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@51822.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@51822.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@51822.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@51822.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@51822.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@51861.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@51861.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@51861.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@51861.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@51861.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@51861.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@51861.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@51861.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@51861.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@51861.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@51861.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@51893.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@51893.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@51893.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@51893.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@51893.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_io_in_x289_TVALID; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_io_in_x289_TREADY; // @[sm_RootController.scala 91:24:@51955.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x289_TDATA; // @[sm_RootController.scala 91:24:@51955.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x289_TID; // @[sm_RootController.scala 91:24:@51955.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x289_TDEST; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_io_in_x558_ready; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_io_in_x558_valid; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_io_in_x557_ready; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_io_in_x557_valid; // @[sm_RootController.scala 91:24:@51955.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x557_bits_wdata_0; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_io_in_x557_bits_wstrb; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_io_in_x556_ready; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_io_in_x556_valid; // @[sm_RootController.scala 91:24:@51955.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x556_bits_addr; // @[sm_RootController.scala 91:24:@51955.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x556_bits_size; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_io_in_x290_TVALID; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_io_in_x290_TREADY; // @[sm_RootController.scala 91:24:@51955.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x290_TDATA; // @[sm_RootController.scala 91:24:@51955.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x287_outdram_number; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@51955.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@51955.4]
  wire  _T_599; // @[package.scala 96:25:@51818.4 package.scala 96:25:@51819.4]
  wire  _T_664; // @[Main.scala 46:50:@51889.4]
  wire  _T_665; // @[Main.scala 46:59:@51890.4]
  wire  _T_677; // @[package.scala 100:49:@51910.4]
  reg  _T_680; // @[package.scala 48:56:@51911.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@51795.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@51813.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@51822.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@51861.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@51893.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@51955.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x289_TVALID(RootController_kernelRootController_concrete1_io_in_x289_TVALID),
    .io_in_x289_TREADY(RootController_kernelRootController_concrete1_io_in_x289_TREADY),
    .io_in_x289_TDATA(RootController_kernelRootController_concrete1_io_in_x289_TDATA),
    .io_in_x289_TID(RootController_kernelRootController_concrete1_io_in_x289_TID),
    .io_in_x289_TDEST(RootController_kernelRootController_concrete1_io_in_x289_TDEST),
    .io_in_x558_ready(RootController_kernelRootController_concrete1_io_in_x558_ready),
    .io_in_x558_valid(RootController_kernelRootController_concrete1_io_in_x558_valid),
    .io_in_x557_ready(RootController_kernelRootController_concrete1_io_in_x557_ready),
    .io_in_x557_valid(RootController_kernelRootController_concrete1_io_in_x557_valid),
    .io_in_x557_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x557_bits_wdata_0),
    .io_in_x557_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x557_bits_wstrb),
    .io_in_x556_ready(RootController_kernelRootController_concrete1_io_in_x556_ready),
    .io_in_x556_valid(RootController_kernelRootController_concrete1_io_in_x556_valid),
    .io_in_x556_bits_addr(RootController_kernelRootController_concrete1_io_in_x556_bits_addr),
    .io_in_x556_bits_size(RootController_kernelRootController_concrete1_io_in_x556_bits_size),
    .io_in_x290_TVALID(RootController_kernelRootController_concrete1_io_in_x290_TVALID),
    .io_in_x290_TREADY(RootController_kernelRootController_concrete1_io_in_x290_TREADY),
    .io_in_x290_TDATA(RootController_kernelRootController_concrete1_io_in_x290_TDATA),
    .io_in_x287_outdram_number(RootController_kernelRootController_concrete1_io_in_x287_outdram_number),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@51818.4 package.scala 96:25:@51819.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@51889.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@51890.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@51910.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@51909.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x556_valid; // @[sm_RootController.scala 63:23:@52034.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x556_bits_addr; // @[sm_RootController.scala 63:23:@52033.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x556_bits_size; // @[sm_RootController.scala 63:23:@52032.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x557_valid; // @[sm_RootController.scala 62:23:@52030.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x557_bits_wdata_0; // @[sm_RootController.scala 62:23:@52029.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x557_bits_wstrb; // @[sm_RootController.scala 62:23:@52028.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x558_ready; // @[sm_RootController.scala 61:23:@52027.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x289_TREADY; // @[sm_RootController.scala 60:23:@52023.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x290_TVALID; // @[sm_RootController.scala 64:23:@52044.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x290_TDATA; // @[sm_RootController.scala 64:23:@52042.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 64:23:@52041.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 64:23:@52040.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 64:23:@52039.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 64:23:@52038.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 64:23:@52037.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 64:23:@52036.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@51796.4]
  assign SingleCounter_reset = reset; // @[:@51797.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@51811.4]
  assign RetimeWrapper_clock = clock; // @[:@51814.4]
  assign RetimeWrapper_reset = reset; // @[:@51815.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@51817.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@51816.4]
  assign SRFF_clock = clock; // @[:@51823.4]
  assign SRFF_reset = reset; // @[:@51824.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@52073.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@51907.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@51908.4]
  assign RootController_sm_clock = clock; // @[:@51862.4]
  assign RootController_sm_reset = reset; // @[:@51863.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@51906.4 SpatialBlocks.scala 140:18:@51940.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@51934.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@51914.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@51902.4 SpatialBlocks.scala 142:21:@51942.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@51931.4]
  assign RetimeWrapper_1_clock = clock; // @[:@51894.4]
  assign RetimeWrapper_1_reset = reset; // @[:@51895.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@51897.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@51896.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@51956.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@51957.4]
  assign RootController_kernelRootController_concrete1_io_in_x289_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 60:23:@52024.4]
  assign RootController_kernelRootController_concrete1_io_in_x289_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 60:23:@52022.4]
  assign RootController_kernelRootController_concrete1_io_in_x289_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 60:23:@52018.4]
  assign RootController_kernelRootController_concrete1_io_in_x289_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 60:23:@52017.4]
  assign RootController_kernelRootController_concrete1_io_in_x558_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 61:23:@52026.4]
  assign RootController_kernelRootController_concrete1_io_in_x557_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 62:23:@52031.4]
  assign RootController_kernelRootController_concrete1_io_in_x556_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 63:23:@52035.4]
  assign RootController_kernelRootController_concrete1_io_in_x290_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 64:23:@52043.4]
  assign RootController_kernelRootController_concrete1_io_in_x287_outdram_number = io_argIns_1; // @[sm_RootController.scala 65:31:@52045.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@52054.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@52052.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@52046.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module Counter( // @[:@52075.2]
  input        clock, // @[:@52076.4]
  input        reset, // @[:@52077.4]
  input        io_enable, // @[:@52078.4]
  output [5:0] io_out, // @[:@52078.4]
  output [5:0] io_next // @[:@52078.4]
);
  reg [5:0] count; // @[Counter.scala 15:22:@52080.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_17; // @[Counter.scala 17:24:@52081.4]
  wire [5:0] newCount; // @[Counter.scala 17:24:@52082.4]
  wire [5:0] _GEN_0; // @[Counter.scala 21:26:@52087.6]
  assign _T_17 = count + 6'h1; // @[Counter.scala 17:24:@52081.4]
  assign newCount = count + 6'h1; // @[Counter.scala 17:24:@52082.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@52087.6]
  assign io_out = count; // @[Counter.scala 25:10:@52090.4]
  assign io_next = count + 6'h1; // @[Counter.scala 26:11:@52091.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module SRAM_25( // @[:@52127.2]
  input         clock, // @[:@52128.4]
  input         reset, // @[:@52129.4]
  input  [5:0]  io_raddr, // @[:@52130.4]
  input         io_wen, // @[:@52130.4]
  input  [5:0]  io_waddr, // @[:@52130.4]
  input  [63:0] io_wdata_addr, // @[:@52130.4]
  input  [31:0] io_wdata_size, // @[:@52130.4]
  output [63:0] io_rdata_addr, // @[:@52130.4]
  output [31:0] io_rdata_size // @[:@52130.4]
);
  wire [95:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@52132.4]
  wire [95:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@52132.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@52132.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@52132.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@52132.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@52132.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@52132.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@52132.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@52132.4]
  wire [95:0] _T_17; // @[SRAM.scala 175:38:@52146.4]
  wire  _T_20; // @[SRAM.scala 182:49:@52151.4]
  wire  _T_21; // @[SRAM.scala 182:37:@52152.4]
  reg  _T_24; // @[SRAM.scala 182:29:@52153.4]
  reg [31:0] _RAND_0;
  reg [95:0] _T_28; // @[SRAM.scala 183:29:@52156.4]
  reg [95:0] _RAND_1;
  wire [95:0] _T_29; // @[SRAM.scala 184:22:@52158.4]
  SRAMVerilogAWS #(.DWIDTH(96), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@52132.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_17 = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:38:@52146.4]
  assign _T_20 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@52151.4]
  assign _T_21 = io_wen & _T_20; // @[SRAM.scala 182:37:@52152.4]
  assign _T_29 = _T_24 ? _T_28 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:22:@52158.4]
  assign io_rdata_addr = _T_29[95:32]; // @[SRAM.scala 184:16:@52167.4]
  assign io_rdata_size = _T_29[31:0]; // @[SRAM.scala 184:16:@52166.4]
  assign SRAMVerilogAWS_wdata = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:20:@52147.4]
  assign SRAMVerilogAWS_backpressure = 1'h1; // @[SRAM.scala 176:27:@52148.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@52144.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@52150.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@52149.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@52145.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@52143.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@52142.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_24 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _T_28 = _RAND_1[95:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_21;
    end
    if (reset) begin
      _T_28 <= 96'h0;
    end else begin
      _T_28 <= _T_17;
    end
  end
endmodule
module FIFO( // @[:@52169.2]
  input         clock, // @[:@52170.4]
  input         reset, // @[:@52171.4]
  output        io_in_ready, // @[:@52172.4]
  input         io_in_valid, // @[:@52172.4]
  input  [63:0] io_in_bits_addr, // @[:@52172.4]
  input  [31:0] io_in_bits_size, // @[:@52172.4]
  input         io_out_ready, // @[:@52172.4]
  output        io_out_valid, // @[:@52172.4]
  output [63:0] io_out_bits_addr, // @[:@52172.4]
  output [31:0] io_out_bits_size // @[:@52172.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@52568.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@52568.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@52568.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@52568.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@52568.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@52578.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@52578.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@52578.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@52578.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@52578.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@52593.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@52593.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@52593.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@52593.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@52593.4]
  wire [63:0] SRAM_io_wdata_addr; // @[FIFO.scala 73:19:@52593.4]
  wire [31:0] SRAM_io_wdata_size; // @[FIFO.scala 73:19:@52593.4]
  wire [63:0] SRAM_io_rdata_addr; // @[FIFO.scala 73:19:@52593.4]
  wire [31:0] SRAM_io_rdata_size; // @[FIFO.scala 73:19:@52593.4]
  wire  writeEn; // @[FIFO.scala 30:29:@52566.4]
  wire  readEn; // @[FIFO.scala 31:29:@52567.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@52588.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@52589.4]
  wire  _T_824; // @[FIFO.scala 45:27:@52590.4]
  wire  empty; // @[FIFO.scala 45:24:@52591.4]
  wire  full; // @[FIFO.scala 46:23:@52592.4]
  wire  _T_827; // @[FIFO.scala 83:17:@52605.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@52606.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@52568.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@52578.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_25 SRAM ( // @[FIFO.scala 73:19:@52593.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata_addr(SRAM_io_wdata_addr),
    .io_wdata_size(SRAM_io_wdata_size),
    .io_rdata_addr(SRAM_io_rdata_addr),
    .io_rdata_size(SRAM_io_rdata_size)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@52566.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@52567.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@52589.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@52590.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@52591.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@52592.4]
  assign _T_827 = writeEn != readEn; // @[FIFO.scala 83:17:@52605.4]
  assign _GEN_0 = _T_827 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@52606.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@52612.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@52610.4]
  assign io_out_bits_addr = SRAM_io_rdata_addr; // @[FIFO.scala 79:17:@52603.4]
  assign io_out_bits_size = SRAM_io_rdata_size; // @[FIFO.scala 79:17:@52602.4]
  assign enqCounter_clock = clock; // @[:@52569.4]
  assign enqCounter_reset = reset; // @[:@52570.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@52576.4]
  assign deqCounter_clock = clock; // @[:@52579.4]
  assign deqCounter_reset = reset; // @[:@52580.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@52586.4]
  assign SRAM_clock = clock; // @[:@52594.4]
  assign SRAM_reset = reset; // @[:@52595.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@52597.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@52598.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@52599.4]
  assign SRAM_io_wdata_addr = io_in_bits_addr; // @[FIFO.scala 78:16:@52601.4]
  assign SRAM_io_wdata_size = io_in_bits_size; // @[FIFO.scala 78:16:@52600.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_827) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module Counter_2( // @[:@52614.2]
  input        clock, // @[:@52615.4]
  input        reset, // @[:@52616.4]
  input        io_enable, // @[:@52617.4]
  output [3:0] io_out // @[:@52617.4]
);
  reg [3:0] count; // @[Counter.scala 15:22:@52619.4]
  reg [31:0] _RAND_0;
  wire [4:0] _T_17; // @[Counter.scala 17:24:@52620.4]
  wire [3:0] newCount; // @[Counter.scala 17:24:@52621.4]
  wire [3:0] _GEN_0; // @[Counter.scala 21:26:@52626.6]
  assign _T_17 = count + 4'h1; // @[Counter.scala 17:24:@52620.4]
  assign newCount = count + 4'h1; // @[Counter.scala 17:24:@52621.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@52626.6]
  assign io_out = count; // @[Counter.scala 25:10:@52629.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module Counter_4( // @[:@52650.2]
  input        clock, // @[:@52651.4]
  input        reset, // @[:@52652.4]
  input        io_reset, // @[:@52653.4]
  input        io_enable, // @[:@52653.4]
  input  [1:0] io_stride, // @[:@52653.4]
  output [1:0] io_out, // @[:@52653.4]
  output [1:0] io_next // @[:@52653.4]
);
  reg [1:0] count; // @[Counter.scala 15:22:@52655.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_17; // @[Counter.scala 17:24:@52656.4]
  wire [1:0] newCount; // @[Counter.scala 17:24:@52657.4]
  wire [1:0] _GEN_0; // @[Counter.scala 21:26:@52662.6]
  wire [1:0] _GEN_1; // @[Counter.scala 19:18:@52658.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@52656.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@52657.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@52662.6]
  assign _GEN_1 = io_reset ? 2'h0 : _GEN_0; // @[Counter.scala 19:18:@52658.4]
  assign io_out = count; // @[Counter.scala 25:10:@52665.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@52666.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 2'h0;
    end else begin
      if (io_reset) begin
        count <= 2'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_26( // @[:@52702.2]
  input         clock, // @[:@52703.4]
  input         reset, // @[:@52704.4]
  input  [1:0]  io_raddr, // @[:@52705.4]
  input         io_wen, // @[:@52705.4]
  input  [1:0]  io_waddr, // @[:@52705.4]
  input  [31:0] io_wdata, // @[:@52705.4]
  output [31:0] io_rdata, // @[:@52705.4]
  input         io_backpressure // @[:@52705.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@52707.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@52707.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@52707.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@52707.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@52707.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@52707.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@52707.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@52707.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@52707.4]
  wire  _T_19; // @[SRAM.scala 182:49:@52725.4]
  wire  _T_20; // @[SRAM.scala 182:37:@52726.4]
  reg  _T_23; // @[SRAM.scala 182:29:@52727.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@52729.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(4), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@52707.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@52725.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@52726.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@52734.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@52721.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@52722.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@52719.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@52724.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@52723.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@52720.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@52718.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@52717.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module FIFO_1( // @[:@52736.2]
  input         clock, // @[:@52737.4]
  input         reset, // @[:@52738.4]
  output        io_in_ready, // @[:@52739.4]
  input         io_in_valid, // @[:@52739.4]
  input  [31:0] io_in_bits, // @[:@52739.4]
  input         io_out_ready, // @[:@52739.4]
  output        io_out_valid, // @[:@52739.4]
  output [31:0] io_out_bits // @[:@52739.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@52765.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@52765.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@52765.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@52765.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@52765.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@52765.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@52765.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@52775.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@52775.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@52775.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@52775.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@52775.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@52775.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@52775.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@52790.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@52790.4]
  wire [1:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@52790.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@52790.4]
  wire [1:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@52790.4]
  wire [31:0] SRAM_io_wdata; // @[FIFO.scala 73:19:@52790.4]
  wire [31:0] SRAM_io_rdata; // @[FIFO.scala 73:19:@52790.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@52790.4]
  wire  writeEn; // @[FIFO.scala 30:29:@52763.4]
  wire  readEn; // @[FIFO.scala 31:29:@52764.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@52785.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@52786.4]
  wire  _T_104; // @[FIFO.scala 45:27:@52787.4]
  wire  empty; // @[FIFO.scala 45:24:@52788.4]
  wire  full; // @[FIFO.scala 46:23:@52789.4]
  wire  _T_107; // @[FIFO.scala 83:17:@52800.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@52801.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@52765.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@52775.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_26 SRAM ( // @[FIFO.scala 73:19:@52790.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@52763.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@52764.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@52786.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@52787.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@52788.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@52789.4]
  assign _T_107 = writeEn != readEn; // @[FIFO.scala 83:17:@52800.4]
  assign _GEN_0 = _T_107 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@52801.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@52807.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@52805.4]
  assign io_out_bits = SRAM_io_rdata; // @[FIFO.scala 79:17:@52798.4]
  assign enqCounter_clock = clock; // @[:@52766.4]
  assign enqCounter_reset = reset; // @[:@52767.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@52773.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@52774.4]
  assign deqCounter_clock = clock; // @[:@52776.4]
  assign deqCounter_reset = reset; // @[:@52777.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@52783.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@52784.4]
  assign SRAM_clock = clock; // @[:@52791.4]
  assign SRAM_reset = reset; // @[:@52792.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@52794.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@52795.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@52796.4]
  assign SRAM_io_wdata = io_in_bits; // @[FIFO.scala 78:16:@52797.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@52799.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_107) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec( // @[:@55194.2]
  input         clock, // @[:@55195.4]
  input         reset, // @[:@55196.4]
  output        io_in_ready, // @[:@55197.4]
  input         io_in_valid, // @[:@55197.4]
  input  [31:0] io_in_bits_0, // @[:@55197.4]
  input         io_out_ready, // @[:@55197.4]
  output        io_out_valid, // @[:@55197.4]
  output [31:0] io_out_bits_0, // @[:@55197.4]
  output [31:0] io_out_bits_1, // @[:@55197.4]
  output [31:0] io_out_bits_2, // @[:@55197.4]
  output [31:0] io_out_bits_3, // @[:@55197.4]
  output [31:0] io_out_bits_4, // @[:@55197.4]
  output [31:0] io_out_bits_5, // @[:@55197.4]
  output [31:0] io_out_bits_6, // @[:@55197.4]
  output [31:0] io_out_bits_7, // @[:@55197.4]
  output [31:0] io_out_bits_8, // @[:@55197.4]
  output [31:0] io_out_bits_9, // @[:@55197.4]
  output [31:0] io_out_bits_10, // @[:@55197.4]
  output [31:0] io_out_bits_11, // @[:@55197.4]
  output [31:0] io_out_bits_12, // @[:@55197.4]
  output [31:0] io_out_bits_13, // @[:@55197.4]
  output [31:0] io_out_bits_14, // @[:@55197.4]
  output [31:0] io_out_bits_15 // @[:@55197.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@55201.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@55201.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@55201.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@55201.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@55212.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@55212.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@55212.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@55212.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@55225.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@55225.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@55225.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@55225.4]
  wire [31:0] fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@55225.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@55225.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@55225.4]
  wire [31:0] fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@55225.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@55260.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@55260.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@55260.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@55260.4]
  wire [31:0] fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@55260.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@55260.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@55260.4]
  wire [31:0] fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@55260.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@55295.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@55295.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@55295.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@55295.4]
  wire [31:0] fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@55295.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@55295.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@55295.4]
  wire [31:0] fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@55295.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@55330.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@55330.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@55330.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@55330.4]
  wire [31:0] fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@55330.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@55330.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@55330.4]
  wire [31:0] fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@55330.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@55365.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@55365.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@55365.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@55365.4]
  wire [31:0] fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@55365.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@55365.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@55365.4]
  wire [31:0] fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@55365.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@55400.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@55400.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@55400.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@55400.4]
  wire [31:0] fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@55400.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@55400.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@55400.4]
  wire [31:0] fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@55400.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@55435.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@55435.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@55435.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@55435.4]
  wire [31:0] fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@55435.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@55435.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@55435.4]
  wire [31:0] fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@55435.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@55470.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@55470.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@55470.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@55470.4]
  wire [31:0] fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@55470.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@55470.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@55470.4]
  wire [31:0] fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@55470.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@55505.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@55505.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@55505.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@55505.4]
  wire [31:0] fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@55505.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@55505.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@55505.4]
  wire [31:0] fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@55505.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@55540.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@55540.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@55540.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@55540.4]
  wire [31:0] fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@55540.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@55540.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@55540.4]
  wire [31:0] fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@55540.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@55575.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@55575.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@55575.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@55575.4]
  wire [31:0] fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@55575.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@55575.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@55575.4]
  wire [31:0] fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@55575.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@55610.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@55610.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@55610.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@55610.4]
  wire [31:0] fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@55610.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@55610.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@55610.4]
  wire [31:0] fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@55610.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@55645.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@55645.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@55645.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@55645.4]
  wire [31:0] fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@55645.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@55645.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@55645.4]
  wire [31:0] fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@55645.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@55680.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@55680.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@55680.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@55680.4]
  wire [31:0] fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@55680.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@55680.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@55680.4]
  wire [31:0] fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@55680.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@55715.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@55715.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@55715.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@55715.4]
  wire [31:0] fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@55715.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@55715.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@55715.4]
  wire [31:0] fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@55715.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@55750.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@55750.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@55750.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@55750.4]
  wire [31:0] fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@55750.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@55750.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@55750.4]
  wire [31:0] fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@55750.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@55200.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@55223.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@55250.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@55285.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@55320.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@55355.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@55390.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@55425.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@55460.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@55495.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@55530.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@55565.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@55600.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@55635.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@55670.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@55705.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@55740.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@55775.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55786.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55787.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@55817.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55788.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@55817.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55789.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@55817.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55790.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@55817.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55791.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@55817.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55792.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@55817.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55793.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@55817.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55794.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@55817.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55795.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@55817.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55796.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@55817.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55797.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@55817.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55798.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@55817.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55799.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@55817.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55800.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@55817.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55801.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@55836.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@55837.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@55838.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@55839.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@55840.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@55841.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@55842.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@55843.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@55844.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@55845.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@55846.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@55847.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@55848.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@55849.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@55201.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@55212.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_1 fifos_0 ( // @[FIFOVec.scala 40:19:@55225.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_1 fifos_1 ( // @[FIFOVec.scala 40:19:@55260.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_1 fifos_2 ( // @[FIFOVec.scala 40:19:@55295.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_1 fifos_3 ( // @[FIFOVec.scala 40:19:@55330.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_1 fifos_4 ( // @[FIFOVec.scala 40:19:@55365.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_1 fifos_5 ( // @[FIFOVec.scala 40:19:@55400.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_1 fifos_6 ( // @[FIFOVec.scala 40:19:@55435.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_1 fifos_7 ( // @[FIFOVec.scala 40:19:@55470.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_1 fifos_8 ( // @[FIFOVec.scala 40:19:@55505.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_1 fifos_9 ( // @[FIFOVec.scala 40:19:@55540.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_1 fifos_10 ( // @[FIFOVec.scala 40:19:@55575.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_1 fifos_11 ( // @[FIFOVec.scala 40:19:@55610.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_1 fifos_12 ( // @[FIFOVec.scala 40:19:@55645.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_1 fifos_13 ( // @[FIFOVec.scala 40:19:@55680.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_1 fifos_14 ( // @[FIFOVec.scala 40:19:@55715.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_1 fifos_15 ( // @[FIFOVec.scala 40:19:@55750.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@55200.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@55223.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@55250.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@55285.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@55320.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@55355.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@55390.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@55425.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@55460.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@55495.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@55530.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@55565.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@55600.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@55635.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@55670.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@55705.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@55740.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@55775.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55786.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55787.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@55817.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55788.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@55817.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55789.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@55817.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55790.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@55817.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55791.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@55817.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55792.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@55817.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55793.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@55817.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55794.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@55817.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55795.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@55817.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55796.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@55817.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55797.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@55817.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55798.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@55817.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55799.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@55817.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55800.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@55817.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@55785.4 FIFOVec.scala 49:42:@55801.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@55836.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@55837.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@55838.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@55839.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@55840.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@55841.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@55842.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@55843.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@55844.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@55845.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@55846.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@55847.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@55848.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@55849.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@55818.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@55852.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@56160.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@56161.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@56162.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@56163.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@56164.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@56165.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@56166.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@56167.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@56168.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@56169.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@56170.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@56171.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@56172.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@56173.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@56174.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@56175.4]
  assign enqCounter_clock = clock; // @[:@55202.4]
  assign enqCounter_reset = reset; // @[:@55203.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@55210.4]
  assign deqCounter_clock = clock; // @[:@55213.4]
  assign deqCounter_reset = reset; // @[:@55214.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@55221.4]
  assign fifos_0_clock = clock; // @[:@55226.4]
  assign fifos_0_reset = reset; // @[:@55227.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@55253.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55255.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55259.4]
  assign fifos_1_clock = clock; // @[:@55261.4]
  assign fifos_1_reset = reset; // @[:@55262.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@55288.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55290.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55294.4]
  assign fifos_2_clock = clock; // @[:@55296.4]
  assign fifos_2_reset = reset; // @[:@55297.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@55323.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55325.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55329.4]
  assign fifos_3_clock = clock; // @[:@55331.4]
  assign fifos_3_reset = reset; // @[:@55332.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@55358.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55360.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55364.4]
  assign fifos_4_clock = clock; // @[:@55366.4]
  assign fifos_4_reset = reset; // @[:@55367.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@55393.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55395.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55399.4]
  assign fifos_5_clock = clock; // @[:@55401.4]
  assign fifos_5_reset = reset; // @[:@55402.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@55428.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55430.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55434.4]
  assign fifos_6_clock = clock; // @[:@55436.4]
  assign fifos_6_reset = reset; // @[:@55437.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@55463.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55465.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55469.4]
  assign fifos_7_clock = clock; // @[:@55471.4]
  assign fifos_7_reset = reset; // @[:@55472.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@55498.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55500.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55504.4]
  assign fifos_8_clock = clock; // @[:@55506.4]
  assign fifos_8_reset = reset; // @[:@55507.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@55533.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55535.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55539.4]
  assign fifos_9_clock = clock; // @[:@55541.4]
  assign fifos_9_reset = reset; // @[:@55542.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@55568.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55570.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55574.4]
  assign fifos_10_clock = clock; // @[:@55576.4]
  assign fifos_10_reset = reset; // @[:@55577.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@55603.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55605.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55609.4]
  assign fifos_11_clock = clock; // @[:@55611.4]
  assign fifos_11_reset = reset; // @[:@55612.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@55638.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55640.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55644.4]
  assign fifos_12_clock = clock; // @[:@55646.4]
  assign fifos_12_reset = reset; // @[:@55647.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@55673.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55675.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55679.4]
  assign fifos_13_clock = clock; // @[:@55681.4]
  assign fifos_13_reset = reset; // @[:@55682.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@55708.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55710.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55714.4]
  assign fifos_14_clock = clock; // @[:@55716.4]
  assign fifos_14_reset = reset; // @[:@55717.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@55743.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55745.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55749.4]
  assign fifos_15_clock = clock; // @[:@55751.4]
  assign fifos_15_reset = reset; // @[:@55752.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@55778.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@55780.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@55784.4]
endmodule
module FFRAM( // @[:@56249.2]
  input        clock, // @[:@56250.4]
  input        reset, // @[:@56251.4]
  input  [1:0] io_raddr, // @[:@56252.4]
  input        io_wen, // @[:@56252.4]
  input  [1:0] io_waddr, // @[:@56252.4]
  input        io_wdata, // @[:@56252.4]
  output       io_rdata, // @[:@56252.4]
  input        io_banks_0_wdata_valid, // @[:@56252.4]
  input        io_banks_0_wdata_bits, // @[:@56252.4]
  input        io_banks_1_wdata_valid, // @[:@56252.4]
  input        io_banks_1_wdata_bits, // @[:@56252.4]
  input        io_banks_2_wdata_valid, // @[:@56252.4]
  input        io_banks_2_wdata_bits, // @[:@56252.4]
  input        io_banks_3_wdata_valid, // @[:@56252.4]
  input        io_banks_3_wdata_bits // @[:@56252.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@56256.4]
  reg [31:0] _RAND_0;
  wire  _T_88; // @[SRAM.scala 148:37:@56257.4]
  wire  _T_89; // @[SRAM.scala 148:25:@56258.4]
  wire  _T_90; // @[SRAM.scala 148:15:@56259.4]
  wire  _T_91; // @[SRAM.scala 149:15:@56261.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@56260.4]
  reg  regs_1; // @[SRAM.scala 145:20:@56267.4]
  reg [31:0] _RAND_1;
  wire  _T_97; // @[SRAM.scala 148:37:@56268.4]
  wire  _T_98; // @[SRAM.scala 148:25:@56269.4]
  wire  _T_99; // @[SRAM.scala 148:15:@56270.4]
  wire  _T_100; // @[SRAM.scala 149:15:@56272.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@56271.4]
  reg  regs_2; // @[SRAM.scala 145:20:@56278.4]
  reg [31:0] _RAND_2;
  wire  _T_106; // @[SRAM.scala 148:37:@56279.4]
  wire  _T_107; // @[SRAM.scala 148:25:@56280.4]
  wire  _T_108; // @[SRAM.scala 148:15:@56281.4]
  wire  _T_109; // @[SRAM.scala 149:15:@56283.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@56282.4]
  reg  regs_3; // @[SRAM.scala 145:20:@56289.4]
  reg [31:0] _RAND_3;
  wire  _T_115; // @[SRAM.scala 148:37:@56290.4]
  wire  _T_116; // @[SRAM.scala 148:25:@56291.4]
  wire  _T_117; // @[SRAM.scala 148:15:@56292.4]
  wire  _T_118; // @[SRAM.scala 149:15:@56294.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@56293.4]
  wire  _GEN_5; // @[SRAM.scala 155:12:@56303.4]
  wire  _GEN_6; // @[SRAM.scala 155:12:@56303.4]
  assign _T_88 = io_waddr == 2'h0; // @[SRAM.scala 148:37:@56257.4]
  assign _T_89 = io_wen & _T_88; // @[SRAM.scala 148:25:@56258.4]
  assign _T_90 = io_banks_0_wdata_valid | _T_89; // @[SRAM.scala 148:15:@56259.4]
  assign _T_91 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@56261.6]
  assign _GEN_0 = _T_90 ? _T_91 : regs_0; // @[SRAM.scala 148:48:@56260.4]
  assign _T_97 = io_waddr == 2'h1; // @[SRAM.scala 148:37:@56268.4]
  assign _T_98 = io_wen & _T_97; // @[SRAM.scala 148:25:@56269.4]
  assign _T_99 = io_banks_1_wdata_valid | _T_98; // @[SRAM.scala 148:15:@56270.4]
  assign _T_100 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@56272.6]
  assign _GEN_1 = _T_99 ? _T_100 : regs_1; // @[SRAM.scala 148:48:@56271.4]
  assign _T_106 = io_waddr == 2'h2; // @[SRAM.scala 148:37:@56279.4]
  assign _T_107 = io_wen & _T_106; // @[SRAM.scala 148:25:@56280.4]
  assign _T_108 = io_banks_2_wdata_valid | _T_107; // @[SRAM.scala 148:15:@56281.4]
  assign _T_109 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@56283.6]
  assign _GEN_2 = _T_108 ? _T_109 : regs_2; // @[SRAM.scala 148:48:@56282.4]
  assign _T_115 = io_waddr == 2'h3; // @[SRAM.scala 148:37:@56290.4]
  assign _T_116 = io_wen & _T_115; // @[SRAM.scala 148:25:@56291.4]
  assign _T_117 = io_banks_3_wdata_valid | _T_116; // @[SRAM.scala 148:15:@56292.4]
  assign _T_118 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@56294.6]
  assign _GEN_3 = _T_117 ? _T_118 : regs_3; // @[SRAM.scala 148:48:@56293.4]
  assign _GEN_5 = 2'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@56303.4]
  assign _GEN_6 = 2'h2 == io_raddr ? regs_2 : _GEN_5; // @[SRAM.scala 155:12:@56303.4]
  assign io_rdata = 2'h3 == io_raddr ? regs_3 : _GEN_6; // @[SRAM.scala 155:12:@56303.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_90) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_99) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_108) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_117) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_17( // @[:@56305.2]
  input   clock, // @[:@56306.4]
  input   reset, // @[:@56307.4]
  output  io_in_ready, // @[:@56308.4]
  input   io_in_valid, // @[:@56308.4]
  input   io_in_bits, // @[:@56308.4]
  input   io_out_ready, // @[:@56308.4]
  output  io_out_valid, // @[:@56308.4]
  output  io_out_bits // @[:@56308.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@56334.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@56334.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@56334.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@56334.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@56334.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@56334.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@56334.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@56344.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@56344.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@56344.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@56344.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@56344.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@56344.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@56344.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@56359.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@56359.4]
  wire [1:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@56359.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@56359.4]
  wire [1:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@56359.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@56359.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@56359.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@56359.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@56359.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@56359.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@56359.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@56359.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@56359.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@56359.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@56359.4]
  wire  writeEn; // @[FIFO.scala 30:29:@56332.4]
  wire  readEn; // @[FIFO.scala 31:29:@56333.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@56354.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@56355.4]
  wire  _T_104; // @[FIFO.scala 45:27:@56356.4]
  wire  empty; // @[FIFO.scala 45:24:@56357.4]
  wire  full; // @[FIFO.scala 46:23:@56358.4]
  wire  _T_157; // @[FIFO.scala 83:17:@56445.4]
  wire  _GEN_4; // @[FIFO.scala 83:29:@56446.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@56334.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@56344.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM FFRAM ( // @[FIFO.scala 49:19:@56359.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@56332.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@56333.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@56355.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@56356.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@56357.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@56358.4]
  assign _T_157 = writeEn != readEn; // @[FIFO.scala 83:17:@56445.4]
  assign _GEN_4 = _T_157 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@56446.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@56452.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@56450.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@56384.4]
  assign enqCounter_clock = clock; // @[:@56335.4]
  assign enqCounter_reset = reset; // @[:@56336.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@56342.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@56343.4]
  assign deqCounter_clock = clock; // @[:@56345.4]
  assign deqCounter_reset = reset; // @[:@56346.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@56352.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@56353.4]
  assign FFRAM_clock = clock; // @[:@56360.4]
  assign FFRAM_reset = reset; // @[:@56361.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@56380.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@56381.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@56382.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@56383.4]
  assign FFRAM_io_banks_0_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@56386.4]
  assign FFRAM_io_banks_0_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@56385.4]
  assign FFRAM_io_banks_1_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@56389.4]
  assign FFRAM_io_banks_1_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@56388.4]
  assign FFRAM_io_banks_2_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@56392.4]
  assign FFRAM_io_banks_2_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@56391.4]
  assign FFRAM_io_banks_3_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@56395.4]
  assign FFRAM_io_banks_3_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@56394.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_157) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_1( // @[:@60069.2]
  input   clock, // @[:@60070.4]
  input   reset, // @[:@60071.4]
  output  io_in_ready, // @[:@60072.4]
  input   io_in_valid, // @[:@60072.4]
  input   io_in_bits_0, // @[:@60072.4]
  input   io_out_ready, // @[:@60072.4]
  output  io_out_valid, // @[:@60072.4]
  output  io_out_bits_0, // @[:@60072.4]
  output  io_out_bits_1, // @[:@60072.4]
  output  io_out_bits_2, // @[:@60072.4]
  output  io_out_bits_3, // @[:@60072.4]
  output  io_out_bits_4, // @[:@60072.4]
  output  io_out_bits_5, // @[:@60072.4]
  output  io_out_bits_6, // @[:@60072.4]
  output  io_out_bits_7, // @[:@60072.4]
  output  io_out_bits_8, // @[:@60072.4]
  output  io_out_bits_9, // @[:@60072.4]
  output  io_out_bits_10, // @[:@60072.4]
  output  io_out_bits_11, // @[:@60072.4]
  output  io_out_bits_12, // @[:@60072.4]
  output  io_out_bits_13, // @[:@60072.4]
  output  io_out_bits_14, // @[:@60072.4]
  output  io_out_bits_15 // @[:@60072.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@60076.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@60076.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@60076.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@60076.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@60087.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@60087.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@60087.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@60087.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@60100.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@60100.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@60100.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@60100.4]
  wire  fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@60100.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@60100.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@60100.4]
  wire  fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@60100.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@60135.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@60135.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@60135.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@60135.4]
  wire  fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@60135.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@60135.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@60135.4]
  wire  fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@60135.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@60170.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@60170.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@60170.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@60170.4]
  wire  fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@60170.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@60170.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@60170.4]
  wire  fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@60170.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@60205.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@60205.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@60205.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@60205.4]
  wire  fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@60205.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@60205.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@60205.4]
  wire  fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@60205.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@60240.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@60240.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@60240.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@60240.4]
  wire  fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@60240.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@60240.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@60240.4]
  wire  fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@60240.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@60275.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@60275.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@60275.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@60275.4]
  wire  fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@60275.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@60275.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@60275.4]
  wire  fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@60275.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@60310.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@60310.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@60310.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@60310.4]
  wire  fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@60310.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@60310.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@60310.4]
  wire  fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@60310.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@60345.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@60345.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@60345.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@60345.4]
  wire  fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@60345.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@60345.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@60345.4]
  wire  fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@60345.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@60380.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@60380.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@60380.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@60380.4]
  wire  fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@60380.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@60380.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@60380.4]
  wire  fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@60380.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@60415.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@60415.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@60415.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@60415.4]
  wire  fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@60415.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@60415.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@60415.4]
  wire  fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@60415.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@60450.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@60450.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@60450.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@60450.4]
  wire  fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@60450.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@60450.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@60450.4]
  wire  fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@60450.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@60485.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@60485.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@60485.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@60485.4]
  wire  fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@60485.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@60485.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@60485.4]
  wire  fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@60485.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@60520.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@60520.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@60520.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@60520.4]
  wire  fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@60520.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@60520.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@60520.4]
  wire  fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@60520.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@60555.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@60555.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@60555.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@60555.4]
  wire  fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@60555.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@60555.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@60555.4]
  wire  fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@60555.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@60590.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@60590.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@60590.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@60590.4]
  wire  fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@60590.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@60590.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@60590.4]
  wire  fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@60590.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@60625.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@60625.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@60625.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@60625.4]
  wire  fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@60625.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@60625.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@60625.4]
  wire  fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@60625.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@60075.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@60098.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@60125.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@60160.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@60195.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@60230.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@60265.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@60300.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@60335.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@60370.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@60405.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@60440.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@60475.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@60510.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@60545.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@60580.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@60615.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@60650.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60661.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60662.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@60692.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60663.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@60692.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60664.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@60692.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60665.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@60692.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60666.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@60692.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60667.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@60692.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60668.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@60692.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60669.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@60692.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60670.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@60692.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60671.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@60692.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60672.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@60692.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60673.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@60692.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60674.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@60692.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60675.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@60692.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60676.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@60711.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@60712.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@60713.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@60714.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@60715.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@60716.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@60717.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@60718.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@60719.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@60720.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@60721.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@60722.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@60723.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@60724.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@60076.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@60087.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_17 fifos_0 ( // @[FIFOVec.scala 40:19:@60100.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_17 fifos_1 ( // @[FIFOVec.scala 40:19:@60135.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_17 fifos_2 ( // @[FIFOVec.scala 40:19:@60170.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_17 fifos_3 ( // @[FIFOVec.scala 40:19:@60205.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_17 fifos_4 ( // @[FIFOVec.scala 40:19:@60240.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_17 fifos_5 ( // @[FIFOVec.scala 40:19:@60275.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_17 fifos_6 ( // @[FIFOVec.scala 40:19:@60310.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_17 fifos_7 ( // @[FIFOVec.scala 40:19:@60345.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_17 fifos_8 ( // @[FIFOVec.scala 40:19:@60380.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_17 fifos_9 ( // @[FIFOVec.scala 40:19:@60415.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_17 fifos_10 ( // @[FIFOVec.scala 40:19:@60450.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_17 fifos_11 ( // @[FIFOVec.scala 40:19:@60485.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_17 fifos_12 ( // @[FIFOVec.scala 40:19:@60520.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_17 fifos_13 ( // @[FIFOVec.scala 40:19:@60555.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_17 fifos_14 ( // @[FIFOVec.scala 40:19:@60590.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_17 fifos_15 ( // @[FIFOVec.scala 40:19:@60625.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@60075.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@60098.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@60125.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@60160.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@60195.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@60230.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@60265.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@60300.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@60335.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@60370.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@60405.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@60440.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@60475.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@60510.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@60545.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@60580.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@60615.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@60650.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60661.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60662.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@60692.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60663.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@60692.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60664.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@60692.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60665.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@60692.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60666.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@60692.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60667.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@60692.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60668.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@60692.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60669.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@60692.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60670.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@60692.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60671.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@60692.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60672.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@60692.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60673.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@60692.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60674.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@60692.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60675.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@60692.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@60660.4 FIFOVec.scala 49:42:@60676.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@60711.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@60712.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@60713.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@60714.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@60715.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@60716.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@60717.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@60718.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@60719.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@60720.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@60721.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@60722.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@60723.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@60724.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@60693.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@60727.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@61035.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@61036.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@61037.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@61038.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@61039.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@61040.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@61041.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@61042.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@61043.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@61044.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@61045.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@61046.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@61047.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@61048.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@61049.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@61050.4]
  assign enqCounter_clock = clock; // @[:@60077.4]
  assign enqCounter_reset = reset; // @[:@60078.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@60085.4]
  assign deqCounter_clock = clock; // @[:@60088.4]
  assign deqCounter_reset = reset; // @[:@60089.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@60096.4]
  assign fifos_0_clock = clock; // @[:@60101.4]
  assign fifos_0_reset = reset; // @[:@60102.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@60128.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60130.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60134.4]
  assign fifos_1_clock = clock; // @[:@60136.4]
  assign fifos_1_reset = reset; // @[:@60137.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@60163.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60165.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60169.4]
  assign fifos_2_clock = clock; // @[:@60171.4]
  assign fifos_2_reset = reset; // @[:@60172.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@60198.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60200.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60204.4]
  assign fifos_3_clock = clock; // @[:@60206.4]
  assign fifos_3_reset = reset; // @[:@60207.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@60233.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60235.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60239.4]
  assign fifos_4_clock = clock; // @[:@60241.4]
  assign fifos_4_reset = reset; // @[:@60242.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@60268.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60270.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60274.4]
  assign fifos_5_clock = clock; // @[:@60276.4]
  assign fifos_5_reset = reset; // @[:@60277.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@60303.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60305.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60309.4]
  assign fifos_6_clock = clock; // @[:@60311.4]
  assign fifos_6_reset = reset; // @[:@60312.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@60338.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60340.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60344.4]
  assign fifos_7_clock = clock; // @[:@60346.4]
  assign fifos_7_reset = reset; // @[:@60347.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@60373.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60375.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60379.4]
  assign fifos_8_clock = clock; // @[:@60381.4]
  assign fifos_8_reset = reset; // @[:@60382.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@60408.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60410.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60414.4]
  assign fifos_9_clock = clock; // @[:@60416.4]
  assign fifos_9_reset = reset; // @[:@60417.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@60443.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60445.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60449.4]
  assign fifos_10_clock = clock; // @[:@60451.4]
  assign fifos_10_reset = reset; // @[:@60452.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@60478.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60480.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60484.4]
  assign fifos_11_clock = clock; // @[:@60486.4]
  assign fifos_11_reset = reset; // @[:@60487.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@60513.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60515.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60519.4]
  assign fifos_12_clock = clock; // @[:@60521.4]
  assign fifos_12_reset = reset; // @[:@60522.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@60548.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60550.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60554.4]
  assign fifos_13_clock = clock; // @[:@60556.4]
  assign fifos_13_reset = reset; // @[:@60557.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@60583.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60585.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60589.4]
  assign fifos_14_clock = clock; // @[:@60591.4]
  assign fifos_14_reset = reset; // @[:@60592.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@60618.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60620.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60624.4]
  assign fifos_15_clock = clock; // @[:@60626.4]
  assign fifos_15_reset = reset; // @[:@60627.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@60653.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@60655.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@60659.4]
endmodule
module FIFOWidthConvert( // @[:@61052.2]
  input         clock, // @[:@61053.4]
  input         reset, // @[:@61054.4]
  output        io_in_ready, // @[:@61055.4]
  input         io_in_valid, // @[:@61055.4]
  input  [31:0] io_in_bits_data_0, // @[:@61055.4]
  input         io_in_bits_strobe, // @[:@61055.4]
  input         io_out_ready, // @[:@61055.4]
  output        io_out_valid, // @[:@61055.4]
  output [31:0] io_out_bits_data_0, // @[:@61055.4]
  output [31:0] io_out_bits_data_1, // @[:@61055.4]
  output [31:0] io_out_bits_data_2, // @[:@61055.4]
  output [31:0] io_out_bits_data_3, // @[:@61055.4]
  output [31:0] io_out_bits_data_4, // @[:@61055.4]
  output [31:0] io_out_bits_data_5, // @[:@61055.4]
  output [31:0] io_out_bits_data_6, // @[:@61055.4]
  output [31:0] io_out_bits_data_7, // @[:@61055.4]
  output [31:0] io_out_bits_data_8, // @[:@61055.4]
  output [31:0] io_out_bits_data_9, // @[:@61055.4]
  output [31:0] io_out_bits_data_10, // @[:@61055.4]
  output [31:0] io_out_bits_data_11, // @[:@61055.4]
  output [31:0] io_out_bits_data_12, // @[:@61055.4]
  output [31:0] io_out_bits_data_13, // @[:@61055.4]
  output [31:0] io_out_bits_data_14, // @[:@61055.4]
  output [31:0] io_out_bits_data_15, // @[:@61055.4]
  output [63:0] io_out_bits_strobe // @[:@61055.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 61:22:@61057.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_in_bits_0; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_ready; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_valid; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_0; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_1; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_2; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_3; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_4; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_5; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_6; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_7; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_8; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_9; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_10; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_11; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_12; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_13; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_14; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire  FIFOVec_1_io_out_bits_15; // @[FIFOWidthConvert.scala 62:26:@61098.4]
  wire [319:0] _T_55; // @[Cat.scala 30:58:@61157.4]
  wire [511:0] _T_61; // @[Cat.scala 30:58:@61163.4]
  wire [9:0] _T_108; // @[Cat.scala 30:58:@61221.4]
  wire [15:0] _T_114; // @[Cat.scala 30:58:@61227.4]
  wire  _T_115; // @[FIFOWidthConvert.scala 36:14:@61228.4]
  wire  _T_119; // @[FIFOWidthConvert.scala 36:14:@61232.4]
  wire  _T_123; // @[FIFOWidthConvert.scala 36:14:@61236.4]
  wire  _T_127; // @[FIFOWidthConvert.scala 36:14:@61240.4]
  wire  _T_131; // @[FIFOWidthConvert.scala 36:14:@61244.4]
  wire  _T_135; // @[FIFOWidthConvert.scala 36:14:@61248.4]
  wire  _T_139; // @[FIFOWidthConvert.scala 36:14:@61252.4]
  wire  _T_143; // @[FIFOWidthConvert.scala 36:14:@61256.4]
  wire  _T_147; // @[FIFOWidthConvert.scala 36:14:@61260.4]
  wire  _T_151; // @[FIFOWidthConvert.scala 36:14:@61264.4]
  wire  _T_155; // @[FIFOWidthConvert.scala 36:14:@61268.4]
  wire  _T_159; // @[FIFOWidthConvert.scala 36:14:@61272.4]
  wire  _T_163; // @[FIFOWidthConvert.scala 36:14:@61276.4]
  wire  _T_167; // @[FIFOWidthConvert.scala 36:14:@61280.4]
  wire  _T_171; // @[FIFOWidthConvert.scala 36:14:@61284.4]
  wire  _T_175; // @[FIFOWidthConvert.scala 36:14:@61288.4]
  wire [9:0] _T_257; // @[Cat.scala 30:58:@61365.4]
  wire [18:0] _T_266; // @[Cat.scala 30:58:@61374.4]
  wire [27:0] _T_275; // @[Cat.scala 30:58:@61383.4]
  wire [36:0] _T_284; // @[Cat.scala 30:58:@61392.4]
  wire [45:0] _T_293; // @[Cat.scala 30:58:@61401.4]
  wire [54:0] _T_302; // @[Cat.scala 30:58:@61410.4]
  wire [62:0] _T_310; // @[Cat.scala 30:58:@61418.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 61:22:@61057.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15)
  );
  FIFOVec_1 FIFOVec_1 ( // @[FIFOWidthConvert.scala 62:26:@61098.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid),
    .io_in_bits_0(FIFOVec_1_io_in_bits_0),
    .io_out_ready(FIFOVec_1_io_out_ready),
    .io_out_valid(FIFOVec_1_io_out_valid),
    .io_out_bits_0(FIFOVec_1_io_out_bits_0),
    .io_out_bits_1(FIFOVec_1_io_out_bits_1),
    .io_out_bits_2(FIFOVec_1_io_out_bits_2),
    .io_out_bits_3(FIFOVec_1_io_out_bits_3),
    .io_out_bits_4(FIFOVec_1_io_out_bits_4),
    .io_out_bits_5(FIFOVec_1_io_out_bits_5),
    .io_out_bits_6(FIFOVec_1_io_out_bits_6),
    .io_out_bits_7(FIFOVec_1_io_out_bits_7),
    .io_out_bits_8(FIFOVec_1_io_out_bits_8),
    .io_out_bits_9(FIFOVec_1_io_out_bits_9),
    .io_out_bits_10(FIFOVec_1_io_out_bits_10),
    .io_out_bits_11(FIFOVec_1_io_out_bits_11),
    .io_out_bits_12(FIFOVec_1_io_out_bits_12),
    .io_out_bits_13(FIFOVec_1_io_out_bits_13),
    .io_out_bits_14(FIFOVec_1_io_out_bits_14),
    .io_out_bits_15(FIFOVec_1_io_out_bits_15)
  );
  assign _T_55 = {FIFOVec_io_out_bits_15,FIFOVec_io_out_bits_14,FIFOVec_io_out_bits_13,FIFOVec_io_out_bits_12,FIFOVec_io_out_bits_11,FIFOVec_io_out_bits_10,FIFOVec_io_out_bits_9,FIFOVec_io_out_bits_8,FIFOVec_io_out_bits_7,FIFOVec_io_out_bits_6}; // @[Cat.scala 30:58:@61157.4]
  assign _T_61 = {_T_55,FIFOVec_io_out_bits_5,FIFOVec_io_out_bits_4,FIFOVec_io_out_bits_3,FIFOVec_io_out_bits_2,FIFOVec_io_out_bits_1,FIFOVec_io_out_bits_0}; // @[Cat.scala 30:58:@61163.4]
  assign _T_108 = {FIFOVec_1_io_out_bits_0,FIFOVec_1_io_out_bits_1,FIFOVec_1_io_out_bits_2,FIFOVec_1_io_out_bits_3,FIFOVec_1_io_out_bits_4,FIFOVec_1_io_out_bits_5,FIFOVec_1_io_out_bits_6,FIFOVec_1_io_out_bits_7,FIFOVec_1_io_out_bits_8,FIFOVec_1_io_out_bits_9}; // @[Cat.scala 30:58:@61221.4]
  assign _T_114 = {_T_108,FIFOVec_1_io_out_bits_10,FIFOVec_1_io_out_bits_11,FIFOVec_1_io_out_bits_12,FIFOVec_1_io_out_bits_13,FIFOVec_1_io_out_bits_14,FIFOVec_1_io_out_bits_15}; // @[Cat.scala 30:58:@61227.4]
  assign _T_115 = _T_114[0]; // @[FIFOWidthConvert.scala 36:14:@61228.4]
  assign _T_119 = _T_114[1]; // @[FIFOWidthConvert.scala 36:14:@61232.4]
  assign _T_123 = _T_114[2]; // @[FIFOWidthConvert.scala 36:14:@61236.4]
  assign _T_127 = _T_114[3]; // @[FIFOWidthConvert.scala 36:14:@61240.4]
  assign _T_131 = _T_114[4]; // @[FIFOWidthConvert.scala 36:14:@61244.4]
  assign _T_135 = _T_114[5]; // @[FIFOWidthConvert.scala 36:14:@61248.4]
  assign _T_139 = _T_114[6]; // @[FIFOWidthConvert.scala 36:14:@61252.4]
  assign _T_143 = _T_114[7]; // @[FIFOWidthConvert.scala 36:14:@61256.4]
  assign _T_147 = _T_114[8]; // @[FIFOWidthConvert.scala 36:14:@61260.4]
  assign _T_151 = _T_114[9]; // @[FIFOWidthConvert.scala 36:14:@61264.4]
  assign _T_155 = _T_114[10]; // @[FIFOWidthConvert.scala 36:14:@61268.4]
  assign _T_159 = _T_114[11]; // @[FIFOWidthConvert.scala 36:14:@61272.4]
  assign _T_163 = _T_114[12]; // @[FIFOWidthConvert.scala 36:14:@61276.4]
  assign _T_167 = _T_114[13]; // @[FIFOWidthConvert.scala 36:14:@61280.4]
  assign _T_171 = _T_114[14]; // @[FIFOWidthConvert.scala 36:14:@61284.4]
  assign _T_175 = _T_114[15]; // @[FIFOWidthConvert.scala 36:14:@61288.4]
  assign _T_257 = {_T_175,_T_175,_T_175,_T_175,_T_171,_T_171,_T_171,_T_171,_T_167,_T_167}; // @[Cat.scala 30:58:@61365.4]
  assign _T_266 = {_T_257,_T_167,_T_167,_T_163,_T_163,_T_163,_T_163,_T_159,_T_159,_T_159}; // @[Cat.scala 30:58:@61374.4]
  assign _T_275 = {_T_266,_T_159,_T_155,_T_155,_T_155,_T_155,_T_151,_T_151,_T_151,_T_151}; // @[Cat.scala 30:58:@61383.4]
  assign _T_284 = {_T_275,_T_147,_T_147,_T_147,_T_147,_T_143,_T_143,_T_143,_T_143,_T_139}; // @[Cat.scala 30:58:@61392.4]
  assign _T_293 = {_T_284,_T_139,_T_139,_T_139,_T_135,_T_135,_T_135,_T_135,_T_131,_T_131}; // @[Cat.scala 30:58:@61401.4]
  assign _T_302 = {_T_293,_T_131,_T_131,_T_127,_T_127,_T_127,_T_127,_T_123,_T_123,_T_123}; // @[Cat.scala 30:58:@61410.4]
  assign _T_310 = {_T_302,_T_123,_T_119,_T_119,_T_119,_T_119,_T_115,_T_115,_T_115}; // @[Cat.scala 30:58:@61418.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 71:17:@61147.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 72:18:@61148.4]
  assign io_out_bits_data_0 = _T_61[31:0]; // @[FIFOWidthConvert.scala 73:22:@61197.4]
  assign io_out_bits_data_1 = _T_61[63:32]; // @[FIFOWidthConvert.scala 73:22:@61198.4]
  assign io_out_bits_data_2 = _T_61[95:64]; // @[FIFOWidthConvert.scala 73:22:@61199.4]
  assign io_out_bits_data_3 = _T_61[127:96]; // @[FIFOWidthConvert.scala 73:22:@61200.4]
  assign io_out_bits_data_4 = _T_61[159:128]; // @[FIFOWidthConvert.scala 73:22:@61201.4]
  assign io_out_bits_data_5 = _T_61[191:160]; // @[FIFOWidthConvert.scala 73:22:@61202.4]
  assign io_out_bits_data_6 = _T_61[223:192]; // @[FIFOWidthConvert.scala 73:22:@61203.4]
  assign io_out_bits_data_7 = _T_61[255:224]; // @[FIFOWidthConvert.scala 73:22:@61204.4]
  assign io_out_bits_data_8 = _T_61[287:256]; // @[FIFOWidthConvert.scala 73:22:@61205.4]
  assign io_out_bits_data_9 = _T_61[319:288]; // @[FIFOWidthConvert.scala 73:22:@61206.4]
  assign io_out_bits_data_10 = _T_61[351:320]; // @[FIFOWidthConvert.scala 73:22:@61207.4]
  assign io_out_bits_data_11 = _T_61[383:352]; // @[FIFOWidthConvert.scala 73:22:@61208.4]
  assign io_out_bits_data_12 = _T_61[415:384]; // @[FIFOWidthConvert.scala 73:22:@61209.4]
  assign io_out_bits_data_13 = _T_61[447:416]; // @[FIFOWidthConvert.scala 73:22:@61210.4]
  assign io_out_bits_data_14 = _T_61[479:448]; // @[FIFOWidthConvert.scala 73:22:@61211.4]
  assign io_out_bits_data_15 = _T_61[511:480]; // @[FIFOWidthConvert.scala 73:22:@61212.4]
  assign io_out_bits_strobe = {_T_310,_T_115}; // @[FIFOWidthConvert.scala 74:24:@61420.4]
  assign FIFOVec_clock = clock; // @[:@61058.4]
  assign FIFOVec_reset = reset; // @[:@61059.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 68:22:@61144.4]
  assign FIFOVec_io_in_bits_0 = io_in_bits_data_0; // @[FIFOWidthConvert.scala 67:24:@61143.4]
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 75:23:@61421.4]
  assign FIFOVec_1_clock = clock; // @[:@61099.4]
  assign FIFOVec_1_reset = reset; // @[:@61100.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 70:26:@61146.4]
  assign FIFOVec_1_io_in_bits_0 = io_in_bits_strobe; // @[FIFOWidthConvert.scala 69:28:@61145.4]
  assign FIFOVec_1_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 76:27:@61422.4]
endmodule
module FFRAM_16( // @[:@61460.2]
  input        clock, // @[:@61461.4]
  input        reset, // @[:@61462.4]
  input  [5:0] io_raddr, // @[:@61463.4]
  input        io_wen, // @[:@61463.4]
  input  [5:0] io_waddr, // @[:@61463.4]
  input        io_wdata, // @[:@61463.4]
  output       io_rdata, // @[:@61463.4]
  input        io_banks_0_wdata_valid, // @[:@61463.4]
  input        io_banks_0_wdata_bits, // @[:@61463.4]
  input        io_banks_1_wdata_valid, // @[:@61463.4]
  input        io_banks_1_wdata_bits, // @[:@61463.4]
  input        io_banks_2_wdata_valid, // @[:@61463.4]
  input        io_banks_2_wdata_bits, // @[:@61463.4]
  input        io_banks_3_wdata_valid, // @[:@61463.4]
  input        io_banks_3_wdata_bits, // @[:@61463.4]
  input        io_banks_4_wdata_valid, // @[:@61463.4]
  input        io_banks_4_wdata_bits, // @[:@61463.4]
  input        io_banks_5_wdata_valid, // @[:@61463.4]
  input        io_banks_5_wdata_bits, // @[:@61463.4]
  input        io_banks_6_wdata_valid, // @[:@61463.4]
  input        io_banks_6_wdata_bits, // @[:@61463.4]
  input        io_banks_7_wdata_valid, // @[:@61463.4]
  input        io_banks_7_wdata_bits, // @[:@61463.4]
  input        io_banks_8_wdata_valid, // @[:@61463.4]
  input        io_banks_8_wdata_bits, // @[:@61463.4]
  input        io_banks_9_wdata_valid, // @[:@61463.4]
  input        io_banks_9_wdata_bits, // @[:@61463.4]
  input        io_banks_10_wdata_valid, // @[:@61463.4]
  input        io_banks_10_wdata_bits, // @[:@61463.4]
  input        io_banks_11_wdata_valid, // @[:@61463.4]
  input        io_banks_11_wdata_bits, // @[:@61463.4]
  input        io_banks_12_wdata_valid, // @[:@61463.4]
  input        io_banks_12_wdata_bits, // @[:@61463.4]
  input        io_banks_13_wdata_valid, // @[:@61463.4]
  input        io_banks_13_wdata_bits, // @[:@61463.4]
  input        io_banks_14_wdata_valid, // @[:@61463.4]
  input        io_banks_14_wdata_bits, // @[:@61463.4]
  input        io_banks_15_wdata_valid, // @[:@61463.4]
  input        io_banks_15_wdata_bits, // @[:@61463.4]
  input        io_banks_16_wdata_valid, // @[:@61463.4]
  input        io_banks_16_wdata_bits, // @[:@61463.4]
  input        io_banks_17_wdata_valid, // @[:@61463.4]
  input        io_banks_17_wdata_bits, // @[:@61463.4]
  input        io_banks_18_wdata_valid, // @[:@61463.4]
  input        io_banks_18_wdata_bits, // @[:@61463.4]
  input        io_banks_19_wdata_valid, // @[:@61463.4]
  input        io_banks_19_wdata_bits, // @[:@61463.4]
  input        io_banks_20_wdata_valid, // @[:@61463.4]
  input        io_banks_20_wdata_bits, // @[:@61463.4]
  input        io_banks_21_wdata_valid, // @[:@61463.4]
  input        io_banks_21_wdata_bits, // @[:@61463.4]
  input        io_banks_22_wdata_valid, // @[:@61463.4]
  input        io_banks_22_wdata_bits, // @[:@61463.4]
  input        io_banks_23_wdata_valid, // @[:@61463.4]
  input        io_banks_23_wdata_bits, // @[:@61463.4]
  input        io_banks_24_wdata_valid, // @[:@61463.4]
  input        io_banks_24_wdata_bits, // @[:@61463.4]
  input        io_banks_25_wdata_valid, // @[:@61463.4]
  input        io_banks_25_wdata_bits, // @[:@61463.4]
  input        io_banks_26_wdata_valid, // @[:@61463.4]
  input        io_banks_26_wdata_bits, // @[:@61463.4]
  input        io_banks_27_wdata_valid, // @[:@61463.4]
  input        io_banks_27_wdata_bits, // @[:@61463.4]
  input        io_banks_28_wdata_valid, // @[:@61463.4]
  input        io_banks_28_wdata_bits, // @[:@61463.4]
  input        io_banks_29_wdata_valid, // @[:@61463.4]
  input        io_banks_29_wdata_bits, // @[:@61463.4]
  input        io_banks_30_wdata_valid, // @[:@61463.4]
  input        io_banks_30_wdata_bits, // @[:@61463.4]
  input        io_banks_31_wdata_valid, // @[:@61463.4]
  input        io_banks_31_wdata_bits, // @[:@61463.4]
  input        io_banks_32_wdata_valid, // @[:@61463.4]
  input        io_banks_32_wdata_bits, // @[:@61463.4]
  input        io_banks_33_wdata_valid, // @[:@61463.4]
  input        io_banks_33_wdata_bits, // @[:@61463.4]
  input        io_banks_34_wdata_valid, // @[:@61463.4]
  input        io_banks_34_wdata_bits, // @[:@61463.4]
  input        io_banks_35_wdata_valid, // @[:@61463.4]
  input        io_banks_35_wdata_bits, // @[:@61463.4]
  input        io_banks_36_wdata_valid, // @[:@61463.4]
  input        io_banks_36_wdata_bits, // @[:@61463.4]
  input        io_banks_37_wdata_valid, // @[:@61463.4]
  input        io_banks_37_wdata_bits, // @[:@61463.4]
  input        io_banks_38_wdata_valid, // @[:@61463.4]
  input        io_banks_38_wdata_bits, // @[:@61463.4]
  input        io_banks_39_wdata_valid, // @[:@61463.4]
  input        io_banks_39_wdata_bits, // @[:@61463.4]
  input        io_banks_40_wdata_valid, // @[:@61463.4]
  input        io_banks_40_wdata_bits, // @[:@61463.4]
  input        io_banks_41_wdata_valid, // @[:@61463.4]
  input        io_banks_41_wdata_bits, // @[:@61463.4]
  input        io_banks_42_wdata_valid, // @[:@61463.4]
  input        io_banks_42_wdata_bits, // @[:@61463.4]
  input        io_banks_43_wdata_valid, // @[:@61463.4]
  input        io_banks_43_wdata_bits, // @[:@61463.4]
  input        io_banks_44_wdata_valid, // @[:@61463.4]
  input        io_banks_44_wdata_bits, // @[:@61463.4]
  input        io_banks_45_wdata_valid, // @[:@61463.4]
  input        io_banks_45_wdata_bits, // @[:@61463.4]
  input        io_banks_46_wdata_valid, // @[:@61463.4]
  input        io_banks_46_wdata_bits, // @[:@61463.4]
  input        io_banks_47_wdata_valid, // @[:@61463.4]
  input        io_banks_47_wdata_bits, // @[:@61463.4]
  input        io_banks_48_wdata_valid, // @[:@61463.4]
  input        io_banks_48_wdata_bits, // @[:@61463.4]
  input        io_banks_49_wdata_valid, // @[:@61463.4]
  input        io_banks_49_wdata_bits, // @[:@61463.4]
  input        io_banks_50_wdata_valid, // @[:@61463.4]
  input        io_banks_50_wdata_bits, // @[:@61463.4]
  input        io_banks_51_wdata_valid, // @[:@61463.4]
  input        io_banks_51_wdata_bits, // @[:@61463.4]
  input        io_banks_52_wdata_valid, // @[:@61463.4]
  input        io_banks_52_wdata_bits, // @[:@61463.4]
  input        io_banks_53_wdata_valid, // @[:@61463.4]
  input        io_banks_53_wdata_bits, // @[:@61463.4]
  input        io_banks_54_wdata_valid, // @[:@61463.4]
  input        io_banks_54_wdata_bits, // @[:@61463.4]
  input        io_banks_55_wdata_valid, // @[:@61463.4]
  input        io_banks_55_wdata_bits, // @[:@61463.4]
  input        io_banks_56_wdata_valid, // @[:@61463.4]
  input        io_banks_56_wdata_bits, // @[:@61463.4]
  input        io_banks_57_wdata_valid, // @[:@61463.4]
  input        io_banks_57_wdata_bits, // @[:@61463.4]
  input        io_banks_58_wdata_valid, // @[:@61463.4]
  input        io_banks_58_wdata_bits, // @[:@61463.4]
  input        io_banks_59_wdata_valid, // @[:@61463.4]
  input        io_banks_59_wdata_bits, // @[:@61463.4]
  input        io_banks_60_wdata_valid, // @[:@61463.4]
  input        io_banks_60_wdata_bits, // @[:@61463.4]
  input        io_banks_61_wdata_valid, // @[:@61463.4]
  input        io_banks_61_wdata_bits, // @[:@61463.4]
  input        io_banks_62_wdata_valid, // @[:@61463.4]
  input        io_banks_62_wdata_bits, // @[:@61463.4]
  input        io_banks_63_wdata_valid, // @[:@61463.4]
  input        io_banks_63_wdata_bits // @[:@61463.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@61467.4]
  reg [31:0] _RAND_0;
  wire  _T_688; // @[SRAM.scala 148:37:@61468.4]
  wire  _T_689; // @[SRAM.scala 148:25:@61469.4]
  wire  _T_690; // @[SRAM.scala 148:15:@61470.4]
  wire  _T_691; // @[SRAM.scala 149:15:@61472.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@61471.4]
  reg  regs_1; // @[SRAM.scala 145:20:@61478.4]
  reg [31:0] _RAND_1;
  wire  _T_697; // @[SRAM.scala 148:37:@61479.4]
  wire  _T_698; // @[SRAM.scala 148:25:@61480.4]
  wire  _T_699; // @[SRAM.scala 148:15:@61481.4]
  wire  _T_700; // @[SRAM.scala 149:15:@61483.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@61482.4]
  reg  regs_2; // @[SRAM.scala 145:20:@61489.4]
  reg [31:0] _RAND_2;
  wire  _T_706; // @[SRAM.scala 148:37:@61490.4]
  wire  _T_707; // @[SRAM.scala 148:25:@61491.4]
  wire  _T_708; // @[SRAM.scala 148:15:@61492.4]
  wire  _T_709; // @[SRAM.scala 149:15:@61494.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@61493.4]
  reg  regs_3; // @[SRAM.scala 145:20:@61500.4]
  reg [31:0] _RAND_3;
  wire  _T_715; // @[SRAM.scala 148:37:@61501.4]
  wire  _T_716; // @[SRAM.scala 148:25:@61502.4]
  wire  _T_717; // @[SRAM.scala 148:15:@61503.4]
  wire  _T_718; // @[SRAM.scala 149:15:@61505.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@61504.4]
  reg  regs_4; // @[SRAM.scala 145:20:@61511.4]
  reg [31:0] _RAND_4;
  wire  _T_724; // @[SRAM.scala 148:37:@61512.4]
  wire  _T_725; // @[SRAM.scala 148:25:@61513.4]
  wire  _T_726; // @[SRAM.scala 148:15:@61514.4]
  wire  _T_727; // @[SRAM.scala 149:15:@61516.6]
  wire  _GEN_4; // @[SRAM.scala 148:48:@61515.4]
  reg  regs_5; // @[SRAM.scala 145:20:@61522.4]
  reg [31:0] _RAND_5;
  wire  _T_733; // @[SRAM.scala 148:37:@61523.4]
  wire  _T_734; // @[SRAM.scala 148:25:@61524.4]
  wire  _T_735; // @[SRAM.scala 148:15:@61525.4]
  wire  _T_736; // @[SRAM.scala 149:15:@61527.6]
  wire  _GEN_5; // @[SRAM.scala 148:48:@61526.4]
  reg  regs_6; // @[SRAM.scala 145:20:@61533.4]
  reg [31:0] _RAND_6;
  wire  _T_742; // @[SRAM.scala 148:37:@61534.4]
  wire  _T_743; // @[SRAM.scala 148:25:@61535.4]
  wire  _T_744; // @[SRAM.scala 148:15:@61536.4]
  wire  _T_745; // @[SRAM.scala 149:15:@61538.6]
  wire  _GEN_6; // @[SRAM.scala 148:48:@61537.4]
  reg  regs_7; // @[SRAM.scala 145:20:@61544.4]
  reg [31:0] _RAND_7;
  wire  _T_751; // @[SRAM.scala 148:37:@61545.4]
  wire  _T_752; // @[SRAM.scala 148:25:@61546.4]
  wire  _T_753; // @[SRAM.scala 148:15:@61547.4]
  wire  _T_754; // @[SRAM.scala 149:15:@61549.6]
  wire  _GEN_7; // @[SRAM.scala 148:48:@61548.4]
  reg  regs_8; // @[SRAM.scala 145:20:@61555.4]
  reg [31:0] _RAND_8;
  wire  _T_760; // @[SRAM.scala 148:37:@61556.4]
  wire  _T_761; // @[SRAM.scala 148:25:@61557.4]
  wire  _T_762; // @[SRAM.scala 148:15:@61558.4]
  wire  _T_763; // @[SRAM.scala 149:15:@61560.6]
  wire  _GEN_8; // @[SRAM.scala 148:48:@61559.4]
  reg  regs_9; // @[SRAM.scala 145:20:@61566.4]
  reg [31:0] _RAND_9;
  wire  _T_769; // @[SRAM.scala 148:37:@61567.4]
  wire  _T_770; // @[SRAM.scala 148:25:@61568.4]
  wire  _T_771; // @[SRAM.scala 148:15:@61569.4]
  wire  _T_772; // @[SRAM.scala 149:15:@61571.6]
  wire  _GEN_9; // @[SRAM.scala 148:48:@61570.4]
  reg  regs_10; // @[SRAM.scala 145:20:@61577.4]
  reg [31:0] _RAND_10;
  wire  _T_778; // @[SRAM.scala 148:37:@61578.4]
  wire  _T_779; // @[SRAM.scala 148:25:@61579.4]
  wire  _T_780; // @[SRAM.scala 148:15:@61580.4]
  wire  _T_781; // @[SRAM.scala 149:15:@61582.6]
  wire  _GEN_10; // @[SRAM.scala 148:48:@61581.4]
  reg  regs_11; // @[SRAM.scala 145:20:@61588.4]
  reg [31:0] _RAND_11;
  wire  _T_787; // @[SRAM.scala 148:37:@61589.4]
  wire  _T_788; // @[SRAM.scala 148:25:@61590.4]
  wire  _T_789; // @[SRAM.scala 148:15:@61591.4]
  wire  _T_790; // @[SRAM.scala 149:15:@61593.6]
  wire  _GEN_11; // @[SRAM.scala 148:48:@61592.4]
  reg  regs_12; // @[SRAM.scala 145:20:@61599.4]
  reg [31:0] _RAND_12;
  wire  _T_796; // @[SRAM.scala 148:37:@61600.4]
  wire  _T_797; // @[SRAM.scala 148:25:@61601.4]
  wire  _T_798; // @[SRAM.scala 148:15:@61602.4]
  wire  _T_799; // @[SRAM.scala 149:15:@61604.6]
  wire  _GEN_12; // @[SRAM.scala 148:48:@61603.4]
  reg  regs_13; // @[SRAM.scala 145:20:@61610.4]
  reg [31:0] _RAND_13;
  wire  _T_805; // @[SRAM.scala 148:37:@61611.4]
  wire  _T_806; // @[SRAM.scala 148:25:@61612.4]
  wire  _T_807; // @[SRAM.scala 148:15:@61613.4]
  wire  _T_808; // @[SRAM.scala 149:15:@61615.6]
  wire  _GEN_13; // @[SRAM.scala 148:48:@61614.4]
  reg  regs_14; // @[SRAM.scala 145:20:@61621.4]
  reg [31:0] _RAND_14;
  wire  _T_814; // @[SRAM.scala 148:37:@61622.4]
  wire  _T_815; // @[SRAM.scala 148:25:@61623.4]
  wire  _T_816; // @[SRAM.scala 148:15:@61624.4]
  wire  _T_817; // @[SRAM.scala 149:15:@61626.6]
  wire  _GEN_14; // @[SRAM.scala 148:48:@61625.4]
  reg  regs_15; // @[SRAM.scala 145:20:@61632.4]
  reg [31:0] _RAND_15;
  wire  _T_823; // @[SRAM.scala 148:37:@61633.4]
  wire  _T_824; // @[SRAM.scala 148:25:@61634.4]
  wire  _T_825; // @[SRAM.scala 148:15:@61635.4]
  wire  _T_826; // @[SRAM.scala 149:15:@61637.6]
  wire  _GEN_15; // @[SRAM.scala 148:48:@61636.4]
  reg  regs_16; // @[SRAM.scala 145:20:@61643.4]
  reg [31:0] _RAND_16;
  wire  _T_832; // @[SRAM.scala 148:37:@61644.4]
  wire  _T_833; // @[SRAM.scala 148:25:@61645.4]
  wire  _T_834; // @[SRAM.scala 148:15:@61646.4]
  wire  _T_835; // @[SRAM.scala 149:15:@61648.6]
  wire  _GEN_16; // @[SRAM.scala 148:48:@61647.4]
  reg  regs_17; // @[SRAM.scala 145:20:@61654.4]
  reg [31:0] _RAND_17;
  wire  _T_841; // @[SRAM.scala 148:37:@61655.4]
  wire  _T_842; // @[SRAM.scala 148:25:@61656.4]
  wire  _T_843; // @[SRAM.scala 148:15:@61657.4]
  wire  _T_844; // @[SRAM.scala 149:15:@61659.6]
  wire  _GEN_17; // @[SRAM.scala 148:48:@61658.4]
  reg  regs_18; // @[SRAM.scala 145:20:@61665.4]
  reg [31:0] _RAND_18;
  wire  _T_850; // @[SRAM.scala 148:37:@61666.4]
  wire  _T_851; // @[SRAM.scala 148:25:@61667.4]
  wire  _T_852; // @[SRAM.scala 148:15:@61668.4]
  wire  _T_853; // @[SRAM.scala 149:15:@61670.6]
  wire  _GEN_18; // @[SRAM.scala 148:48:@61669.4]
  reg  regs_19; // @[SRAM.scala 145:20:@61676.4]
  reg [31:0] _RAND_19;
  wire  _T_859; // @[SRAM.scala 148:37:@61677.4]
  wire  _T_860; // @[SRAM.scala 148:25:@61678.4]
  wire  _T_861; // @[SRAM.scala 148:15:@61679.4]
  wire  _T_862; // @[SRAM.scala 149:15:@61681.6]
  wire  _GEN_19; // @[SRAM.scala 148:48:@61680.4]
  reg  regs_20; // @[SRAM.scala 145:20:@61687.4]
  reg [31:0] _RAND_20;
  wire  _T_868; // @[SRAM.scala 148:37:@61688.4]
  wire  _T_869; // @[SRAM.scala 148:25:@61689.4]
  wire  _T_870; // @[SRAM.scala 148:15:@61690.4]
  wire  _T_871; // @[SRAM.scala 149:15:@61692.6]
  wire  _GEN_20; // @[SRAM.scala 148:48:@61691.4]
  reg  regs_21; // @[SRAM.scala 145:20:@61698.4]
  reg [31:0] _RAND_21;
  wire  _T_877; // @[SRAM.scala 148:37:@61699.4]
  wire  _T_878; // @[SRAM.scala 148:25:@61700.4]
  wire  _T_879; // @[SRAM.scala 148:15:@61701.4]
  wire  _T_880; // @[SRAM.scala 149:15:@61703.6]
  wire  _GEN_21; // @[SRAM.scala 148:48:@61702.4]
  reg  regs_22; // @[SRAM.scala 145:20:@61709.4]
  reg [31:0] _RAND_22;
  wire  _T_886; // @[SRAM.scala 148:37:@61710.4]
  wire  _T_887; // @[SRAM.scala 148:25:@61711.4]
  wire  _T_888; // @[SRAM.scala 148:15:@61712.4]
  wire  _T_889; // @[SRAM.scala 149:15:@61714.6]
  wire  _GEN_22; // @[SRAM.scala 148:48:@61713.4]
  reg  regs_23; // @[SRAM.scala 145:20:@61720.4]
  reg [31:0] _RAND_23;
  wire  _T_895; // @[SRAM.scala 148:37:@61721.4]
  wire  _T_896; // @[SRAM.scala 148:25:@61722.4]
  wire  _T_897; // @[SRAM.scala 148:15:@61723.4]
  wire  _T_898; // @[SRAM.scala 149:15:@61725.6]
  wire  _GEN_23; // @[SRAM.scala 148:48:@61724.4]
  reg  regs_24; // @[SRAM.scala 145:20:@61731.4]
  reg [31:0] _RAND_24;
  wire  _T_904; // @[SRAM.scala 148:37:@61732.4]
  wire  _T_905; // @[SRAM.scala 148:25:@61733.4]
  wire  _T_906; // @[SRAM.scala 148:15:@61734.4]
  wire  _T_907; // @[SRAM.scala 149:15:@61736.6]
  wire  _GEN_24; // @[SRAM.scala 148:48:@61735.4]
  reg  regs_25; // @[SRAM.scala 145:20:@61742.4]
  reg [31:0] _RAND_25;
  wire  _T_913; // @[SRAM.scala 148:37:@61743.4]
  wire  _T_914; // @[SRAM.scala 148:25:@61744.4]
  wire  _T_915; // @[SRAM.scala 148:15:@61745.4]
  wire  _T_916; // @[SRAM.scala 149:15:@61747.6]
  wire  _GEN_25; // @[SRAM.scala 148:48:@61746.4]
  reg  regs_26; // @[SRAM.scala 145:20:@61753.4]
  reg [31:0] _RAND_26;
  wire  _T_922; // @[SRAM.scala 148:37:@61754.4]
  wire  _T_923; // @[SRAM.scala 148:25:@61755.4]
  wire  _T_924; // @[SRAM.scala 148:15:@61756.4]
  wire  _T_925; // @[SRAM.scala 149:15:@61758.6]
  wire  _GEN_26; // @[SRAM.scala 148:48:@61757.4]
  reg  regs_27; // @[SRAM.scala 145:20:@61764.4]
  reg [31:0] _RAND_27;
  wire  _T_931; // @[SRAM.scala 148:37:@61765.4]
  wire  _T_932; // @[SRAM.scala 148:25:@61766.4]
  wire  _T_933; // @[SRAM.scala 148:15:@61767.4]
  wire  _T_934; // @[SRAM.scala 149:15:@61769.6]
  wire  _GEN_27; // @[SRAM.scala 148:48:@61768.4]
  reg  regs_28; // @[SRAM.scala 145:20:@61775.4]
  reg [31:0] _RAND_28;
  wire  _T_940; // @[SRAM.scala 148:37:@61776.4]
  wire  _T_941; // @[SRAM.scala 148:25:@61777.4]
  wire  _T_942; // @[SRAM.scala 148:15:@61778.4]
  wire  _T_943; // @[SRAM.scala 149:15:@61780.6]
  wire  _GEN_28; // @[SRAM.scala 148:48:@61779.4]
  reg  regs_29; // @[SRAM.scala 145:20:@61786.4]
  reg [31:0] _RAND_29;
  wire  _T_949; // @[SRAM.scala 148:37:@61787.4]
  wire  _T_950; // @[SRAM.scala 148:25:@61788.4]
  wire  _T_951; // @[SRAM.scala 148:15:@61789.4]
  wire  _T_952; // @[SRAM.scala 149:15:@61791.6]
  wire  _GEN_29; // @[SRAM.scala 148:48:@61790.4]
  reg  regs_30; // @[SRAM.scala 145:20:@61797.4]
  reg [31:0] _RAND_30;
  wire  _T_958; // @[SRAM.scala 148:37:@61798.4]
  wire  _T_959; // @[SRAM.scala 148:25:@61799.4]
  wire  _T_960; // @[SRAM.scala 148:15:@61800.4]
  wire  _T_961; // @[SRAM.scala 149:15:@61802.6]
  wire  _GEN_30; // @[SRAM.scala 148:48:@61801.4]
  reg  regs_31; // @[SRAM.scala 145:20:@61808.4]
  reg [31:0] _RAND_31;
  wire  _T_967; // @[SRAM.scala 148:37:@61809.4]
  wire  _T_968; // @[SRAM.scala 148:25:@61810.4]
  wire  _T_969; // @[SRAM.scala 148:15:@61811.4]
  wire  _T_970; // @[SRAM.scala 149:15:@61813.6]
  wire  _GEN_31; // @[SRAM.scala 148:48:@61812.4]
  reg  regs_32; // @[SRAM.scala 145:20:@61819.4]
  reg [31:0] _RAND_32;
  wire  _T_976; // @[SRAM.scala 148:37:@61820.4]
  wire  _T_977; // @[SRAM.scala 148:25:@61821.4]
  wire  _T_978; // @[SRAM.scala 148:15:@61822.4]
  wire  _T_979; // @[SRAM.scala 149:15:@61824.6]
  wire  _GEN_32; // @[SRAM.scala 148:48:@61823.4]
  reg  regs_33; // @[SRAM.scala 145:20:@61830.4]
  reg [31:0] _RAND_33;
  wire  _T_985; // @[SRAM.scala 148:37:@61831.4]
  wire  _T_986; // @[SRAM.scala 148:25:@61832.4]
  wire  _T_987; // @[SRAM.scala 148:15:@61833.4]
  wire  _T_988; // @[SRAM.scala 149:15:@61835.6]
  wire  _GEN_33; // @[SRAM.scala 148:48:@61834.4]
  reg  regs_34; // @[SRAM.scala 145:20:@61841.4]
  reg [31:0] _RAND_34;
  wire  _T_994; // @[SRAM.scala 148:37:@61842.4]
  wire  _T_995; // @[SRAM.scala 148:25:@61843.4]
  wire  _T_996; // @[SRAM.scala 148:15:@61844.4]
  wire  _T_997; // @[SRAM.scala 149:15:@61846.6]
  wire  _GEN_34; // @[SRAM.scala 148:48:@61845.4]
  reg  regs_35; // @[SRAM.scala 145:20:@61852.4]
  reg [31:0] _RAND_35;
  wire  _T_1003; // @[SRAM.scala 148:37:@61853.4]
  wire  _T_1004; // @[SRAM.scala 148:25:@61854.4]
  wire  _T_1005; // @[SRAM.scala 148:15:@61855.4]
  wire  _T_1006; // @[SRAM.scala 149:15:@61857.6]
  wire  _GEN_35; // @[SRAM.scala 148:48:@61856.4]
  reg  regs_36; // @[SRAM.scala 145:20:@61863.4]
  reg [31:0] _RAND_36;
  wire  _T_1012; // @[SRAM.scala 148:37:@61864.4]
  wire  _T_1013; // @[SRAM.scala 148:25:@61865.4]
  wire  _T_1014; // @[SRAM.scala 148:15:@61866.4]
  wire  _T_1015; // @[SRAM.scala 149:15:@61868.6]
  wire  _GEN_36; // @[SRAM.scala 148:48:@61867.4]
  reg  regs_37; // @[SRAM.scala 145:20:@61874.4]
  reg [31:0] _RAND_37;
  wire  _T_1021; // @[SRAM.scala 148:37:@61875.4]
  wire  _T_1022; // @[SRAM.scala 148:25:@61876.4]
  wire  _T_1023; // @[SRAM.scala 148:15:@61877.4]
  wire  _T_1024; // @[SRAM.scala 149:15:@61879.6]
  wire  _GEN_37; // @[SRAM.scala 148:48:@61878.4]
  reg  regs_38; // @[SRAM.scala 145:20:@61885.4]
  reg [31:0] _RAND_38;
  wire  _T_1030; // @[SRAM.scala 148:37:@61886.4]
  wire  _T_1031; // @[SRAM.scala 148:25:@61887.4]
  wire  _T_1032; // @[SRAM.scala 148:15:@61888.4]
  wire  _T_1033; // @[SRAM.scala 149:15:@61890.6]
  wire  _GEN_38; // @[SRAM.scala 148:48:@61889.4]
  reg  regs_39; // @[SRAM.scala 145:20:@61896.4]
  reg [31:0] _RAND_39;
  wire  _T_1039; // @[SRAM.scala 148:37:@61897.4]
  wire  _T_1040; // @[SRAM.scala 148:25:@61898.4]
  wire  _T_1041; // @[SRAM.scala 148:15:@61899.4]
  wire  _T_1042; // @[SRAM.scala 149:15:@61901.6]
  wire  _GEN_39; // @[SRAM.scala 148:48:@61900.4]
  reg  regs_40; // @[SRAM.scala 145:20:@61907.4]
  reg [31:0] _RAND_40;
  wire  _T_1048; // @[SRAM.scala 148:37:@61908.4]
  wire  _T_1049; // @[SRAM.scala 148:25:@61909.4]
  wire  _T_1050; // @[SRAM.scala 148:15:@61910.4]
  wire  _T_1051; // @[SRAM.scala 149:15:@61912.6]
  wire  _GEN_40; // @[SRAM.scala 148:48:@61911.4]
  reg  regs_41; // @[SRAM.scala 145:20:@61918.4]
  reg [31:0] _RAND_41;
  wire  _T_1057; // @[SRAM.scala 148:37:@61919.4]
  wire  _T_1058; // @[SRAM.scala 148:25:@61920.4]
  wire  _T_1059; // @[SRAM.scala 148:15:@61921.4]
  wire  _T_1060; // @[SRAM.scala 149:15:@61923.6]
  wire  _GEN_41; // @[SRAM.scala 148:48:@61922.4]
  reg  regs_42; // @[SRAM.scala 145:20:@61929.4]
  reg [31:0] _RAND_42;
  wire  _T_1066; // @[SRAM.scala 148:37:@61930.4]
  wire  _T_1067; // @[SRAM.scala 148:25:@61931.4]
  wire  _T_1068; // @[SRAM.scala 148:15:@61932.4]
  wire  _T_1069; // @[SRAM.scala 149:15:@61934.6]
  wire  _GEN_42; // @[SRAM.scala 148:48:@61933.4]
  reg  regs_43; // @[SRAM.scala 145:20:@61940.4]
  reg [31:0] _RAND_43;
  wire  _T_1075; // @[SRAM.scala 148:37:@61941.4]
  wire  _T_1076; // @[SRAM.scala 148:25:@61942.4]
  wire  _T_1077; // @[SRAM.scala 148:15:@61943.4]
  wire  _T_1078; // @[SRAM.scala 149:15:@61945.6]
  wire  _GEN_43; // @[SRAM.scala 148:48:@61944.4]
  reg  regs_44; // @[SRAM.scala 145:20:@61951.4]
  reg [31:0] _RAND_44;
  wire  _T_1084; // @[SRAM.scala 148:37:@61952.4]
  wire  _T_1085; // @[SRAM.scala 148:25:@61953.4]
  wire  _T_1086; // @[SRAM.scala 148:15:@61954.4]
  wire  _T_1087; // @[SRAM.scala 149:15:@61956.6]
  wire  _GEN_44; // @[SRAM.scala 148:48:@61955.4]
  reg  regs_45; // @[SRAM.scala 145:20:@61962.4]
  reg [31:0] _RAND_45;
  wire  _T_1093; // @[SRAM.scala 148:37:@61963.4]
  wire  _T_1094; // @[SRAM.scala 148:25:@61964.4]
  wire  _T_1095; // @[SRAM.scala 148:15:@61965.4]
  wire  _T_1096; // @[SRAM.scala 149:15:@61967.6]
  wire  _GEN_45; // @[SRAM.scala 148:48:@61966.4]
  reg  regs_46; // @[SRAM.scala 145:20:@61973.4]
  reg [31:0] _RAND_46;
  wire  _T_1102; // @[SRAM.scala 148:37:@61974.4]
  wire  _T_1103; // @[SRAM.scala 148:25:@61975.4]
  wire  _T_1104; // @[SRAM.scala 148:15:@61976.4]
  wire  _T_1105; // @[SRAM.scala 149:15:@61978.6]
  wire  _GEN_46; // @[SRAM.scala 148:48:@61977.4]
  reg  regs_47; // @[SRAM.scala 145:20:@61984.4]
  reg [31:0] _RAND_47;
  wire  _T_1111; // @[SRAM.scala 148:37:@61985.4]
  wire  _T_1112; // @[SRAM.scala 148:25:@61986.4]
  wire  _T_1113; // @[SRAM.scala 148:15:@61987.4]
  wire  _T_1114; // @[SRAM.scala 149:15:@61989.6]
  wire  _GEN_47; // @[SRAM.scala 148:48:@61988.4]
  reg  regs_48; // @[SRAM.scala 145:20:@61995.4]
  reg [31:0] _RAND_48;
  wire  _T_1120; // @[SRAM.scala 148:37:@61996.4]
  wire  _T_1121; // @[SRAM.scala 148:25:@61997.4]
  wire  _T_1122; // @[SRAM.scala 148:15:@61998.4]
  wire  _T_1123; // @[SRAM.scala 149:15:@62000.6]
  wire  _GEN_48; // @[SRAM.scala 148:48:@61999.4]
  reg  regs_49; // @[SRAM.scala 145:20:@62006.4]
  reg [31:0] _RAND_49;
  wire  _T_1129; // @[SRAM.scala 148:37:@62007.4]
  wire  _T_1130; // @[SRAM.scala 148:25:@62008.4]
  wire  _T_1131; // @[SRAM.scala 148:15:@62009.4]
  wire  _T_1132; // @[SRAM.scala 149:15:@62011.6]
  wire  _GEN_49; // @[SRAM.scala 148:48:@62010.4]
  reg  regs_50; // @[SRAM.scala 145:20:@62017.4]
  reg [31:0] _RAND_50;
  wire  _T_1138; // @[SRAM.scala 148:37:@62018.4]
  wire  _T_1139; // @[SRAM.scala 148:25:@62019.4]
  wire  _T_1140; // @[SRAM.scala 148:15:@62020.4]
  wire  _T_1141; // @[SRAM.scala 149:15:@62022.6]
  wire  _GEN_50; // @[SRAM.scala 148:48:@62021.4]
  reg  regs_51; // @[SRAM.scala 145:20:@62028.4]
  reg [31:0] _RAND_51;
  wire  _T_1147; // @[SRAM.scala 148:37:@62029.4]
  wire  _T_1148; // @[SRAM.scala 148:25:@62030.4]
  wire  _T_1149; // @[SRAM.scala 148:15:@62031.4]
  wire  _T_1150; // @[SRAM.scala 149:15:@62033.6]
  wire  _GEN_51; // @[SRAM.scala 148:48:@62032.4]
  reg  regs_52; // @[SRAM.scala 145:20:@62039.4]
  reg [31:0] _RAND_52;
  wire  _T_1156; // @[SRAM.scala 148:37:@62040.4]
  wire  _T_1157; // @[SRAM.scala 148:25:@62041.4]
  wire  _T_1158; // @[SRAM.scala 148:15:@62042.4]
  wire  _T_1159; // @[SRAM.scala 149:15:@62044.6]
  wire  _GEN_52; // @[SRAM.scala 148:48:@62043.4]
  reg  regs_53; // @[SRAM.scala 145:20:@62050.4]
  reg [31:0] _RAND_53;
  wire  _T_1165; // @[SRAM.scala 148:37:@62051.4]
  wire  _T_1166; // @[SRAM.scala 148:25:@62052.4]
  wire  _T_1167; // @[SRAM.scala 148:15:@62053.4]
  wire  _T_1168; // @[SRAM.scala 149:15:@62055.6]
  wire  _GEN_53; // @[SRAM.scala 148:48:@62054.4]
  reg  regs_54; // @[SRAM.scala 145:20:@62061.4]
  reg [31:0] _RAND_54;
  wire  _T_1174; // @[SRAM.scala 148:37:@62062.4]
  wire  _T_1175; // @[SRAM.scala 148:25:@62063.4]
  wire  _T_1176; // @[SRAM.scala 148:15:@62064.4]
  wire  _T_1177; // @[SRAM.scala 149:15:@62066.6]
  wire  _GEN_54; // @[SRAM.scala 148:48:@62065.4]
  reg  regs_55; // @[SRAM.scala 145:20:@62072.4]
  reg [31:0] _RAND_55;
  wire  _T_1183; // @[SRAM.scala 148:37:@62073.4]
  wire  _T_1184; // @[SRAM.scala 148:25:@62074.4]
  wire  _T_1185; // @[SRAM.scala 148:15:@62075.4]
  wire  _T_1186; // @[SRAM.scala 149:15:@62077.6]
  wire  _GEN_55; // @[SRAM.scala 148:48:@62076.4]
  reg  regs_56; // @[SRAM.scala 145:20:@62083.4]
  reg [31:0] _RAND_56;
  wire  _T_1192; // @[SRAM.scala 148:37:@62084.4]
  wire  _T_1193; // @[SRAM.scala 148:25:@62085.4]
  wire  _T_1194; // @[SRAM.scala 148:15:@62086.4]
  wire  _T_1195; // @[SRAM.scala 149:15:@62088.6]
  wire  _GEN_56; // @[SRAM.scala 148:48:@62087.4]
  reg  regs_57; // @[SRAM.scala 145:20:@62094.4]
  reg [31:0] _RAND_57;
  wire  _T_1201; // @[SRAM.scala 148:37:@62095.4]
  wire  _T_1202; // @[SRAM.scala 148:25:@62096.4]
  wire  _T_1203; // @[SRAM.scala 148:15:@62097.4]
  wire  _T_1204; // @[SRAM.scala 149:15:@62099.6]
  wire  _GEN_57; // @[SRAM.scala 148:48:@62098.4]
  reg  regs_58; // @[SRAM.scala 145:20:@62105.4]
  reg [31:0] _RAND_58;
  wire  _T_1210; // @[SRAM.scala 148:37:@62106.4]
  wire  _T_1211; // @[SRAM.scala 148:25:@62107.4]
  wire  _T_1212; // @[SRAM.scala 148:15:@62108.4]
  wire  _T_1213; // @[SRAM.scala 149:15:@62110.6]
  wire  _GEN_58; // @[SRAM.scala 148:48:@62109.4]
  reg  regs_59; // @[SRAM.scala 145:20:@62116.4]
  reg [31:0] _RAND_59;
  wire  _T_1219; // @[SRAM.scala 148:37:@62117.4]
  wire  _T_1220; // @[SRAM.scala 148:25:@62118.4]
  wire  _T_1221; // @[SRAM.scala 148:15:@62119.4]
  wire  _T_1222; // @[SRAM.scala 149:15:@62121.6]
  wire  _GEN_59; // @[SRAM.scala 148:48:@62120.4]
  reg  regs_60; // @[SRAM.scala 145:20:@62127.4]
  reg [31:0] _RAND_60;
  wire  _T_1228; // @[SRAM.scala 148:37:@62128.4]
  wire  _T_1229; // @[SRAM.scala 148:25:@62129.4]
  wire  _T_1230; // @[SRAM.scala 148:15:@62130.4]
  wire  _T_1231; // @[SRAM.scala 149:15:@62132.6]
  wire  _GEN_60; // @[SRAM.scala 148:48:@62131.4]
  reg  regs_61; // @[SRAM.scala 145:20:@62138.4]
  reg [31:0] _RAND_61;
  wire  _T_1237; // @[SRAM.scala 148:37:@62139.4]
  wire  _T_1238; // @[SRAM.scala 148:25:@62140.4]
  wire  _T_1239; // @[SRAM.scala 148:15:@62141.4]
  wire  _T_1240; // @[SRAM.scala 149:15:@62143.6]
  wire  _GEN_61; // @[SRAM.scala 148:48:@62142.4]
  reg  regs_62; // @[SRAM.scala 145:20:@62149.4]
  reg [31:0] _RAND_62;
  wire  _T_1246; // @[SRAM.scala 148:37:@62150.4]
  wire  _T_1247; // @[SRAM.scala 148:25:@62151.4]
  wire  _T_1248; // @[SRAM.scala 148:15:@62152.4]
  wire  _T_1249; // @[SRAM.scala 149:15:@62154.6]
  wire  _GEN_62; // @[SRAM.scala 148:48:@62153.4]
  reg  regs_63; // @[SRAM.scala 145:20:@62160.4]
  reg [31:0] _RAND_63;
  wire  _T_1255; // @[SRAM.scala 148:37:@62161.4]
  wire  _T_1256; // @[SRAM.scala 148:25:@62162.4]
  wire  _T_1257; // @[SRAM.scala 148:15:@62163.4]
  wire  _T_1258; // @[SRAM.scala 149:15:@62165.6]
  wire  _GEN_63; // @[SRAM.scala 148:48:@62164.4]
  wire  _GEN_65; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_66; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_67; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_68; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_69; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_70; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_71; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_72; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_73; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_74; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_75; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_76; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_77; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_78; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_79; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_80; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_81; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_82; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_83; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_84; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_85; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_86; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_87; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_88; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_89; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_90; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_91; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_92; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_93; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_94; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_95; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_96; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_97; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_98; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_99; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_100; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_101; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_102; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_103; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_104; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_105; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_106; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_107; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_108; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_109; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_110; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_111; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_112; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_113; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_114; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_115; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_116; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_117; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_118; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_119; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_120; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_121; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_122; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_123; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_124; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_125; // @[SRAM.scala 155:12:@62234.4]
  wire  _GEN_126; // @[SRAM.scala 155:12:@62234.4]
  assign _T_688 = io_waddr == 6'h0; // @[SRAM.scala 148:37:@61468.4]
  assign _T_689 = io_wen & _T_688; // @[SRAM.scala 148:25:@61469.4]
  assign _T_690 = io_banks_0_wdata_valid | _T_689; // @[SRAM.scala 148:15:@61470.4]
  assign _T_691 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61472.6]
  assign _GEN_0 = _T_690 ? _T_691 : regs_0; // @[SRAM.scala 148:48:@61471.4]
  assign _T_697 = io_waddr == 6'h1; // @[SRAM.scala 148:37:@61479.4]
  assign _T_698 = io_wen & _T_697; // @[SRAM.scala 148:25:@61480.4]
  assign _T_699 = io_banks_1_wdata_valid | _T_698; // @[SRAM.scala 148:15:@61481.4]
  assign _T_700 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61483.6]
  assign _GEN_1 = _T_699 ? _T_700 : regs_1; // @[SRAM.scala 148:48:@61482.4]
  assign _T_706 = io_waddr == 6'h2; // @[SRAM.scala 148:37:@61490.4]
  assign _T_707 = io_wen & _T_706; // @[SRAM.scala 148:25:@61491.4]
  assign _T_708 = io_banks_2_wdata_valid | _T_707; // @[SRAM.scala 148:15:@61492.4]
  assign _T_709 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61494.6]
  assign _GEN_2 = _T_708 ? _T_709 : regs_2; // @[SRAM.scala 148:48:@61493.4]
  assign _T_715 = io_waddr == 6'h3; // @[SRAM.scala 148:37:@61501.4]
  assign _T_716 = io_wen & _T_715; // @[SRAM.scala 148:25:@61502.4]
  assign _T_717 = io_banks_3_wdata_valid | _T_716; // @[SRAM.scala 148:15:@61503.4]
  assign _T_718 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61505.6]
  assign _GEN_3 = _T_717 ? _T_718 : regs_3; // @[SRAM.scala 148:48:@61504.4]
  assign _T_724 = io_waddr == 6'h4; // @[SRAM.scala 148:37:@61512.4]
  assign _T_725 = io_wen & _T_724; // @[SRAM.scala 148:25:@61513.4]
  assign _T_726 = io_banks_4_wdata_valid | _T_725; // @[SRAM.scala 148:15:@61514.4]
  assign _T_727 = io_banks_4_wdata_valid ? io_banks_4_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61516.6]
  assign _GEN_4 = _T_726 ? _T_727 : regs_4; // @[SRAM.scala 148:48:@61515.4]
  assign _T_733 = io_waddr == 6'h5; // @[SRAM.scala 148:37:@61523.4]
  assign _T_734 = io_wen & _T_733; // @[SRAM.scala 148:25:@61524.4]
  assign _T_735 = io_banks_5_wdata_valid | _T_734; // @[SRAM.scala 148:15:@61525.4]
  assign _T_736 = io_banks_5_wdata_valid ? io_banks_5_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61527.6]
  assign _GEN_5 = _T_735 ? _T_736 : regs_5; // @[SRAM.scala 148:48:@61526.4]
  assign _T_742 = io_waddr == 6'h6; // @[SRAM.scala 148:37:@61534.4]
  assign _T_743 = io_wen & _T_742; // @[SRAM.scala 148:25:@61535.4]
  assign _T_744 = io_banks_6_wdata_valid | _T_743; // @[SRAM.scala 148:15:@61536.4]
  assign _T_745 = io_banks_6_wdata_valid ? io_banks_6_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61538.6]
  assign _GEN_6 = _T_744 ? _T_745 : regs_6; // @[SRAM.scala 148:48:@61537.4]
  assign _T_751 = io_waddr == 6'h7; // @[SRAM.scala 148:37:@61545.4]
  assign _T_752 = io_wen & _T_751; // @[SRAM.scala 148:25:@61546.4]
  assign _T_753 = io_banks_7_wdata_valid | _T_752; // @[SRAM.scala 148:15:@61547.4]
  assign _T_754 = io_banks_7_wdata_valid ? io_banks_7_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61549.6]
  assign _GEN_7 = _T_753 ? _T_754 : regs_7; // @[SRAM.scala 148:48:@61548.4]
  assign _T_760 = io_waddr == 6'h8; // @[SRAM.scala 148:37:@61556.4]
  assign _T_761 = io_wen & _T_760; // @[SRAM.scala 148:25:@61557.4]
  assign _T_762 = io_banks_8_wdata_valid | _T_761; // @[SRAM.scala 148:15:@61558.4]
  assign _T_763 = io_banks_8_wdata_valid ? io_banks_8_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61560.6]
  assign _GEN_8 = _T_762 ? _T_763 : regs_8; // @[SRAM.scala 148:48:@61559.4]
  assign _T_769 = io_waddr == 6'h9; // @[SRAM.scala 148:37:@61567.4]
  assign _T_770 = io_wen & _T_769; // @[SRAM.scala 148:25:@61568.4]
  assign _T_771 = io_banks_9_wdata_valid | _T_770; // @[SRAM.scala 148:15:@61569.4]
  assign _T_772 = io_banks_9_wdata_valid ? io_banks_9_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61571.6]
  assign _GEN_9 = _T_771 ? _T_772 : regs_9; // @[SRAM.scala 148:48:@61570.4]
  assign _T_778 = io_waddr == 6'ha; // @[SRAM.scala 148:37:@61578.4]
  assign _T_779 = io_wen & _T_778; // @[SRAM.scala 148:25:@61579.4]
  assign _T_780 = io_banks_10_wdata_valid | _T_779; // @[SRAM.scala 148:15:@61580.4]
  assign _T_781 = io_banks_10_wdata_valid ? io_banks_10_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61582.6]
  assign _GEN_10 = _T_780 ? _T_781 : regs_10; // @[SRAM.scala 148:48:@61581.4]
  assign _T_787 = io_waddr == 6'hb; // @[SRAM.scala 148:37:@61589.4]
  assign _T_788 = io_wen & _T_787; // @[SRAM.scala 148:25:@61590.4]
  assign _T_789 = io_banks_11_wdata_valid | _T_788; // @[SRAM.scala 148:15:@61591.4]
  assign _T_790 = io_banks_11_wdata_valid ? io_banks_11_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61593.6]
  assign _GEN_11 = _T_789 ? _T_790 : regs_11; // @[SRAM.scala 148:48:@61592.4]
  assign _T_796 = io_waddr == 6'hc; // @[SRAM.scala 148:37:@61600.4]
  assign _T_797 = io_wen & _T_796; // @[SRAM.scala 148:25:@61601.4]
  assign _T_798 = io_banks_12_wdata_valid | _T_797; // @[SRAM.scala 148:15:@61602.4]
  assign _T_799 = io_banks_12_wdata_valid ? io_banks_12_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61604.6]
  assign _GEN_12 = _T_798 ? _T_799 : regs_12; // @[SRAM.scala 148:48:@61603.4]
  assign _T_805 = io_waddr == 6'hd; // @[SRAM.scala 148:37:@61611.4]
  assign _T_806 = io_wen & _T_805; // @[SRAM.scala 148:25:@61612.4]
  assign _T_807 = io_banks_13_wdata_valid | _T_806; // @[SRAM.scala 148:15:@61613.4]
  assign _T_808 = io_banks_13_wdata_valid ? io_banks_13_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61615.6]
  assign _GEN_13 = _T_807 ? _T_808 : regs_13; // @[SRAM.scala 148:48:@61614.4]
  assign _T_814 = io_waddr == 6'he; // @[SRAM.scala 148:37:@61622.4]
  assign _T_815 = io_wen & _T_814; // @[SRAM.scala 148:25:@61623.4]
  assign _T_816 = io_banks_14_wdata_valid | _T_815; // @[SRAM.scala 148:15:@61624.4]
  assign _T_817 = io_banks_14_wdata_valid ? io_banks_14_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61626.6]
  assign _GEN_14 = _T_816 ? _T_817 : regs_14; // @[SRAM.scala 148:48:@61625.4]
  assign _T_823 = io_waddr == 6'hf; // @[SRAM.scala 148:37:@61633.4]
  assign _T_824 = io_wen & _T_823; // @[SRAM.scala 148:25:@61634.4]
  assign _T_825 = io_banks_15_wdata_valid | _T_824; // @[SRAM.scala 148:15:@61635.4]
  assign _T_826 = io_banks_15_wdata_valid ? io_banks_15_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61637.6]
  assign _GEN_15 = _T_825 ? _T_826 : regs_15; // @[SRAM.scala 148:48:@61636.4]
  assign _T_832 = io_waddr == 6'h10; // @[SRAM.scala 148:37:@61644.4]
  assign _T_833 = io_wen & _T_832; // @[SRAM.scala 148:25:@61645.4]
  assign _T_834 = io_banks_16_wdata_valid | _T_833; // @[SRAM.scala 148:15:@61646.4]
  assign _T_835 = io_banks_16_wdata_valid ? io_banks_16_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61648.6]
  assign _GEN_16 = _T_834 ? _T_835 : regs_16; // @[SRAM.scala 148:48:@61647.4]
  assign _T_841 = io_waddr == 6'h11; // @[SRAM.scala 148:37:@61655.4]
  assign _T_842 = io_wen & _T_841; // @[SRAM.scala 148:25:@61656.4]
  assign _T_843 = io_banks_17_wdata_valid | _T_842; // @[SRAM.scala 148:15:@61657.4]
  assign _T_844 = io_banks_17_wdata_valid ? io_banks_17_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61659.6]
  assign _GEN_17 = _T_843 ? _T_844 : regs_17; // @[SRAM.scala 148:48:@61658.4]
  assign _T_850 = io_waddr == 6'h12; // @[SRAM.scala 148:37:@61666.4]
  assign _T_851 = io_wen & _T_850; // @[SRAM.scala 148:25:@61667.4]
  assign _T_852 = io_banks_18_wdata_valid | _T_851; // @[SRAM.scala 148:15:@61668.4]
  assign _T_853 = io_banks_18_wdata_valid ? io_banks_18_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61670.6]
  assign _GEN_18 = _T_852 ? _T_853 : regs_18; // @[SRAM.scala 148:48:@61669.4]
  assign _T_859 = io_waddr == 6'h13; // @[SRAM.scala 148:37:@61677.4]
  assign _T_860 = io_wen & _T_859; // @[SRAM.scala 148:25:@61678.4]
  assign _T_861 = io_banks_19_wdata_valid | _T_860; // @[SRAM.scala 148:15:@61679.4]
  assign _T_862 = io_banks_19_wdata_valid ? io_banks_19_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61681.6]
  assign _GEN_19 = _T_861 ? _T_862 : regs_19; // @[SRAM.scala 148:48:@61680.4]
  assign _T_868 = io_waddr == 6'h14; // @[SRAM.scala 148:37:@61688.4]
  assign _T_869 = io_wen & _T_868; // @[SRAM.scala 148:25:@61689.4]
  assign _T_870 = io_banks_20_wdata_valid | _T_869; // @[SRAM.scala 148:15:@61690.4]
  assign _T_871 = io_banks_20_wdata_valid ? io_banks_20_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61692.6]
  assign _GEN_20 = _T_870 ? _T_871 : regs_20; // @[SRAM.scala 148:48:@61691.4]
  assign _T_877 = io_waddr == 6'h15; // @[SRAM.scala 148:37:@61699.4]
  assign _T_878 = io_wen & _T_877; // @[SRAM.scala 148:25:@61700.4]
  assign _T_879 = io_banks_21_wdata_valid | _T_878; // @[SRAM.scala 148:15:@61701.4]
  assign _T_880 = io_banks_21_wdata_valid ? io_banks_21_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61703.6]
  assign _GEN_21 = _T_879 ? _T_880 : regs_21; // @[SRAM.scala 148:48:@61702.4]
  assign _T_886 = io_waddr == 6'h16; // @[SRAM.scala 148:37:@61710.4]
  assign _T_887 = io_wen & _T_886; // @[SRAM.scala 148:25:@61711.4]
  assign _T_888 = io_banks_22_wdata_valid | _T_887; // @[SRAM.scala 148:15:@61712.4]
  assign _T_889 = io_banks_22_wdata_valid ? io_banks_22_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61714.6]
  assign _GEN_22 = _T_888 ? _T_889 : regs_22; // @[SRAM.scala 148:48:@61713.4]
  assign _T_895 = io_waddr == 6'h17; // @[SRAM.scala 148:37:@61721.4]
  assign _T_896 = io_wen & _T_895; // @[SRAM.scala 148:25:@61722.4]
  assign _T_897 = io_banks_23_wdata_valid | _T_896; // @[SRAM.scala 148:15:@61723.4]
  assign _T_898 = io_banks_23_wdata_valid ? io_banks_23_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61725.6]
  assign _GEN_23 = _T_897 ? _T_898 : regs_23; // @[SRAM.scala 148:48:@61724.4]
  assign _T_904 = io_waddr == 6'h18; // @[SRAM.scala 148:37:@61732.4]
  assign _T_905 = io_wen & _T_904; // @[SRAM.scala 148:25:@61733.4]
  assign _T_906 = io_banks_24_wdata_valid | _T_905; // @[SRAM.scala 148:15:@61734.4]
  assign _T_907 = io_banks_24_wdata_valid ? io_banks_24_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61736.6]
  assign _GEN_24 = _T_906 ? _T_907 : regs_24; // @[SRAM.scala 148:48:@61735.4]
  assign _T_913 = io_waddr == 6'h19; // @[SRAM.scala 148:37:@61743.4]
  assign _T_914 = io_wen & _T_913; // @[SRAM.scala 148:25:@61744.4]
  assign _T_915 = io_banks_25_wdata_valid | _T_914; // @[SRAM.scala 148:15:@61745.4]
  assign _T_916 = io_banks_25_wdata_valid ? io_banks_25_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61747.6]
  assign _GEN_25 = _T_915 ? _T_916 : regs_25; // @[SRAM.scala 148:48:@61746.4]
  assign _T_922 = io_waddr == 6'h1a; // @[SRAM.scala 148:37:@61754.4]
  assign _T_923 = io_wen & _T_922; // @[SRAM.scala 148:25:@61755.4]
  assign _T_924 = io_banks_26_wdata_valid | _T_923; // @[SRAM.scala 148:15:@61756.4]
  assign _T_925 = io_banks_26_wdata_valid ? io_banks_26_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61758.6]
  assign _GEN_26 = _T_924 ? _T_925 : regs_26; // @[SRAM.scala 148:48:@61757.4]
  assign _T_931 = io_waddr == 6'h1b; // @[SRAM.scala 148:37:@61765.4]
  assign _T_932 = io_wen & _T_931; // @[SRAM.scala 148:25:@61766.4]
  assign _T_933 = io_banks_27_wdata_valid | _T_932; // @[SRAM.scala 148:15:@61767.4]
  assign _T_934 = io_banks_27_wdata_valid ? io_banks_27_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61769.6]
  assign _GEN_27 = _T_933 ? _T_934 : regs_27; // @[SRAM.scala 148:48:@61768.4]
  assign _T_940 = io_waddr == 6'h1c; // @[SRAM.scala 148:37:@61776.4]
  assign _T_941 = io_wen & _T_940; // @[SRAM.scala 148:25:@61777.4]
  assign _T_942 = io_banks_28_wdata_valid | _T_941; // @[SRAM.scala 148:15:@61778.4]
  assign _T_943 = io_banks_28_wdata_valid ? io_banks_28_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61780.6]
  assign _GEN_28 = _T_942 ? _T_943 : regs_28; // @[SRAM.scala 148:48:@61779.4]
  assign _T_949 = io_waddr == 6'h1d; // @[SRAM.scala 148:37:@61787.4]
  assign _T_950 = io_wen & _T_949; // @[SRAM.scala 148:25:@61788.4]
  assign _T_951 = io_banks_29_wdata_valid | _T_950; // @[SRAM.scala 148:15:@61789.4]
  assign _T_952 = io_banks_29_wdata_valid ? io_banks_29_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61791.6]
  assign _GEN_29 = _T_951 ? _T_952 : regs_29; // @[SRAM.scala 148:48:@61790.4]
  assign _T_958 = io_waddr == 6'h1e; // @[SRAM.scala 148:37:@61798.4]
  assign _T_959 = io_wen & _T_958; // @[SRAM.scala 148:25:@61799.4]
  assign _T_960 = io_banks_30_wdata_valid | _T_959; // @[SRAM.scala 148:15:@61800.4]
  assign _T_961 = io_banks_30_wdata_valid ? io_banks_30_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61802.6]
  assign _GEN_30 = _T_960 ? _T_961 : regs_30; // @[SRAM.scala 148:48:@61801.4]
  assign _T_967 = io_waddr == 6'h1f; // @[SRAM.scala 148:37:@61809.4]
  assign _T_968 = io_wen & _T_967; // @[SRAM.scala 148:25:@61810.4]
  assign _T_969 = io_banks_31_wdata_valid | _T_968; // @[SRAM.scala 148:15:@61811.4]
  assign _T_970 = io_banks_31_wdata_valid ? io_banks_31_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61813.6]
  assign _GEN_31 = _T_969 ? _T_970 : regs_31; // @[SRAM.scala 148:48:@61812.4]
  assign _T_976 = io_waddr == 6'h20; // @[SRAM.scala 148:37:@61820.4]
  assign _T_977 = io_wen & _T_976; // @[SRAM.scala 148:25:@61821.4]
  assign _T_978 = io_banks_32_wdata_valid | _T_977; // @[SRAM.scala 148:15:@61822.4]
  assign _T_979 = io_banks_32_wdata_valid ? io_banks_32_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61824.6]
  assign _GEN_32 = _T_978 ? _T_979 : regs_32; // @[SRAM.scala 148:48:@61823.4]
  assign _T_985 = io_waddr == 6'h21; // @[SRAM.scala 148:37:@61831.4]
  assign _T_986 = io_wen & _T_985; // @[SRAM.scala 148:25:@61832.4]
  assign _T_987 = io_banks_33_wdata_valid | _T_986; // @[SRAM.scala 148:15:@61833.4]
  assign _T_988 = io_banks_33_wdata_valid ? io_banks_33_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61835.6]
  assign _GEN_33 = _T_987 ? _T_988 : regs_33; // @[SRAM.scala 148:48:@61834.4]
  assign _T_994 = io_waddr == 6'h22; // @[SRAM.scala 148:37:@61842.4]
  assign _T_995 = io_wen & _T_994; // @[SRAM.scala 148:25:@61843.4]
  assign _T_996 = io_banks_34_wdata_valid | _T_995; // @[SRAM.scala 148:15:@61844.4]
  assign _T_997 = io_banks_34_wdata_valid ? io_banks_34_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61846.6]
  assign _GEN_34 = _T_996 ? _T_997 : regs_34; // @[SRAM.scala 148:48:@61845.4]
  assign _T_1003 = io_waddr == 6'h23; // @[SRAM.scala 148:37:@61853.4]
  assign _T_1004 = io_wen & _T_1003; // @[SRAM.scala 148:25:@61854.4]
  assign _T_1005 = io_banks_35_wdata_valid | _T_1004; // @[SRAM.scala 148:15:@61855.4]
  assign _T_1006 = io_banks_35_wdata_valid ? io_banks_35_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61857.6]
  assign _GEN_35 = _T_1005 ? _T_1006 : regs_35; // @[SRAM.scala 148:48:@61856.4]
  assign _T_1012 = io_waddr == 6'h24; // @[SRAM.scala 148:37:@61864.4]
  assign _T_1013 = io_wen & _T_1012; // @[SRAM.scala 148:25:@61865.4]
  assign _T_1014 = io_banks_36_wdata_valid | _T_1013; // @[SRAM.scala 148:15:@61866.4]
  assign _T_1015 = io_banks_36_wdata_valid ? io_banks_36_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61868.6]
  assign _GEN_36 = _T_1014 ? _T_1015 : regs_36; // @[SRAM.scala 148:48:@61867.4]
  assign _T_1021 = io_waddr == 6'h25; // @[SRAM.scala 148:37:@61875.4]
  assign _T_1022 = io_wen & _T_1021; // @[SRAM.scala 148:25:@61876.4]
  assign _T_1023 = io_banks_37_wdata_valid | _T_1022; // @[SRAM.scala 148:15:@61877.4]
  assign _T_1024 = io_banks_37_wdata_valid ? io_banks_37_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61879.6]
  assign _GEN_37 = _T_1023 ? _T_1024 : regs_37; // @[SRAM.scala 148:48:@61878.4]
  assign _T_1030 = io_waddr == 6'h26; // @[SRAM.scala 148:37:@61886.4]
  assign _T_1031 = io_wen & _T_1030; // @[SRAM.scala 148:25:@61887.4]
  assign _T_1032 = io_banks_38_wdata_valid | _T_1031; // @[SRAM.scala 148:15:@61888.4]
  assign _T_1033 = io_banks_38_wdata_valid ? io_banks_38_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61890.6]
  assign _GEN_38 = _T_1032 ? _T_1033 : regs_38; // @[SRAM.scala 148:48:@61889.4]
  assign _T_1039 = io_waddr == 6'h27; // @[SRAM.scala 148:37:@61897.4]
  assign _T_1040 = io_wen & _T_1039; // @[SRAM.scala 148:25:@61898.4]
  assign _T_1041 = io_banks_39_wdata_valid | _T_1040; // @[SRAM.scala 148:15:@61899.4]
  assign _T_1042 = io_banks_39_wdata_valid ? io_banks_39_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61901.6]
  assign _GEN_39 = _T_1041 ? _T_1042 : regs_39; // @[SRAM.scala 148:48:@61900.4]
  assign _T_1048 = io_waddr == 6'h28; // @[SRAM.scala 148:37:@61908.4]
  assign _T_1049 = io_wen & _T_1048; // @[SRAM.scala 148:25:@61909.4]
  assign _T_1050 = io_banks_40_wdata_valid | _T_1049; // @[SRAM.scala 148:15:@61910.4]
  assign _T_1051 = io_banks_40_wdata_valid ? io_banks_40_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61912.6]
  assign _GEN_40 = _T_1050 ? _T_1051 : regs_40; // @[SRAM.scala 148:48:@61911.4]
  assign _T_1057 = io_waddr == 6'h29; // @[SRAM.scala 148:37:@61919.4]
  assign _T_1058 = io_wen & _T_1057; // @[SRAM.scala 148:25:@61920.4]
  assign _T_1059 = io_banks_41_wdata_valid | _T_1058; // @[SRAM.scala 148:15:@61921.4]
  assign _T_1060 = io_banks_41_wdata_valid ? io_banks_41_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61923.6]
  assign _GEN_41 = _T_1059 ? _T_1060 : regs_41; // @[SRAM.scala 148:48:@61922.4]
  assign _T_1066 = io_waddr == 6'h2a; // @[SRAM.scala 148:37:@61930.4]
  assign _T_1067 = io_wen & _T_1066; // @[SRAM.scala 148:25:@61931.4]
  assign _T_1068 = io_banks_42_wdata_valid | _T_1067; // @[SRAM.scala 148:15:@61932.4]
  assign _T_1069 = io_banks_42_wdata_valid ? io_banks_42_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61934.6]
  assign _GEN_42 = _T_1068 ? _T_1069 : regs_42; // @[SRAM.scala 148:48:@61933.4]
  assign _T_1075 = io_waddr == 6'h2b; // @[SRAM.scala 148:37:@61941.4]
  assign _T_1076 = io_wen & _T_1075; // @[SRAM.scala 148:25:@61942.4]
  assign _T_1077 = io_banks_43_wdata_valid | _T_1076; // @[SRAM.scala 148:15:@61943.4]
  assign _T_1078 = io_banks_43_wdata_valid ? io_banks_43_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61945.6]
  assign _GEN_43 = _T_1077 ? _T_1078 : regs_43; // @[SRAM.scala 148:48:@61944.4]
  assign _T_1084 = io_waddr == 6'h2c; // @[SRAM.scala 148:37:@61952.4]
  assign _T_1085 = io_wen & _T_1084; // @[SRAM.scala 148:25:@61953.4]
  assign _T_1086 = io_banks_44_wdata_valid | _T_1085; // @[SRAM.scala 148:15:@61954.4]
  assign _T_1087 = io_banks_44_wdata_valid ? io_banks_44_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61956.6]
  assign _GEN_44 = _T_1086 ? _T_1087 : regs_44; // @[SRAM.scala 148:48:@61955.4]
  assign _T_1093 = io_waddr == 6'h2d; // @[SRAM.scala 148:37:@61963.4]
  assign _T_1094 = io_wen & _T_1093; // @[SRAM.scala 148:25:@61964.4]
  assign _T_1095 = io_banks_45_wdata_valid | _T_1094; // @[SRAM.scala 148:15:@61965.4]
  assign _T_1096 = io_banks_45_wdata_valid ? io_banks_45_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61967.6]
  assign _GEN_45 = _T_1095 ? _T_1096 : regs_45; // @[SRAM.scala 148:48:@61966.4]
  assign _T_1102 = io_waddr == 6'h2e; // @[SRAM.scala 148:37:@61974.4]
  assign _T_1103 = io_wen & _T_1102; // @[SRAM.scala 148:25:@61975.4]
  assign _T_1104 = io_banks_46_wdata_valid | _T_1103; // @[SRAM.scala 148:15:@61976.4]
  assign _T_1105 = io_banks_46_wdata_valid ? io_banks_46_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61978.6]
  assign _GEN_46 = _T_1104 ? _T_1105 : regs_46; // @[SRAM.scala 148:48:@61977.4]
  assign _T_1111 = io_waddr == 6'h2f; // @[SRAM.scala 148:37:@61985.4]
  assign _T_1112 = io_wen & _T_1111; // @[SRAM.scala 148:25:@61986.4]
  assign _T_1113 = io_banks_47_wdata_valid | _T_1112; // @[SRAM.scala 148:15:@61987.4]
  assign _T_1114 = io_banks_47_wdata_valid ? io_banks_47_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@61989.6]
  assign _GEN_47 = _T_1113 ? _T_1114 : regs_47; // @[SRAM.scala 148:48:@61988.4]
  assign _T_1120 = io_waddr == 6'h30; // @[SRAM.scala 148:37:@61996.4]
  assign _T_1121 = io_wen & _T_1120; // @[SRAM.scala 148:25:@61997.4]
  assign _T_1122 = io_banks_48_wdata_valid | _T_1121; // @[SRAM.scala 148:15:@61998.4]
  assign _T_1123 = io_banks_48_wdata_valid ? io_banks_48_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62000.6]
  assign _GEN_48 = _T_1122 ? _T_1123 : regs_48; // @[SRAM.scala 148:48:@61999.4]
  assign _T_1129 = io_waddr == 6'h31; // @[SRAM.scala 148:37:@62007.4]
  assign _T_1130 = io_wen & _T_1129; // @[SRAM.scala 148:25:@62008.4]
  assign _T_1131 = io_banks_49_wdata_valid | _T_1130; // @[SRAM.scala 148:15:@62009.4]
  assign _T_1132 = io_banks_49_wdata_valid ? io_banks_49_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62011.6]
  assign _GEN_49 = _T_1131 ? _T_1132 : regs_49; // @[SRAM.scala 148:48:@62010.4]
  assign _T_1138 = io_waddr == 6'h32; // @[SRAM.scala 148:37:@62018.4]
  assign _T_1139 = io_wen & _T_1138; // @[SRAM.scala 148:25:@62019.4]
  assign _T_1140 = io_banks_50_wdata_valid | _T_1139; // @[SRAM.scala 148:15:@62020.4]
  assign _T_1141 = io_banks_50_wdata_valid ? io_banks_50_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62022.6]
  assign _GEN_50 = _T_1140 ? _T_1141 : regs_50; // @[SRAM.scala 148:48:@62021.4]
  assign _T_1147 = io_waddr == 6'h33; // @[SRAM.scala 148:37:@62029.4]
  assign _T_1148 = io_wen & _T_1147; // @[SRAM.scala 148:25:@62030.4]
  assign _T_1149 = io_banks_51_wdata_valid | _T_1148; // @[SRAM.scala 148:15:@62031.4]
  assign _T_1150 = io_banks_51_wdata_valid ? io_banks_51_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62033.6]
  assign _GEN_51 = _T_1149 ? _T_1150 : regs_51; // @[SRAM.scala 148:48:@62032.4]
  assign _T_1156 = io_waddr == 6'h34; // @[SRAM.scala 148:37:@62040.4]
  assign _T_1157 = io_wen & _T_1156; // @[SRAM.scala 148:25:@62041.4]
  assign _T_1158 = io_banks_52_wdata_valid | _T_1157; // @[SRAM.scala 148:15:@62042.4]
  assign _T_1159 = io_banks_52_wdata_valid ? io_banks_52_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62044.6]
  assign _GEN_52 = _T_1158 ? _T_1159 : regs_52; // @[SRAM.scala 148:48:@62043.4]
  assign _T_1165 = io_waddr == 6'h35; // @[SRAM.scala 148:37:@62051.4]
  assign _T_1166 = io_wen & _T_1165; // @[SRAM.scala 148:25:@62052.4]
  assign _T_1167 = io_banks_53_wdata_valid | _T_1166; // @[SRAM.scala 148:15:@62053.4]
  assign _T_1168 = io_banks_53_wdata_valid ? io_banks_53_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62055.6]
  assign _GEN_53 = _T_1167 ? _T_1168 : regs_53; // @[SRAM.scala 148:48:@62054.4]
  assign _T_1174 = io_waddr == 6'h36; // @[SRAM.scala 148:37:@62062.4]
  assign _T_1175 = io_wen & _T_1174; // @[SRAM.scala 148:25:@62063.4]
  assign _T_1176 = io_banks_54_wdata_valid | _T_1175; // @[SRAM.scala 148:15:@62064.4]
  assign _T_1177 = io_banks_54_wdata_valid ? io_banks_54_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62066.6]
  assign _GEN_54 = _T_1176 ? _T_1177 : regs_54; // @[SRAM.scala 148:48:@62065.4]
  assign _T_1183 = io_waddr == 6'h37; // @[SRAM.scala 148:37:@62073.4]
  assign _T_1184 = io_wen & _T_1183; // @[SRAM.scala 148:25:@62074.4]
  assign _T_1185 = io_banks_55_wdata_valid | _T_1184; // @[SRAM.scala 148:15:@62075.4]
  assign _T_1186 = io_banks_55_wdata_valid ? io_banks_55_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62077.6]
  assign _GEN_55 = _T_1185 ? _T_1186 : regs_55; // @[SRAM.scala 148:48:@62076.4]
  assign _T_1192 = io_waddr == 6'h38; // @[SRAM.scala 148:37:@62084.4]
  assign _T_1193 = io_wen & _T_1192; // @[SRAM.scala 148:25:@62085.4]
  assign _T_1194 = io_banks_56_wdata_valid | _T_1193; // @[SRAM.scala 148:15:@62086.4]
  assign _T_1195 = io_banks_56_wdata_valid ? io_banks_56_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62088.6]
  assign _GEN_56 = _T_1194 ? _T_1195 : regs_56; // @[SRAM.scala 148:48:@62087.4]
  assign _T_1201 = io_waddr == 6'h39; // @[SRAM.scala 148:37:@62095.4]
  assign _T_1202 = io_wen & _T_1201; // @[SRAM.scala 148:25:@62096.4]
  assign _T_1203 = io_banks_57_wdata_valid | _T_1202; // @[SRAM.scala 148:15:@62097.4]
  assign _T_1204 = io_banks_57_wdata_valid ? io_banks_57_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62099.6]
  assign _GEN_57 = _T_1203 ? _T_1204 : regs_57; // @[SRAM.scala 148:48:@62098.4]
  assign _T_1210 = io_waddr == 6'h3a; // @[SRAM.scala 148:37:@62106.4]
  assign _T_1211 = io_wen & _T_1210; // @[SRAM.scala 148:25:@62107.4]
  assign _T_1212 = io_banks_58_wdata_valid | _T_1211; // @[SRAM.scala 148:15:@62108.4]
  assign _T_1213 = io_banks_58_wdata_valid ? io_banks_58_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62110.6]
  assign _GEN_58 = _T_1212 ? _T_1213 : regs_58; // @[SRAM.scala 148:48:@62109.4]
  assign _T_1219 = io_waddr == 6'h3b; // @[SRAM.scala 148:37:@62117.4]
  assign _T_1220 = io_wen & _T_1219; // @[SRAM.scala 148:25:@62118.4]
  assign _T_1221 = io_banks_59_wdata_valid | _T_1220; // @[SRAM.scala 148:15:@62119.4]
  assign _T_1222 = io_banks_59_wdata_valid ? io_banks_59_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62121.6]
  assign _GEN_59 = _T_1221 ? _T_1222 : regs_59; // @[SRAM.scala 148:48:@62120.4]
  assign _T_1228 = io_waddr == 6'h3c; // @[SRAM.scala 148:37:@62128.4]
  assign _T_1229 = io_wen & _T_1228; // @[SRAM.scala 148:25:@62129.4]
  assign _T_1230 = io_banks_60_wdata_valid | _T_1229; // @[SRAM.scala 148:15:@62130.4]
  assign _T_1231 = io_banks_60_wdata_valid ? io_banks_60_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62132.6]
  assign _GEN_60 = _T_1230 ? _T_1231 : regs_60; // @[SRAM.scala 148:48:@62131.4]
  assign _T_1237 = io_waddr == 6'h3d; // @[SRAM.scala 148:37:@62139.4]
  assign _T_1238 = io_wen & _T_1237; // @[SRAM.scala 148:25:@62140.4]
  assign _T_1239 = io_banks_61_wdata_valid | _T_1238; // @[SRAM.scala 148:15:@62141.4]
  assign _T_1240 = io_banks_61_wdata_valid ? io_banks_61_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62143.6]
  assign _GEN_61 = _T_1239 ? _T_1240 : regs_61; // @[SRAM.scala 148:48:@62142.4]
  assign _T_1246 = io_waddr == 6'h3e; // @[SRAM.scala 148:37:@62150.4]
  assign _T_1247 = io_wen & _T_1246; // @[SRAM.scala 148:25:@62151.4]
  assign _T_1248 = io_banks_62_wdata_valid | _T_1247; // @[SRAM.scala 148:15:@62152.4]
  assign _T_1249 = io_banks_62_wdata_valid ? io_banks_62_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62154.6]
  assign _GEN_62 = _T_1248 ? _T_1249 : regs_62; // @[SRAM.scala 148:48:@62153.4]
  assign _T_1255 = io_waddr == 6'h3f; // @[SRAM.scala 148:37:@62161.4]
  assign _T_1256 = io_wen & _T_1255; // @[SRAM.scala 148:25:@62162.4]
  assign _T_1257 = io_banks_63_wdata_valid | _T_1256; // @[SRAM.scala 148:15:@62163.4]
  assign _T_1258 = io_banks_63_wdata_valid ? io_banks_63_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@62165.6]
  assign _GEN_63 = _T_1257 ? _T_1258 : regs_63; // @[SRAM.scala 148:48:@62164.4]
  assign _GEN_65 = 6'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_66 = 6'h2 == io_raddr ? regs_2 : _GEN_65; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_67 = 6'h3 == io_raddr ? regs_3 : _GEN_66; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_68 = 6'h4 == io_raddr ? regs_4 : _GEN_67; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_69 = 6'h5 == io_raddr ? regs_5 : _GEN_68; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_70 = 6'h6 == io_raddr ? regs_6 : _GEN_69; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_71 = 6'h7 == io_raddr ? regs_7 : _GEN_70; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_72 = 6'h8 == io_raddr ? regs_8 : _GEN_71; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_73 = 6'h9 == io_raddr ? regs_9 : _GEN_72; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_74 = 6'ha == io_raddr ? regs_10 : _GEN_73; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_75 = 6'hb == io_raddr ? regs_11 : _GEN_74; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_76 = 6'hc == io_raddr ? regs_12 : _GEN_75; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_77 = 6'hd == io_raddr ? regs_13 : _GEN_76; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_78 = 6'he == io_raddr ? regs_14 : _GEN_77; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_79 = 6'hf == io_raddr ? regs_15 : _GEN_78; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_80 = 6'h10 == io_raddr ? regs_16 : _GEN_79; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_81 = 6'h11 == io_raddr ? regs_17 : _GEN_80; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_82 = 6'h12 == io_raddr ? regs_18 : _GEN_81; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_83 = 6'h13 == io_raddr ? regs_19 : _GEN_82; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_84 = 6'h14 == io_raddr ? regs_20 : _GEN_83; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_85 = 6'h15 == io_raddr ? regs_21 : _GEN_84; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_86 = 6'h16 == io_raddr ? regs_22 : _GEN_85; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_87 = 6'h17 == io_raddr ? regs_23 : _GEN_86; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_88 = 6'h18 == io_raddr ? regs_24 : _GEN_87; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_89 = 6'h19 == io_raddr ? regs_25 : _GEN_88; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_90 = 6'h1a == io_raddr ? regs_26 : _GEN_89; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_91 = 6'h1b == io_raddr ? regs_27 : _GEN_90; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_92 = 6'h1c == io_raddr ? regs_28 : _GEN_91; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_93 = 6'h1d == io_raddr ? regs_29 : _GEN_92; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_94 = 6'h1e == io_raddr ? regs_30 : _GEN_93; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_95 = 6'h1f == io_raddr ? regs_31 : _GEN_94; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_96 = 6'h20 == io_raddr ? regs_32 : _GEN_95; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_97 = 6'h21 == io_raddr ? regs_33 : _GEN_96; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_98 = 6'h22 == io_raddr ? regs_34 : _GEN_97; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_99 = 6'h23 == io_raddr ? regs_35 : _GEN_98; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_100 = 6'h24 == io_raddr ? regs_36 : _GEN_99; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_101 = 6'h25 == io_raddr ? regs_37 : _GEN_100; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_102 = 6'h26 == io_raddr ? regs_38 : _GEN_101; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_103 = 6'h27 == io_raddr ? regs_39 : _GEN_102; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_104 = 6'h28 == io_raddr ? regs_40 : _GEN_103; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_105 = 6'h29 == io_raddr ? regs_41 : _GEN_104; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_106 = 6'h2a == io_raddr ? regs_42 : _GEN_105; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_107 = 6'h2b == io_raddr ? regs_43 : _GEN_106; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_108 = 6'h2c == io_raddr ? regs_44 : _GEN_107; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_109 = 6'h2d == io_raddr ? regs_45 : _GEN_108; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_110 = 6'h2e == io_raddr ? regs_46 : _GEN_109; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_111 = 6'h2f == io_raddr ? regs_47 : _GEN_110; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_112 = 6'h30 == io_raddr ? regs_48 : _GEN_111; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_113 = 6'h31 == io_raddr ? regs_49 : _GEN_112; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_114 = 6'h32 == io_raddr ? regs_50 : _GEN_113; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_115 = 6'h33 == io_raddr ? regs_51 : _GEN_114; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_116 = 6'h34 == io_raddr ? regs_52 : _GEN_115; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_117 = 6'h35 == io_raddr ? regs_53 : _GEN_116; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_118 = 6'h36 == io_raddr ? regs_54 : _GEN_117; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_119 = 6'h37 == io_raddr ? regs_55 : _GEN_118; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_120 = 6'h38 == io_raddr ? regs_56 : _GEN_119; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_121 = 6'h39 == io_raddr ? regs_57 : _GEN_120; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_122 = 6'h3a == io_raddr ? regs_58 : _GEN_121; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_123 = 6'h3b == io_raddr ? regs_59 : _GEN_122; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_124 = 6'h3c == io_raddr ? regs_60 : _GEN_123; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_125 = 6'h3d == io_raddr ? regs_61 : _GEN_124; // @[SRAM.scala 155:12:@62234.4]
  assign _GEN_126 = 6'h3e == io_raddr ? regs_62 : _GEN_125; // @[SRAM.scala 155:12:@62234.4]
  assign io_rdata = 6'h3f == io_raddr ? regs_63 : _GEN_126; // @[SRAM.scala 155:12:@62234.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_690) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_699) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_708) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_717) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_4 <= 1'h0;
    end else begin
      if (_T_726) begin
        if (io_banks_4_wdata_valid) begin
          regs_4 <= io_banks_4_wdata_bits;
        end else begin
          regs_4 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_5 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (io_banks_5_wdata_valid) begin
          regs_5 <= io_banks_5_wdata_bits;
        end else begin
          regs_5 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_6 <= 1'h0;
    end else begin
      if (_T_744) begin
        if (io_banks_6_wdata_valid) begin
          regs_6 <= io_banks_6_wdata_bits;
        end else begin
          regs_6 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_7 <= 1'h0;
    end else begin
      if (_T_753) begin
        if (io_banks_7_wdata_valid) begin
          regs_7 <= io_banks_7_wdata_bits;
        end else begin
          regs_7 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_8 <= 1'h0;
    end else begin
      if (_T_762) begin
        if (io_banks_8_wdata_valid) begin
          regs_8 <= io_banks_8_wdata_bits;
        end else begin
          regs_8 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_9 <= 1'h0;
    end else begin
      if (_T_771) begin
        if (io_banks_9_wdata_valid) begin
          regs_9 <= io_banks_9_wdata_bits;
        end else begin
          regs_9 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_10 <= 1'h0;
    end else begin
      if (_T_780) begin
        if (io_banks_10_wdata_valid) begin
          regs_10 <= io_banks_10_wdata_bits;
        end else begin
          regs_10 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_11 <= 1'h0;
    end else begin
      if (_T_789) begin
        if (io_banks_11_wdata_valid) begin
          regs_11 <= io_banks_11_wdata_bits;
        end else begin
          regs_11 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_12 <= 1'h0;
    end else begin
      if (_T_798) begin
        if (io_banks_12_wdata_valid) begin
          regs_12 <= io_banks_12_wdata_bits;
        end else begin
          regs_12 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_13 <= 1'h0;
    end else begin
      if (_T_807) begin
        if (io_banks_13_wdata_valid) begin
          regs_13 <= io_banks_13_wdata_bits;
        end else begin
          regs_13 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_14 <= 1'h0;
    end else begin
      if (_T_816) begin
        if (io_banks_14_wdata_valid) begin
          regs_14 <= io_banks_14_wdata_bits;
        end else begin
          regs_14 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_15 <= 1'h0;
    end else begin
      if (_T_825) begin
        if (io_banks_15_wdata_valid) begin
          regs_15 <= io_banks_15_wdata_bits;
        end else begin
          regs_15 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_16 <= 1'h0;
    end else begin
      if (_T_834) begin
        if (io_banks_16_wdata_valid) begin
          regs_16 <= io_banks_16_wdata_bits;
        end else begin
          regs_16 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_17 <= 1'h0;
    end else begin
      if (_T_843) begin
        if (io_banks_17_wdata_valid) begin
          regs_17 <= io_banks_17_wdata_bits;
        end else begin
          regs_17 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_18 <= 1'h0;
    end else begin
      if (_T_852) begin
        if (io_banks_18_wdata_valid) begin
          regs_18 <= io_banks_18_wdata_bits;
        end else begin
          regs_18 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_19 <= 1'h0;
    end else begin
      if (_T_861) begin
        if (io_banks_19_wdata_valid) begin
          regs_19 <= io_banks_19_wdata_bits;
        end else begin
          regs_19 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_20 <= 1'h0;
    end else begin
      if (_T_870) begin
        if (io_banks_20_wdata_valid) begin
          regs_20 <= io_banks_20_wdata_bits;
        end else begin
          regs_20 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_21 <= 1'h0;
    end else begin
      if (_T_879) begin
        if (io_banks_21_wdata_valid) begin
          regs_21 <= io_banks_21_wdata_bits;
        end else begin
          regs_21 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_22 <= 1'h0;
    end else begin
      if (_T_888) begin
        if (io_banks_22_wdata_valid) begin
          regs_22 <= io_banks_22_wdata_bits;
        end else begin
          regs_22 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_23 <= 1'h0;
    end else begin
      if (_T_897) begin
        if (io_banks_23_wdata_valid) begin
          regs_23 <= io_banks_23_wdata_bits;
        end else begin
          regs_23 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_24 <= 1'h0;
    end else begin
      if (_T_906) begin
        if (io_banks_24_wdata_valid) begin
          regs_24 <= io_banks_24_wdata_bits;
        end else begin
          regs_24 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_25 <= 1'h0;
    end else begin
      if (_T_915) begin
        if (io_banks_25_wdata_valid) begin
          regs_25 <= io_banks_25_wdata_bits;
        end else begin
          regs_25 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_26 <= 1'h0;
    end else begin
      if (_T_924) begin
        if (io_banks_26_wdata_valid) begin
          regs_26 <= io_banks_26_wdata_bits;
        end else begin
          regs_26 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_27 <= 1'h0;
    end else begin
      if (_T_933) begin
        if (io_banks_27_wdata_valid) begin
          regs_27 <= io_banks_27_wdata_bits;
        end else begin
          regs_27 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_28 <= 1'h0;
    end else begin
      if (_T_942) begin
        if (io_banks_28_wdata_valid) begin
          regs_28 <= io_banks_28_wdata_bits;
        end else begin
          regs_28 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_29 <= 1'h0;
    end else begin
      if (_T_951) begin
        if (io_banks_29_wdata_valid) begin
          regs_29 <= io_banks_29_wdata_bits;
        end else begin
          regs_29 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_30 <= 1'h0;
    end else begin
      if (_T_960) begin
        if (io_banks_30_wdata_valid) begin
          regs_30 <= io_banks_30_wdata_bits;
        end else begin
          regs_30 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_31 <= 1'h0;
    end else begin
      if (_T_969) begin
        if (io_banks_31_wdata_valid) begin
          regs_31 <= io_banks_31_wdata_bits;
        end else begin
          regs_31 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_32 <= 1'h0;
    end else begin
      if (_T_978) begin
        if (io_banks_32_wdata_valid) begin
          regs_32 <= io_banks_32_wdata_bits;
        end else begin
          regs_32 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_33 <= 1'h0;
    end else begin
      if (_T_987) begin
        if (io_banks_33_wdata_valid) begin
          regs_33 <= io_banks_33_wdata_bits;
        end else begin
          regs_33 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_34 <= 1'h0;
    end else begin
      if (_T_996) begin
        if (io_banks_34_wdata_valid) begin
          regs_34 <= io_banks_34_wdata_bits;
        end else begin
          regs_34 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_35 <= 1'h0;
    end else begin
      if (_T_1005) begin
        if (io_banks_35_wdata_valid) begin
          regs_35 <= io_banks_35_wdata_bits;
        end else begin
          regs_35 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_36 <= 1'h0;
    end else begin
      if (_T_1014) begin
        if (io_banks_36_wdata_valid) begin
          regs_36 <= io_banks_36_wdata_bits;
        end else begin
          regs_36 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_37 <= 1'h0;
    end else begin
      if (_T_1023) begin
        if (io_banks_37_wdata_valid) begin
          regs_37 <= io_banks_37_wdata_bits;
        end else begin
          regs_37 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_38 <= 1'h0;
    end else begin
      if (_T_1032) begin
        if (io_banks_38_wdata_valid) begin
          regs_38 <= io_banks_38_wdata_bits;
        end else begin
          regs_38 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_39 <= 1'h0;
    end else begin
      if (_T_1041) begin
        if (io_banks_39_wdata_valid) begin
          regs_39 <= io_banks_39_wdata_bits;
        end else begin
          regs_39 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_40 <= 1'h0;
    end else begin
      if (_T_1050) begin
        if (io_banks_40_wdata_valid) begin
          regs_40 <= io_banks_40_wdata_bits;
        end else begin
          regs_40 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_41 <= 1'h0;
    end else begin
      if (_T_1059) begin
        if (io_banks_41_wdata_valid) begin
          regs_41 <= io_banks_41_wdata_bits;
        end else begin
          regs_41 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_42 <= 1'h0;
    end else begin
      if (_T_1068) begin
        if (io_banks_42_wdata_valid) begin
          regs_42 <= io_banks_42_wdata_bits;
        end else begin
          regs_42 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_43 <= 1'h0;
    end else begin
      if (_T_1077) begin
        if (io_banks_43_wdata_valid) begin
          regs_43 <= io_banks_43_wdata_bits;
        end else begin
          regs_43 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_44 <= 1'h0;
    end else begin
      if (_T_1086) begin
        if (io_banks_44_wdata_valid) begin
          regs_44 <= io_banks_44_wdata_bits;
        end else begin
          regs_44 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_45 <= 1'h0;
    end else begin
      if (_T_1095) begin
        if (io_banks_45_wdata_valid) begin
          regs_45 <= io_banks_45_wdata_bits;
        end else begin
          regs_45 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_46 <= 1'h0;
    end else begin
      if (_T_1104) begin
        if (io_banks_46_wdata_valid) begin
          regs_46 <= io_banks_46_wdata_bits;
        end else begin
          regs_46 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_47 <= 1'h0;
    end else begin
      if (_T_1113) begin
        if (io_banks_47_wdata_valid) begin
          regs_47 <= io_banks_47_wdata_bits;
        end else begin
          regs_47 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_48 <= 1'h0;
    end else begin
      if (_T_1122) begin
        if (io_banks_48_wdata_valid) begin
          regs_48 <= io_banks_48_wdata_bits;
        end else begin
          regs_48 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_49 <= 1'h0;
    end else begin
      if (_T_1131) begin
        if (io_banks_49_wdata_valid) begin
          regs_49 <= io_banks_49_wdata_bits;
        end else begin
          regs_49 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_50 <= 1'h0;
    end else begin
      if (_T_1140) begin
        if (io_banks_50_wdata_valid) begin
          regs_50 <= io_banks_50_wdata_bits;
        end else begin
          regs_50 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_51 <= 1'h0;
    end else begin
      if (_T_1149) begin
        if (io_banks_51_wdata_valid) begin
          regs_51 <= io_banks_51_wdata_bits;
        end else begin
          regs_51 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_52 <= 1'h0;
    end else begin
      if (_T_1158) begin
        if (io_banks_52_wdata_valid) begin
          regs_52 <= io_banks_52_wdata_bits;
        end else begin
          regs_52 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_53 <= 1'h0;
    end else begin
      if (_T_1167) begin
        if (io_banks_53_wdata_valid) begin
          regs_53 <= io_banks_53_wdata_bits;
        end else begin
          regs_53 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_54 <= 1'h0;
    end else begin
      if (_T_1176) begin
        if (io_banks_54_wdata_valid) begin
          regs_54 <= io_banks_54_wdata_bits;
        end else begin
          regs_54 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_55 <= 1'h0;
    end else begin
      if (_T_1185) begin
        if (io_banks_55_wdata_valid) begin
          regs_55 <= io_banks_55_wdata_bits;
        end else begin
          regs_55 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_56 <= 1'h0;
    end else begin
      if (_T_1194) begin
        if (io_banks_56_wdata_valid) begin
          regs_56 <= io_banks_56_wdata_bits;
        end else begin
          regs_56 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_57 <= 1'h0;
    end else begin
      if (_T_1203) begin
        if (io_banks_57_wdata_valid) begin
          regs_57 <= io_banks_57_wdata_bits;
        end else begin
          regs_57 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_58 <= 1'h0;
    end else begin
      if (_T_1212) begin
        if (io_banks_58_wdata_valid) begin
          regs_58 <= io_banks_58_wdata_bits;
        end else begin
          regs_58 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_59 <= 1'h0;
    end else begin
      if (_T_1221) begin
        if (io_banks_59_wdata_valid) begin
          regs_59 <= io_banks_59_wdata_bits;
        end else begin
          regs_59 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_60 <= 1'h0;
    end else begin
      if (_T_1230) begin
        if (io_banks_60_wdata_valid) begin
          regs_60 <= io_banks_60_wdata_bits;
        end else begin
          regs_60 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_61 <= 1'h0;
    end else begin
      if (_T_1239) begin
        if (io_banks_61_wdata_valid) begin
          regs_61 <= io_banks_61_wdata_bits;
        end else begin
          regs_61 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_62 <= 1'h0;
    end else begin
      if (_T_1248) begin
        if (io_banks_62_wdata_valid) begin
          regs_62 <= io_banks_62_wdata_bits;
        end else begin
          regs_62 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_63 <= 1'h0;
    end else begin
      if (_T_1257) begin
        if (io_banks_63_wdata_valid) begin
          regs_63 <= io_banks_63_wdata_bits;
        end else begin
          regs_63 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_33( // @[:@62236.2]
  input   clock, // @[:@62237.4]
  input   reset, // @[:@62238.4]
  output  io_in_ready, // @[:@62239.4]
  input   io_in_valid, // @[:@62239.4]
  input   io_in_bits, // @[:@62239.4]
  input   io_out_ready, // @[:@62239.4]
  output  io_out_valid, // @[:@62239.4]
  output  io_out_bits, // @[:@62239.4]
  input   io_banks_0_wdata_valid, // @[:@62239.4]
  input   io_banks_0_wdata_bits, // @[:@62239.4]
  input   io_banks_1_wdata_valid, // @[:@62239.4]
  input   io_banks_1_wdata_bits, // @[:@62239.4]
  input   io_banks_2_wdata_valid, // @[:@62239.4]
  input   io_banks_2_wdata_bits, // @[:@62239.4]
  input   io_banks_3_wdata_valid, // @[:@62239.4]
  input   io_banks_3_wdata_bits, // @[:@62239.4]
  input   io_banks_4_wdata_valid, // @[:@62239.4]
  input   io_banks_4_wdata_bits, // @[:@62239.4]
  input   io_banks_5_wdata_valid, // @[:@62239.4]
  input   io_banks_5_wdata_bits, // @[:@62239.4]
  input   io_banks_6_wdata_valid, // @[:@62239.4]
  input   io_banks_6_wdata_bits, // @[:@62239.4]
  input   io_banks_7_wdata_valid, // @[:@62239.4]
  input   io_banks_7_wdata_bits, // @[:@62239.4]
  input   io_banks_8_wdata_valid, // @[:@62239.4]
  input   io_banks_8_wdata_bits, // @[:@62239.4]
  input   io_banks_9_wdata_valid, // @[:@62239.4]
  input   io_banks_9_wdata_bits, // @[:@62239.4]
  input   io_banks_10_wdata_valid, // @[:@62239.4]
  input   io_banks_10_wdata_bits, // @[:@62239.4]
  input   io_banks_11_wdata_valid, // @[:@62239.4]
  input   io_banks_11_wdata_bits, // @[:@62239.4]
  input   io_banks_12_wdata_valid, // @[:@62239.4]
  input   io_banks_12_wdata_bits, // @[:@62239.4]
  input   io_banks_13_wdata_valid, // @[:@62239.4]
  input   io_banks_13_wdata_bits, // @[:@62239.4]
  input   io_banks_14_wdata_valid, // @[:@62239.4]
  input   io_banks_14_wdata_bits, // @[:@62239.4]
  input   io_banks_15_wdata_valid, // @[:@62239.4]
  input   io_banks_15_wdata_bits, // @[:@62239.4]
  input   io_banks_16_wdata_valid, // @[:@62239.4]
  input   io_banks_16_wdata_bits, // @[:@62239.4]
  input   io_banks_17_wdata_valid, // @[:@62239.4]
  input   io_banks_17_wdata_bits, // @[:@62239.4]
  input   io_banks_18_wdata_valid, // @[:@62239.4]
  input   io_banks_18_wdata_bits, // @[:@62239.4]
  input   io_banks_19_wdata_valid, // @[:@62239.4]
  input   io_banks_19_wdata_bits, // @[:@62239.4]
  input   io_banks_20_wdata_valid, // @[:@62239.4]
  input   io_banks_20_wdata_bits, // @[:@62239.4]
  input   io_banks_21_wdata_valid, // @[:@62239.4]
  input   io_banks_21_wdata_bits, // @[:@62239.4]
  input   io_banks_22_wdata_valid, // @[:@62239.4]
  input   io_banks_22_wdata_bits, // @[:@62239.4]
  input   io_banks_23_wdata_valid, // @[:@62239.4]
  input   io_banks_23_wdata_bits, // @[:@62239.4]
  input   io_banks_24_wdata_valid, // @[:@62239.4]
  input   io_banks_24_wdata_bits, // @[:@62239.4]
  input   io_banks_25_wdata_valid, // @[:@62239.4]
  input   io_banks_25_wdata_bits, // @[:@62239.4]
  input   io_banks_26_wdata_valid, // @[:@62239.4]
  input   io_banks_26_wdata_bits, // @[:@62239.4]
  input   io_banks_27_wdata_valid, // @[:@62239.4]
  input   io_banks_27_wdata_bits, // @[:@62239.4]
  input   io_banks_28_wdata_valid, // @[:@62239.4]
  input   io_banks_28_wdata_bits, // @[:@62239.4]
  input   io_banks_29_wdata_valid, // @[:@62239.4]
  input   io_banks_29_wdata_bits, // @[:@62239.4]
  input   io_banks_30_wdata_valid, // @[:@62239.4]
  input   io_banks_30_wdata_bits, // @[:@62239.4]
  input   io_banks_31_wdata_valid, // @[:@62239.4]
  input   io_banks_31_wdata_bits, // @[:@62239.4]
  input   io_banks_32_wdata_valid, // @[:@62239.4]
  input   io_banks_32_wdata_bits, // @[:@62239.4]
  input   io_banks_33_wdata_valid, // @[:@62239.4]
  input   io_banks_33_wdata_bits, // @[:@62239.4]
  input   io_banks_34_wdata_valid, // @[:@62239.4]
  input   io_banks_34_wdata_bits, // @[:@62239.4]
  input   io_banks_35_wdata_valid, // @[:@62239.4]
  input   io_banks_35_wdata_bits, // @[:@62239.4]
  input   io_banks_36_wdata_valid, // @[:@62239.4]
  input   io_banks_36_wdata_bits, // @[:@62239.4]
  input   io_banks_37_wdata_valid, // @[:@62239.4]
  input   io_banks_37_wdata_bits, // @[:@62239.4]
  input   io_banks_38_wdata_valid, // @[:@62239.4]
  input   io_banks_38_wdata_bits, // @[:@62239.4]
  input   io_banks_39_wdata_valid, // @[:@62239.4]
  input   io_banks_39_wdata_bits, // @[:@62239.4]
  input   io_banks_40_wdata_valid, // @[:@62239.4]
  input   io_banks_40_wdata_bits, // @[:@62239.4]
  input   io_banks_41_wdata_valid, // @[:@62239.4]
  input   io_banks_41_wdata_bits, // @[:@62239.4]
  input   io_banks_42_wdata_valid, // @[:@62239.4]
  input   io_banks_42_wdata_bits, // @[:@62239.4]
  input   io_banks_43_wdata_valid, // @[:@62239.4]
  input   io_banks_43_wdata_bits, // @[:@62239.4]
  input   io_banks_44_wdata_valid, // @[:@62239.4]
  input   io_banks_44_wdata_bits, // @[:@62239.4]
  input   io_banks_45_wdata_valid, // @[:@62239.4]
  input   io_banks_45_wdata_bits, // @[:@62239.4]
  input   io_banks_46_wdata_valid, // @[:@62239.4]
  input   io_banks_46_wdata_bits, // @[:@62239.4]
  input   io_banks_47_wdata_valid, // @[:@62239.4]
  input   io_banks_47_wdata_bits, // @[:@62239.4]
  input   io_banks_48_wdata_valid, // @[:@62239.4]
  input   io_banks_48_wdata_bits, // @[:@62239.4]
  input   io_banks_49_wdata_valid, // @[:@62239.4]
  input   io_banks_49_wdata_bits, // @[:@62239.4]
  input   io_banks_50_wdata_valid, // @[:@62239.4]
  input   io_banks_50_wdata_bits, // @[:@62239.4]
  input   io_banks_51_wdata_valid, // @[:@62239.4]
  input   io_banks_51_wdata_bits, // @[:@62239.4]
  input   io_banks_52_wdata_valid, // @[:@62239.4]
  input   io_banks_52_wdata_bits, // @[:@62239.4]
  input   io_banks_53_wdata_valid, // @[:@62239.4]
  input   io_banks_53_wdata_bits, // @[:@62239.4]
  input   io_banks_54_wdata_valid, // @[:@62239.4]
  input   io_banks_54_wdata_bits, // @[:@62239.4]
  input   io_banks_55_wdata_valid, // @[:@62239.4]
  input   io_banks_55_wdata_bits, // @[:@62239.4]
  input   io_banks_56_wdata_valid, // @[:@62239.4]
  input   io_banks_56_wdata_bits, // @[:@62239.4]
  input   io_banks_57_wdata_valid, // @[:@62239.4]
  input   io_banks_57_wdata_bits, // @[:@62239.4]
  input   io_banks_58_wdata_valid, // @[:@62239.4]
  input   io_banks_58_wdata_bits, // @[:@62239.4]
  input   io_banks_59_wdata_valid, // @[:@62239.4]
  input   io_banks_59_wdata_bits, // @[:@62239.4]
  input   io_banks_60_wdata_valid, // @[:@62239.4]
  input   io_banks_60_wdata_bits, // @[:@62239.4]
  input   io_banks_61_wdata_valid, // @[:@62239.4]
  input   io_banks_61_wdata_bits, // @[:@62239.4]
  input   io_banks_62_wdata_valid, // @[:@62239.4]
  input   io_banks_62_wdata_bits, // @[:@62239.4]
  input   io_banks_63_wdata_valid, // @[:@62239.4]
  input   io_banks_63_wdata_bits // @[:@62239.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@62505.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@62505.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@62505.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@62505.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@62505.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@62515.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@62515.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@62515.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@62515.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@62515.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@62530.4]
  wire [5:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@62530.4]
  wire [5:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_4_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_4_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_5_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_5_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_6_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_6_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_7_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_7_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_8_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_8_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_9_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_9_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_10_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_10_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_11_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_11_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_12_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_12_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_13_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_13_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_14_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_14_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_15_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_15_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_16_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_16_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_17_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_17_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_18_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_18_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_19_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_19_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_20_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_20_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_21_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_21_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_22_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_22_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_23_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_23_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_24_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_24_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_25_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_25_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_26_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_26_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_27_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_27_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_28_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_28_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_29_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_29_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_30_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_30_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_31_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_31_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_32_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_32_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_33_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_33_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_34_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_34_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_35_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_35_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_36_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_36_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_37_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_37_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_38_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_38_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_39_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_39_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_40_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_40_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_41_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_41_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_42_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_42_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_43_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_43_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_44_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_44_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_45_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_45_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_46_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_46_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_47_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_47_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_48_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_48_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_49_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_49_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_50_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_50_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_51_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_51_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_52_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_52_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_53_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_53_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_54_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_54_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_55_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_55_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_56_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_56_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_57_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_57_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_58_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_58_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_59_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_59_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_60_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_60_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_61_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_61_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_62_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_62_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_63_wdata_valid; // @[FIFO.scala 49:19:@62530.4]
  wire  FFRAM_io_banks_63_wdata_bits; // @[FIFO.scala 49:19:@62530.4]
  wire  writeEn; // @[FIFO.scala 30:29:@62503.4]
  wire  readEn; // @[FIFO.scala 31:29:@62504.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@62525.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@62526.4]
  wire  _T_824; // @[FIFO.scala 45:27:@62527.4]
  wire  empty; // @[FIFO.scala 45:24:@62528.4]
  wire  full; // @[FIFO.scala 46:23:@62529.4]
  wire  _T_1657; // @[FIFO.scala 83:17:@63696.4]
  wire  _GEN_64; // @[FIFO.scala 83:29:@63697.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@62505.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@62515.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM_16 FFRAM ( // @[FIFO.scala 49:19:@62530.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(FFRAM_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(FFRAM_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(FFRAM_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(FFRAM_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(FFRAM_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(FFRAM_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(FFRAM_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(FFRAM_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(FFRAM_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(FFRAM_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(FFRAM_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(FFRAM_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(FFRAM_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(FFRAM_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(FFRAM_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(FFRAM_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(FFRAM_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(FFRAM_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(FFRAM_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(FFRAM_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(FFRAM_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(FFRAM_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(FFRAM_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(FFRAM_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(FFRAM_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(FFRAM_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(FFRAM_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(FFRAM_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(FFRAM_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(FFRAM_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(FFRAM_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(FFRAM_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(FFRAM_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(FFRAM_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(FFRAM_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(FFRAM_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(FFRAM_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(FFRAM_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(FFRAM_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(FFRAM_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(FFRAM_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(FFRAM_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(FFRAM_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(FFRAM_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(FFRAM_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(FFRAM_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(FFRAM_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(FFRAM_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(FFRAM_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(FFRAM_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(FFRAM_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(FFRAM_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(FFRAM_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(FFRAM_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(FFRAM_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(FFRAM_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(FFRAM_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(FFRAM_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(FFRAM_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(FFRAM_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(FFRAM_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(FFRAM_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(FFRAM_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(FFRAM_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(FFRAM_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(FFRAM_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(FFRAM_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(FFRAM_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(FFRAM_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(FFRAM_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(FFRAM_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(FFRAM_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(FFRAM_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(FFRAM_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(FFRAM_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(FFRAM_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(FFRAM_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(FFRAM_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(FFRAM_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(FFRAM_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(FFRAM_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(FFRAM_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(FFRAM_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(FFRAM_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(FFRAM_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(FFRAM_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(FFRAM_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(FFRAM_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(FFRAM_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(FFRAM_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(FFRAM_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(FFRAM_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(FFRAM_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(FFRAM_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(FFRAM_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(FFRAM_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(FFRAM_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(FFRAM_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(FFRAM_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(FFRAM_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(FFRAM_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(FFRAM_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(FFRAM_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(FFRAM_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(FFRAM_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(FFRAM_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(FFRAM_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(FFRAM_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(FFRAM_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(FFRAM_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(FFRAM_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(FFRAM_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(FFRAM_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(FFRAM_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(FFRAM_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(FFRAM_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(FFRAM_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(FFRAM_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(FFRAM_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(FFRAM_io_banks_63_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@62503.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@62504.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@62526.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@62527.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@62528.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@62529.4]
  assign _T_1657 = writeEn != readEn; // @[FIFO.scala 83:17:@63696.4]
  assign _GEN_64 = _T_1657 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@63697.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@63703.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@63701.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@62735.4]
  assign enqCounter_clock = clock; // @[:@62506.4]
  assign enqCounter_reset = reset; // @[:@62507.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@62513.4]
  assign deqCounter_clock = clock; // @[:@62516.4]
  assign deqCounter_reset = reset; // @[:@62517.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@62523.4]
  assign FFRAM_clock = clock; // @[:@62531.4]
  assign FFRAM_reset = reset; // @[:@62532.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@62731.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@62732.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@62733.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@62734.4]
  assign FFRAM_io_banks_0_wdata_valid = io_banks_0_wdata_valid; // @[FIFO.scala 59:15:@62737.4]
  assign FFRAM_io_banks_0_wdata_bits = io_banks_0_wdata_bits; // @[FIFO.scala 59:15:@62736.4]
  assign FFRAM_io_banks_1_wdata_valid = io_banks_1_wdata_valid; // @[FIFO.scala 59:15:@62740.4]
  assign FFRAM_io_banks_1_wdata_bits = io_banks_1_wdata_bits; // @[FIFO.scala 59:15:@62739.4]
  assign FFRAM_io_banks_2_wdata_valid = io_banks_2_wdata_valid; // @[FIFO.scala 59:15:@62743.4]
  assign FFRAM_io_banks_2_wdata_bits = io_banks_2_wdata_bits; // @[FIFO.scala 59:15:@62742.4]
  assign FFRAM_io_banks_3_wdata_valid = io_banks_3_wdata_valid; // @[FIFO.scala 59:15:@62746.4]
  assign FFRAM_io_banks_3_wdata_bits = io_banks_3_wdata_bits; // @[FIFO.scala 59:15:@62745.4]
  assign FFRAM_io_banks_4_wdata_valid = io_banks_4_wdata_valid; // @[FIFO.scala 59:15:@62749.4]
  assign FFRAM_io_banks_4_wdata_bits = io_banks_4_wdata_bits; // @[FIFO.scala 59:15:@62748.4]
  assign FFRAM_io_banks_5_wdata_valid = io_banks_5_wdata_valid; // @[FIFO.scala 59:15:@62752.4]
  assign FFRAM_io_banks_5_wdata_bits = io_banks_5_wdata_bits; // @[FIFO.scala 59:15:@62751.4]
  assign FFRAM_io_banks_6_wdata_valid = io_banks_6_wdata_valid; // @[FIFO.scala 59:15:@62755.4]
  assign FFRAM_io_banks_6_wdata_bits = io_banks_6_wdata_bits; // @[FIFO.scala 59:15:@62754.4]
  assign FFRAM_io_banks_7_wdata_valid = io_banks_7_wdata_valid; // @[FIFO.scala 59:15:@62758.4]
  assign FFRAM_io_banks_7_wdata_bits = io_banks_7_wdata_bits; // @[FIFO.scala 59:15:@62757.4]
  assign FFRAM_io_banks_8_wdata_valid = io_banks_8_wdata_valid; // @[FIFO.scala 59:15:@62761.4]
  assign FFRAM_io_banks_8_wdata_bits = io_banks_8_wdata_bits; // @[FIFO.scala 59:15:@62760.4]
  assign FFRAM_io_banks_9_wdata_valid = io_banks_9_wdata_valid; // @[FIFO.scala 59:15:@62764.4]
  assign FFRAM_io_banks_9_wdata_bits = io_banks_9_wdata_bits; // @[FIFO.scala 59:15:@62763.4]
  assign FFRAM_io_banks_10_wdata_valid = io_banks_10_wdata_valid; // @[FIFO.scala 59:15:@62767.4]
  assign FFRAM_io_banks_10_wdata_bits = io_banks_10_wdata_bits; // @[FIFO.scala 59:15:@62766.4]
  assign FFRAM_io_banks_11_wdata_valid = io_banks_11_wdata_valid; // @[FIFO.scala 59:15:@62770.4]
  assign FFRAM_io_banks_11_wdata_bits = io_banks_11_wdata_bits; // @[FIFO.scala 59:15:@62769.4]
  assign FFRAM_io_banks_12_wdata_valid = io_banks_12_wdata_valid; // @[FIFO.scala 59:15:@62773.4]
  assign FFRAM_io_banks_12_wdata_bits = io_banks_12_wdata_bits; // @[FIFO.scala 59:15:@62772.4]
  assign FFRAM_io_banks_13_wdata_valid = io_banks_13_wdata_valid; // @[FIFO.scala 59:15:@62776.4]
  assign FFRAM_io_banks_13_wdata_bits = io_banks_13_wdata_bits; // @[FIFO.scala 59:15:@62775.4]
  assign FFRAM_io_banks_14_wdata_valid = io_banks_14_wdata_valid; // @[FIFO.scala 59:15:@62779.4]
  assign FFRAM_io_banks_14_wdata_bits = io_banks_14_wdata_bits; // @[FIFO.scala 59:15:@62778.4]
  assign FFRAM_io_banks_15_wdata_valid = io_banks_15_wdata_valid; // @[FIFO.scala 59:15:@62782.4]
  assign FFRAM_io_banks_15_wdata_bits = io_banks_15_wdata_bits; // @[FIFO.scala 59:15:@62781.4]
  assign FFRAM_io_banks_16_wdata_valid = io_banks_16_wdata_valid; // @[FIFO.scala 59:15:@62785.4]
  assign FFRAM_io_banks_16_wdata_bits = io_banks_16_wdata_bits; // @[FIFO.scala 59:15:@62784.4]
  assign FFRAM_io_banks_17_wdata_valid = io_banks_17_wdata_valid; // @[FIFO.scala 59:15:@62788.4]
  assign FFRAM_io_banks_17_wdata_bits = io_banks_17_wdata_bits; // @[FIFO.scala 59:15:@62787.4]
  assign FFRAM_io_banks_18_wdata_valid = io_banks_18_wdata_valid; // @[FIFO.scala 59:15:@62791.4]
  assign FFRAM_io_banks_18_wdata_bits = io_banks_18_wdata_bits; // @[FIFO.scala 59:15:@62790.4]
  assign FFRAM_io_banks_19_wdata_valid = io_banks_19_wdata_valid; // @[FIFO.scala 59:15:@62794.4]
  assign FFRAM_io_banks_19_wdata_bits = io_banks_19_wdata_bits; // @[FIFO.scala 59:15:@62793.4]
  assign FFRAM_io_banks_20_wdata_valid = io_banks_20_wdata_valid; // @[FIFO.scala 59:15:@62797.4]
  assign FFRAM_io_banks_20_wdata_bits = io_banks_20_wdata_bits; // @[FIFO.scala 59:15:@62796.4]
  assign FFRAM_io_banks_21_wdata_valid = io_banks_21_wdata_valid; // @[FIFO.scala 59:15:@62800.4]
  assign FFRAM_io_banks_21_wdata_bits = io_banks_21_wdata_bits; // @[FIFO.scala 59:15:@62799.4]
  assign FFRAM_io_banks_22_wdata_valid = io_banks_22_wdata_valid; // @[FIFO.scala 59:15:@62803.4]
  assign FFRAM_io_banks_22_wdata_bits = io_banks_22_wdata_bits; // @[FIFO.scala 59:15:@62802.4]
  assign FFRAM_io_banks_23_wdata_valid = io_banks_23_wdata_valid; // @[FIFO.scala 59:15:@62806.4]
  assign FFRAM_io_banks_23_wdata_bits = io_banks_23_wdata_bits; // @[FIFO.scala 59:15:@62805.4]
  assign FFRAM_io_banks_24_wdata_valid = io_banks_24_wdata_valid; // @[FIFO.scala 59:15:@62809.4]
  assign FFRAM_io_banks_24_wdata_bits = io_banks_24_wdata_bits; // @[FIFO.scala 59:15:@62808.4]
  assign FFRAM_io_banks_25_wdata_valid = io_banks_25_wdata_valid; // @[FIFO.scala 59:15:@62812.4]
  assign FFRAM_io_banks_25_wdata_bits = io_banks_25_wdata_bits; // @[FIFO.scala 59:15:@62811.4]
  assign FFRAM_io_banks_26_wdata_valid = io_banks_26_wdata_valid; // @[FIFO.scala 59:15:@62815.4]
  assign FFRAM_io_banks_26_wdata_bits = io_banks_26_wdata_bits; // @[FIFO.scala 59:15:@62814.4]
  assign FFRAM_io_banks_27_wdata_valid = io_banks_27_wdata_valid; // @[FIFO.scala 59:15:@62818.4]
  assign FFRAM_io_banks_27_wdata_bits = io_banks_27_wdata_bits; // @[FIFO.scala 59:15:@62817.4]
  assign FFRAM_io_banks_28_wdata_valid = io_banks_28_wdata_valid; // @[FIFO.scala 59:15:@62821.4]
  assign FFRAM_io_banks_28_wdata_bits = io_banks_28_wdata_bits; // @[FIFO.scala 59:15:@62820.4]
  assign FFRAM_io_banks_29_wdata_valid = io_banks_29_wdata_valid; // @[FIFO.scala 59:15:@62824.4]
  assign FFRAM_io_banks_29_wdata_bits = io_banks_29_wdata_bits; // @[FIFO.scala 59:15:@62823.4]
  assign FFRAM_io_banks_30_wdata_valid = io_banks_30_wdata_valid; // @[FIFO.scala 59:15:@62827.4]
  assign FFRAM_io_banks_30_wdata_bits = io_banks_30_wdata_bits; // @[FIFO.scala 59:15:@62826.4]
  assign FFRAM_io_banks_31_wdata_valid = io_banks_31_wdata_valid; // @[FIFO.scala 59:15:@62830.4]
  assign FFRAM_io_banks_31_wdata_bits = io_banks_31_wdata_bits; // @[FIFO.scala 59:15:@62829.4]
  assign FFRAM_io_banks_32_wdata_valid = io_banks_32_wdata_valid; // @[FIFO.scala 59:15:@62833.4]
  assign FFRAM_io_banks_32_wdata_bits = io_banks_32_wdata_bits; // @[FIFO.scala 59:15:@62832.4]
  assign FFRAM_io_banks_33_wdata_valid = io_banks_33_wdata_valid; // @[FIFO.scala 59:15:@62836.4]
  assign FFRAM_io_banks_33_wdata_bits = io_banks_33_wdata_bits; // @[FIFO.scala 59:15:@62835.4]
  assign FFRAM_io_banks_34_wdata_valid = io_banks_34_wdata_valid; // @[FIFO.scala 59:15:@62839.4]
  assign FFRAM_io_banks_34_wdata_bits = io_banks_34_wdata_bits; // @[FIFO.scala 59:15:@62838.4]
  assign FFRAM_io_banks_35_wdata_valid = io_banks_35_wdata_valid; // @[FIFO.scala 59:15:@62842.4]
  assign FFRAM_io_banks_35_wdata_bits = io_banks_35_wdata_bits; // @[FIFO.scala 59:15:@62841.4]
  assign FFRAM_io_banks_36_wdata_valid = io_banks_36_wdata_valid; // @[FIFO.scala 59:15:@62845.4]
  assign FFRAM_io_banks_36_wdata_bits = io_banks_36_wdata_bits; // @[FIFO.scala 59:15:@62844.4]
  assign FFRAM_io_banks_37_wdata_valid = io_banks_37_wdata_valid; // @[FIFO.scala 59:15:@62848.4]
  assign FFRAM_io_banks_37_wdata_bits = io_banks_37_wdata_bits; // @[FIFO.scala 59:15:@62847.4]
  assign FFRAM_io_banks_38_wdata_valid = io_banks_38_wdata_valid; // @[FIFO.scala 59:15:@62851.4]
  assign FFRAM_io_banks_38_wdata_bits = io_banks_38_wdata_bits; // @[FIFO.scala 59:15:@62850.4]
  assign FFRAM_io_banks_39_wdata_valid = io_banks_39_wdata_valid; // @[FIFO.scala 59:15:@62854.4]
  assign FFRAM_io_banks_39_wdata_bits = io_banks_39_wdata_bits; // @[FIFO.scala 59:15:@62853.4]
  assign FFRAM_io_banks_40_wdata_valid = io_banks_40_wdata_valid; // @[FIFO.scala 59:15:@62857.4]
  assign FFRAM_io_banks_40_wdata_bits = io_banks_40_wdata_bits; // @[FIFO.scala 59:15:@62856.4]
  assign FFRAM_io_banks_41_wdata_valid = io_banks_41_wdata_valid; // @[FIFO.scala 59:15:@62860.4]
  assign FFRAM_io_banks_41_wdata_bits = io_banks_41_wdata_bits; // @[FIFO.scala 59:15:@62859.4]
  assign FFRAM_io_banks_42_wdata_valid = io_banks_42_wdata_valid; // @[FIFO.scala 59:15:@62863.4]
  assign FFRAM_io_banks_42_wdata_bits = io_banks_42_wdata_bits; // @[FIFO.scala 59:15:@62862.4]
  assign FFRAM_io_banks_43_wdata_valid = io_banks_43_wdata_valid; // @[FIFO.scala 59:15:@62866.4]
  assign FFRAM_io_banks_43_wdata_bits = io_banks_43_wdata_bits; // @[FIFO.scala 59:15:@62865.4]
  assign FFRAM_io_banks_44_wdata_valid = io_banks_44_wdata_valid; // @[FIFO.scala 59:15:@62869.4]
  assign FFRAM_io_banks_44_wdata_bits = io_banks_44_wdata_bits; // @[FIFO.scala 59:15:@62868.4]
  assign FFRAM_io_banks_45_wdata_valid = io_banks_45_wdata_valid; // @[FIFO.scala 59:15:@62872.4]
  assign FFRAM_io_banks_45_wdata_bits = io_banks_45_wdata_bits; // @[FIFO.scala 59:15:@62871.4]
  assign FFRAM_io_banks_46_wdata_valid = io_banks_46_wdata_valid; // @[FIFO.scala 59:15:@62875.4]
  assign FFRAM_io_banks_46_wdata_bits = io_banks_46_wdata_bits; // @[FIFO.scala 59:15:@62874.4]
  assign FFRAM_io_banks_47_wdata_valid = io_banks_47_wdata_valid; // @[FIFO.scala 59:15:@62878.4]
  assign FFRAM_io_banks_47_wdata_bits = io_banks_47_wdata_bits; // @[FIFO.scala 59:15:@62877.4]
  assign FFRAM_io_banks_48_wdata_valid = io_banks_48_wdata_valid; // @[FIFO.scala 59:15:@62881.4]
  assign FFRAM_io_banks_48_wdata_bits = io_banks_48_wdata_bits; // @[FIFO.scala 59:15:@62880.4]
  assign FFRAM_io_banks_49_wdata_valid = io_banks_49_wdata_valid; // @[FIFO.scala 59:15:@62884.4]
  assign FFRAM_io_banks_49_wdata_bits = io_banks_49_wdata_bits; // @[FIFO.scala 59:15:@62883.4]
  assign FFRAM_io_banks_50_wdata_valid = io_banks_50_wdata_valid; // @[FIFO.scala 59:15:@62887.4]
  assign FFRAM_io_banks_50_wdata_bits = io_banks_50_wdata_bits; // @[FIFO.scala 59:15:@62886.4]
  assign FFRAM_io_banks_51_wdata_valid = io_banks_51_wdata_valid; // @[FIFO.scala 59:15:@62890.4]
  assign FFRAM_io_banks_51_wdata_bits = io_banks_51_wdata_bits; // @[FIFO.scala 59:15:@62889.4]
  assign FFRAM_io_banks_52_wdata_valid = io_banks_52_wdata_valid; // @[FIFO.scala 59:15:@62893.4]
  assign FFRAM_io_banks_52_wdata_bits = io_banks_52_wdata_bits; // @[FIFO.scala 59:15:@62892.4]
  assign FFRAM_io_banks_53_wdata_valid = io_banks_53_wdata_valid; // @[FIFO.scala 59:15:@62896.4]
  assign FFRAM_io_banks_53_wdata_bits = io_banks_53_wdata_bits; // @[FIFO.scala 59:15:@62895.4]
  assign FFRAM_io_banks_54_wdata_valid = io_banks_54_wdata_valid; // @[FIFO.scala 59:15:@62899.4]
  assign FFRAM_io_banks_54_wdata_bits = io_banks_54_wdata_bits; // @[FIFO.scala 59:15:@62898.4]
  assign FFRAM_io_banks_55_wdata_valid = io_banks_55_wdata_valid; // @[FIFO.scala 59:15:@62902.4]
  assign FFRAM_io_banks_55_wdata_bits = io_banks_55_wdata_bits; // @[FIFO.scala 59:15:@62901.4]
  assign FFRAM_io_banks_56_wdata_valid = io_banks_56_wdata_valid; // @[FIFO.scala 59:15:@62905.4]
  assign FFRAM_io_banks_56_wdata_bits = io_banks_56_wdata_bits; // @[FIFO.scala 59:15:@62904.4]
  assign FFRAM_io_banks_57_wdata_valid = io_banks_57_wdata_valid; // @[FIFO.scala 59:15:@62908.4]
  assign FFRAM_io_banks_57_wdata_bits = io_banks_57_wdata_bits; // @[FIFO.scala 59:15:@62907.4]
  assign FFRAM_io_banks_58_wdata_valid = io_banks_58_wdata_valid; // @[FIFO.scala 59:15:@62911.4]
  assign FFRAM_io_banks_58_wdata_bits = io_banks_58_wdata_bits; // @[FIFO.scala 59:15:@62910.4]
  assign FFRAM_io_banks_59_wdata_valid = io_banks_59_wdata_valid; // @[FIFO.scala 59:15:@62914.4]
  assign FFRAM_io_banks_59_wdata_bits = io_banks_59_wdata_bits; // @[FIFO.scala 59:15:@62913.4]
  assign FFRAM_io_banks_60_wdata_valid = io_banks_60_wdata_valid; // @[FIFO.scala 59:15:@62917.4]
  assign FFRAM_io_banks_60_wdata_bits = io_banks_60_wdata_bits; // @[FIFO.scala 59:15:@62916.4]
  assign FFRAM_io_banks_61_wdata_valid = io_banks_61_wdata_valid; // @[FIFO.scala 59:15:@62920.4]
  assign FFRAM_io_banks_61_wdata_bits = io_banks_61_wdata_bits; // @[FIFO.scala 59:15:@62919.4]
  assign FFRAM_io_banks_62_wdata_valid = io_banks_62_wdata_valid; // @[FIFO.scala 59:15:@62923.4]
  assign FFRAM_io_banks_62_wdata_bits = io_banks_62_wdata_bits; // @[FIFO.scala 59:15:@62922.4]
  assign FFRAM_io_banks_63_wdata_valid = io_banks_63_wdata_valid; // @[FIFO.scala 59:15:@62926.4]
  assign FFRAM_io_banks_63_wdata_bits = io_banks_63_wdata_bits; // @[FIFO.scala 59:15:@62925.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_1657) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module StreamControllerStore( // @[:@63705.2]
  input         clock, // @[:@63706.4]
  input         reset, // @[:@63707.4]
  input         io_dram_cmd_ready, // @[:@63708.4]
  output        io_dram_cmd_valid, // @[:@63708.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@63708.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@63708.4]
  input         io_dram_wdata_ready, // @[:@63708.4]
  output        io_dram_wdata_valid, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@63708.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@63708.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@63708.4]
  output        io_dram_wresp_ready, // @[:@63708.4]
  input         io_dram_wresp_valid, // @[:@63708.4]
  output        io_store_cmd_ready, // @[:@63708.4]
  input         io_store_cmd_valid, // @[:@63708.4]
  input  [63:0] io_store_cmd_bits_addr, // @[:@63708.4]
  input  [31:0] io_store_cmd_bits_size, // @[:@63708.4]
  output        io_store_data_ready, // @[:@63708.4]
  input         io_store_data_valid, // @[:@63708.4]
  input  [31:0] io_store_data_bits_wdata_0, // @[:@63708.4]
  input         io_store_data_bits_wstrb, // @[:@63708.4]
  input         io_store_wresp_ready, // @[:@63708.4]
  output        io_store_wresp_valid, // @[:@63708.4]
  output        io_store_wresp_bits // @[:@63708.4]
);
  wire  cmd_clock; // @[StreamController.scala 75:19:@63833.4]
  wire  cmd_reset; // @[StreamController.scala 75:19:@63833.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 75:19:@63833.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 75:19:@63833.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 75:19:@63833.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 75:19:@63833.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 75:19:@63833.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 75:19:@63833.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 75:19:@63833.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 75:19:@63833.4]
  wire  wdata_clock; // @[StreamController.scala 88:21:@64239.4]
  wire  wdata_reset; // @[StreamController.scala 88:21:@64239.4]
  wire  wdata_io_in_ready; // @[StreamController.scala 88:21:@64239.4]
  wire  wdata_io_in_valid; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_in_bits_data_0; // @[StreamController.scala 88:21:@64239.4]
  wire  wdata_io_in_bits_strobe; // @[StreamController.scala 88:21:@64239.4]
  wire  wdata_io_out_ready; // @[StreamController.scala 88:21:@64239.4]
  wire  wdata_io_out_valid; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_0; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_1; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_2; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_3; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_4; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_5; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_6; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_7; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_8; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_9; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_10; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_11; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_12; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_13; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_14; // @[StreamController.scala 88:21:@64239.4]
  wire [31:0] wdata_io_out_bits_data_15; // @[StreamController.scala 88:21:@64239.4]
  wire [63:0] wdata_io_out_bits_strobe; // @[StreamController.scala 88:21:@64239.4]
  wire  wresp_clock; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_reset; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_in_ready; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_in_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_in_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_out_ready; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_out_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_out_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_0_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_0_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_1_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_1_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_2_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_2_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_3_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_3_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_4_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_4_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_5_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_5_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_6_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_6_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_7_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_7_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_8_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_8_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_9_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_9_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_10_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_10_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_11_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_11_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_12_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_12_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_13_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_13_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_14_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_14_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_15_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_15_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_16_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_16_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_17_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_17_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_18_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_18_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_19_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_19_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_20_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_20_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_21_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_21_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_22_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_22_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_23_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_23_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_24_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_24_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_25_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_25_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_26_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_26_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_27_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_27_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_28_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_28_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_29_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_29_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_30_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_30_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_31_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_31_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_32_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_32_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_33_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_33_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_34_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_34_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_35_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_35_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_36_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_36_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_37_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_37_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_38_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_38_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_39_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_39_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_40_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_40_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_41_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_41_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_42_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_42_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_43_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_43_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_44_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_44_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_45_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_45_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_46_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_46_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_47_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_47_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_48_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_48_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_49_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_49_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_50_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_50_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_51_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_51_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_52_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_52_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_53_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_53_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_54_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_54_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_55_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_55_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_56_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_56_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_57_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_57_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_58_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_58_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_59_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_59_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_60_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_60_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_61_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_61_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_62_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_62_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_63_wdata_valid; // @[StreamController.scala 100:21:@64480.4]
  wire  wresp_io_banks_63_wdata_bits; // @[StreamController.scala 100:21:@64480.4]
  wire [25:0] _T_111; // @[StreamController.scala 21:10:@64236.4]
  FIFO cmd ( // @[StreamController.scala 75:19:@63833.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert wdata ( // @[StreamController.scala 88:21:@64239.4]
    .clock(wdata_clock),
    .reset(wdata_reset),
    .io_in_ready(wdata_io_in_ready),
    .io_in_valid(wdata_io_in_valid),
    .io_in_bits_data_0(wdata_io_in_bits_data_0),
    .io_in_bits_strobe(wdata_io_in_bits_strobe),
    .io_out_ready(wdata_io_out_ready),
    .io_out_valid(wdata_io_out_valid),
    .io_out_bits_data_0(wdata_io_out_bits_data_0),
    .io_out_bits_data_1(wdata_io_out_bits_data_1),
    .io_out_bits_data_2(wdata_io_out_bits_data_2),
    .io_out_bits_data_3(wdata_io_out_bits_data_3),
    .io_out_bits_data_4(wdata_io_out_bits_data_4),
    .io_out_bits_data_5(wdata_io_out_bits_data_5),
    .io_out_bits_data_6(wdata_io_out_bits_data_6),
    .io_out_bits_data_7(wdata_io_out_bits_data_7),
    .io_out_bits_data_8(wdata_io_out_bits_data_8),
    .io_out_bits_data_9(wdata_io_out_bits_data_9),
    .io_out_bits_data_10(wdata_io_out_bits_data_10),
    .io_out_bits_data_11(wdata_io_out_bits_data_11),
    .io_out_bits_data_12(wdata_io_out_bits_data_12),
    .io_out_bits_data_13(wdata_io_out_bits_data_13),
    .io_out_bits_data_14(wdata_io_out_bits_data_14),
    .io_out_bits_data_15(wdata_io_out_bits_data_15),
    .io_out_bits_strobe(wdata_io_out_bits_strobe)
  );
  FIFO_33 wresp ( // @[StreamController.scala 100:21:@64480.4]
    .clock(wresp_clock),
    .reset(wresp_reset),
    .io_in_ready(wresp_io_in_ready),
    .io_in_valid(wresp_io_in_valid),
    .io_in_bits(wresp_io_in_bits),
    .io_out_ready(wresp_io_out_ready),
    .io_out_valid(wresp_io_out_valid),
    .io_out_bits(wresp_io_out_bits),
    .io_banks_0_wdata_valid(wresp_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(wresp_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(wresp_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(wresp_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(wresp_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(wresp_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(wresp_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(wresp_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(wresp_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(wresp_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(wresp_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(wresp_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(wresp_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(wresp_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(wresp_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(wresp_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(wresp_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(wresp_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(wresp_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(wresp_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(wresp_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(wresp_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(wresp_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(wresp_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(wresp_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(wresp_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(wresp_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(wresp_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(wresp_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(wresp_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(wresp_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(wresp_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(wresp_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(wresp_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(wresp_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(wresp_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(wresp_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(wresp_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(wresp_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(wresp_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(wresp_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(wresp_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(wresp_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(wresp_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(wresp_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(wresp_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(wresp_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(wresp_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(wresp_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(wresp_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(wresp_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(wresp_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(wresp_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(wresp_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(wresp_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(wresp_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(wresp_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(wresp_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(wresp_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(wresp_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(wresp_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(wresp_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(wresp_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(wresp_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(wresp_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(wresp_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(wresp_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(wresp_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(wresp_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(wresp_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(wresp_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(wresp_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(wresp_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(wresp_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(wresp_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(wresp_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(wresp_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(wresp_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(wresp_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(wresp_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(wresp_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(wresp_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(wresp_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(wresp_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(wresp_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(wresp_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(wresp_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(wresp_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(wresp_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(wresp_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(wresp_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(wresp_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(wresp_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(wresp_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(wresp_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(wresp_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(wresp_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(wresp_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(wresp_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(wresp_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(wresp_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(wresp_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(wresp_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(wresp_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(wresp_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(wresp_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(wresp_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(wresp_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(wresp_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(wresp_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(wresp_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(wresp_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(wresp_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(wresp_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(wresp_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(wresp_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(wresp_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(wresp_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(wresp_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(wresp_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(wresp_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(wresp_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(wresp_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(wresp_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(wresp_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(wresp_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(wresp_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(wresp_io_banks_63_wdata_bits)
  );
  assign _T_111 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@64236.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 81:21:@64233.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 83:25:@64234.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_111}; // @[StreamController.scala 85:25:@64237.4]
  assign io_dram_wdata_valid = wdata_io_out_valid; // @[StreamController.scala 95:23:@64269.4]
  assign io_dram_wdata_bits_wdata_0 = wdata_io_out_bits_data_0; // @[StreamController.scala 96:28:@64270.4]
  assign io_dram_wdata_bits_wdata_1 = wdata_io_out_bits_data_1; // @[StreamController.scala 96:28:@64271.4]
  assign io_dram_wdata_bits_wdata_2 = wdata_io_out_bits_data_2; // @[StreamController.scala 96:28:@64272.4]
  assign io_dram_wdata_bits_wdata_3 = wdata_io_out_bits_data_3; // @[StreamController.scala 96:28:@64273.4]
  assign io_dram_wdata_bits_wdata_4 = wdata_io_out_bits_data_4; // @[StreamController.scala 96:28:@64274.4]
  assign io_dram_wdata_bits_wdata_5 = wdata_io_out_bits_data_5; // @[StreamController.scala 96:28:@64275.4]
  assign io_dram_wdata_bits_wdata_6 = wdata_io_out_bits_data_6; // @[StreamController.scala 96:28:@64276.4]
  assign io_dram_wdata_bits_wdata_7 = wdata_io_out_bits_data_7; // @[StreamController.scala 96:28:@64277.4]
  assign io_dram_wdata_bits_wdata_8 = wdata_io_out_bits_data_8; // @[StreamController.scala 96:28:@64278.4]
  assign io_dram_wdata_bits_wdata_9 = wdata_io_out_bits_data_9; // @[StreamController.scala 96:28:@64279.4]
  assign io_dram_wdata_bits_wdata_10 = wdata_io_out_bits_data_10; // @[StreamController.scala 96:28:@64280.4]
  assign io_dram_wdata_bits_wdata_11 = wdata_io_out_bits_data_11; // @[StreamController.scala 96:28:@64281.4]
  assign io_dram_wdata_bits_wdata_12 = wdata_io_out_bits_data_12; // @[StreamController.scala 96:28:@64282.4]
  assign io_dram_wdata_bits_wdata_13 = wdata_io_out_bits_data_13; // @[StreamController.scala 96:28:@64283.4]
  assign io_dram_wdata_bits_wdata_14 = wdata_io_out_bits_data_14; // @[StreamController.scala 96:28:@64284.4]
  assign io_dram_wdata_bits_wdata_15 = wdata_io_out_bits_data_15; // @[StreamController.scala 96:28:@64285.4]
  assign io_dram_wdata_bits_wstrb_0 = wdata_io_out_bits_strobe[63]; // @[StreamController.scala 97:28:@64415.4]
  assign io_dram_wdata_bits_wstrb_1 = wdata_io_out_bits_strobe[62]; // @[StreamController.scala 97:28:@64416.4]
  assign io_dram_wdata_bits_wstrb_2 = wdata_io_out_bits_strobe[61]; // @[StreamController.scala 97:28:@64417.4]
  assign io_dram_wdata_bits_wstrb_3 = wdata_io_out_bits_strobe[60]; // @[StreamController.scala 97:28:@64418.4]
  assign io_dram_wdata_bits_wstrb_4 = wdata_io_out_bits_strobe[59]; // @[StreamController.scala 97:28:@64419.4]
  assign io_dram_wdata_bits_wstrb_5 = wdata_io_out_bits_strobe[58]; // @[StreamController.scala 97:28:@64420.4]
  assign io_dram_wdata_bits_wstrb_6 = wdata_io_out_bits_strobe[57]; // @[StreamController.scala 97:28:@64421.4]
  assign io_dram_wdata_bits_wstrb_7 = wdata_io_out_bits_strobe[56]; // @[StreamController.scala 97:28:@64422.4]
  assign io_dram_wdata_bits_wstrb_8 = wdata_io_out_bits_strobe[55]; // @[StreamController.scala 97:28:@64423.4]
  assign io_dram_wdata_bits_wstrb_9 = wdata_io_out_bits_strobe[54]; // @[StreamController.scala 97:28:@64424.4]
  assign io_dram_wdata_bits_wstrb_10 = wdata_io_out_bits_strobe[53]; // @[StreamController.scala 97:28:@64425.4]
  assign io_dram_wdata_bits_wstrb_11 = wdata_io_out_bits_strobe[52]; // @[StreamController.scala 97:28:@64426.4]
  assign io_dram_wdata_bits_wstrb_12 = wdata_io_out_bits_strobe[51]; // @[StreamController.scala 97:28:@64427.4]
  assign io_dram_wdata_bits_wstrb_13 = wdata_io_out_bits_strobe[50]; // @[StreamController.scala 97:28:@64428.4]
  assign io_dram_wdata_bits_wstrb_14 = wdata_io_out_bits_strobe[49]; // @[StreamController.scala 97:28:@64429.4]
  assign io_dram_wdata_bits_wstrb_15 = wdata_io_out_bits_strobe[48]; // @[StreamController.scala 97:28:@64430.4]
  assign io_dram_wdata_bits_wstrb_16 = wdata_io_out_bits_strobe[47]; // @[StreamController.scala 97:28:@64431.4]
  assign io_dram_wdata_bits_wstrb_17 = wdata_io_out_bits_strobe[46]; // @[StreamController.scala 97:28:@64432.4]
  assign io_dram_wdata_bits_wstrb_18 = wdata_io_out_bits_strobe[45]; // @[StreamController.scala 97:28:@64433.4]
  assign io_dram_wdata_bits_wstrb_19 = wdata_io_out_bits_strobe[44]; // @[StreamController.scala 97:28:@64434.4]
  assign io_dram_wdata_bits_wstrb_20 = wdata_io_out_bits_strobe[43]; // @[StreamController.scala 97:28:@64435.4]
  assign io_dram_wdata_bits_wstrb_21 = wdata_io_out_bits_strobe[42]; // @[StreamController.scala 97:28:@64436.4]
  assign io_dram_wdata_bits_wstrb_22 = wdata_io_out_bits_strobe[41]; // @[StreamController.scala 97:28:@64437.4]
  assign io_dram_wdata_bits_wstrb_23 = wdata_io_out_bits_strobe[40]; // @[StreamController.scala 97:28:@64438.4]
  assign io_dram_wdata_bits_wstrb_24 = wdata_io_out_bits_strobe[39]; // @[StreamController.scala 97:28:@64439.4]
  assign io_dram_wdata_bits_wstrb_25 = wdata_io_out_bits_strobe[38]; // @[StreamController.scala 97:28:@64440.4]
  assign io_dram_wdata_bits_wstrb_26 = wdata_io_out_bits_strobe[37]; // @[StreamController.scala 97:28:@64441.4]
  assign io_dram_wdata_bits_wstrb_27 = wdata_io_out_bits_strobe[36]; // @[StreamController.scala 97:28:@64442.4]
  assign io_dram_wdata_bits_wstrb_28 = wdata_io_out_bits_strobe[35]; // @[StreamController.scala 97:28:@64443.4]
  assign io_dram_wdata_bits_wstrb_29 = wdata_io_out_bits_strobe[34]; // @[StreamController.scala 97:28:@64444.4]
  assign io_dram_wdata_bits_wstrb_30 = wdata_io_out_bits_strobe[33]; // @[StreamController.scala 97:28:@64445.4]
  assign io_dram_wdata_bits_wstrb_31 = wdata_io_out_bits_strobe[32]; // @[StreamController.scala 97:28:@64446.4]
  assign io_dram_wdata_bits_wstrb_32 = wdata_io_out_bits_strobe[31]; // @[StreamController.scala 97:28:@64447.4]
  assign io_dram_wdata_bits_wstrb_33 = wdata_io_out_bits_strobe[30]; // @[StreamController.scala 97:28:@64448.4]
  assign io_dram_wdata_bits_wstrb_34 = wdata_io_out_bits_strobe[29]; // @[StreamController.scala 97:28:@64449.4]
  assign io_dram_wdata_bits_wstrb_35 = wdata_io_out_bits_strobe[28]; // @[StreamController.scala 97:28:@64450.4]
  assign io_dram_wdata_bits_wstrb_36 = wdata_io_out_bits_strobe[27]; // @[StreamController.scala 97:28:@64451.4]
  assign io_dram_wdata_bits_wstrb_37 = wdata_io_out_bits_strobe[26]; // @[StreamController.scala 97:28:@64452.4]
  assign io_dram_wdata_bits_wstrb_38 = wdata_io_out_bits_strobe[25]; // @[StreamController.scala 97:28:@64453.4]
  assign io_dram_wdata_bits_wstrb_39 = wdata_io_out_bits_strobe[24]; // @[StreamController.scala 97:28:@64454.4]
  assign io_dram_wdata_bits_wstrb_40 = wdata_io_out_bits_strobe[23]; // @[StreamController.scala 97:28:@64455.4]
  assign io_dram_wdata_bits_wstrb_41 = wdata_io_out_bits_strobe[22]; // @[StreamController.scala 97:28:@64456.4]
  assign io_dram_wdata_bits_wstrb_42 = wdata_io_out_bits_strobe[21]; // @[StreamController.scala 97:28:@64457.4]
  assign io_dram_wdata_bits_wstrb_43 = wdata_io_out_bits_strobe[20]; // @[StreamController.scala 97:28:@64458.4]
  assign io_dram_wdata_bits_wstrb_44 = wdata_io_out_bits_strobe[19]; // @[StreamController.scala 97:28:@64459.4]
  assign io_dram_wdata_bits_wstrb_45 = wdata_io_out_bits_strobe[18]; // @[StreamController.scala 97:28:@64460.4]
  assign io_dram_wdata_bits_wstrb_46 = wdata_io_out_bits_strobe[17]; // @[StreamController.scala 97:28:@64461.4]
  assign io_dram_wdata_bits_wstrb_47 = wdata_io_out_bits_strobe[16]; // @[StreamController.scala 97:28:@64462.4]
  assign io_dram_wdata_bits_wstrb_48 = wdata_io_out_bits_strobe[15]; // @[StreamController.scala 97:28:@64463.4]
  assign io_dram_wdata_bits_wstrb_49 = wdata_io_out_bits_strobe[14]; // @[StreamController.scala 97:28:@64464.4]
  assign io_dram_wdata_bits_wstrb_50 = wdata_io_out_bits_strobe[13]; // @[StreamController.scala 97:28:@64465.4]
  assign io_dram_wdata_bits_wstrb_51 = wdata_io_out_bits_strobe[12]; // @[StreamController.scala 97:28:@64466.4]
  assign io_dram_wdata_bits_wstrb_52 = wdata_io_out_bits_strobe[11]; // @[StreamController.scala 97:28:@64467.4]
  assign io_dram_wdata_bits_wstrb_53 = wdata_io_out_bits_strobe[10]; // @[StreamController.scala 97:28:@64468.4]
  assign io_dram_wdata_bits_wstrb_54 = wdata_io_out_bits_strobe[9]; // @[StreamController.scala 97:28:@64469.4]
  assign io_dram_wdata_bits_wstrb_55 = wdata_io_out_bits_strobe[8]; // @[StreamController.scala 97:28:@64470.4]
  assign io_dram_wdata_bits_wstrb_56 = wdata_io_out_bits_strobe[7]; // @[StreamController.scala 97:28:@64471.4]
  assign io_dram_wdata_bits_wstrb_57 = wdata_io_out_bits_strobe[6]; // @[StreamController.scala 97:28:@64472.4]
  assign io_dram_wdata_bits_wstrb_58 = wdata_io_out_bits_strobe[5]; // @[StreamController.scala 97:28:@64473.4]
  assign io_dram_wdata_bits_wstrb_59 = wdata_io_out_bits_strobe[4]; // @[StreamController.scala 97:28:@64474.4]
  assign io_dram_wdata_bits_wstrb_60 = wdata_io_out_bits_strobe[3]; // @[StreamController.scala 97:28:@64475.4]
  assign io_dram_wdata_bits_wstrb_61 = wdata_io_out_bits_strobe[2]; // @[StreamController.scala 97:28:@64476.4]
  assign io_dram_wdata_bits_wstrb_62 = wdata_io_out_bits_strobe[1]; // @[StreamController.scala 97:28:@64477.4]
  assign io_dram_wdata_bits_wstrb_63 = wdata_io_out_bits_strobe[0]; // @[StreamController.scala 97:28:@64478.4]
  assign io_dram_wresp_ready = wresp_io_in_ready; // @[StreamController.scala 104:23:@64747.4]
  assign io_store_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 79:22:@64231.4]
  assign io_store_data_ready = wdata_io_in_ready; // @[StreamController.scala 93:23:@64268.4]
  assign io_store_wresp_valid = wresp_io_out_valid; // @[StreamController.scala 106:24:@64748.4]
  assign io_store_wresp_bits = wresp_io_out_bits; // @[StreamController.scala 107:23:@64749.4]
  assign cmd_clock = clock; // @[:@63834.4]
  assign cmd_reset = reset; // @[:@63835.4]
  assign cmd_io_in_valid = io_store_cmd_valid; // @[StreamController.scala 77:19:@64228.4]
  assign cmd_io_in_bits_addr = io_store_cmd_bits_addr; // @[StreamController.scala 78:18:@64230.4]
  assign cmd_io_in_bits_size = io_store_cmd_bits_size; // @[StreamController.scala 78:18:@64229.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 80:20:@64232.4]
  assign wdata_clock = clock; // @[:@64240.4]
  assign wdata_reset = reset; // @[:@64241.4]
  assign wdata_io_in_valid = io_store_data_valid; // @[StreamController.scala 90:21:@64265.4]
  assign wdata_io_in_bits_data_0 = io_store_data_bits_wdata_0; // @[StreamController.scala 91:25:@64266.4]
  assign wdata_io_in_bits_strobe = io_store_data_bits_wstrb; // @[StreamController.scala 92:27:@64267.4]
  assign wdata_io_out_ready = io_dram_wdata_ready; // @[StreamController.scala 98:22:@64479.4]
  assign wresp_clock = clock; // @[:@64481.4]
  assign wresp_reset = reset; // @[:@64482.4]
  assign wresp_io_in_valid = io_dram_wresp_valid; // @[StreamController.scala 102:21:@64745.4]
  assign wresp_io_in_bits = 1'h1; // @[StreamController.scala 103:20:@64746.4]
  assign wresp_io_out_ready = io_store_wresp_ready; // @[StreamController.scala 108:22:@64750.4]
  assign wresp_io_banks_0_wdata_valid = 1'h0;
  assign wresp_io_banks_0_wdata_bits = 1'h0;
  assign wresp_io_banks_1_wdata_valid = 1'h0;
  assign wresp_io_banks_1_wdata_bits = 1'h0;
  assign wresp_io_banks_2_wdata_valid = 1'h0;
  assign wresp_io_banks_2_wdata_bits = 1'h0;
  assign wresp_io_banks_3_wdata_valid = 1'h0;
  assign wresp_io_banks_3_wdata_bits = 1'h0;
  assign wresp_io_banks_4_wdata_valid = 1'h0;
  assign wresp_io_banks_4_wdata_bits = 1'h0;
  assign wresp_io_banks_5_wdata_valid = 1'h0;
  assign wresp_io_banks_5_wdata_bits = 1'h0;
  assign wresp_io_banks_6_wdata_valid = 1'h0;
  assign wresp_io_banks_6_wdata_bits = 1'h0;
  assign wresp_io_banks_7_wdata_valid = 1'h0;
  assign wresp_io_banks_7_wdata_bits = 1'h0;
  assign wresp_io_banks_8_wdata_valid = 1'h0;
  assign wresp_io_banks_8_wdata_bits = 1'h0;
  assign wresp_io_banks_9_wdata_valid = 1'h0;
  assign wresp_io_banks_9_wdata_bits = 1'h0;
  assign wresp_io_banks_10_wdata_valid = 1'h0;
  assign wresp_io_banks_10_wdata_bits = 1'h0;
  assign wresp_io_banks_11_wdata_valid = 1'h0;
  assign wresp_io_banks_11_wdata_bits = 1'h0;
  assign wresp_io_banks_12_wdata_valid = 1'h0;
  assign wresp_io_banks_12_wdata_bits = 1'h0;
  assign wresp_io_banks_13_wdata_valid = 1'h0;
  assign wresp_io_banks_13_wdata_bits = 1'h0;
  assign wresp_io_banks_14_wdata_valid = 1'h0;
  assign wresp_io_banks_14_wdata_bits = 1'h0;
  assign wresp_io_banks_15_wdata_valid = 1'h0;
  assign wresp_io_banks_15_wdata_bits = 1'h0;
  assign wresp_io_banks_16_wdata_valid = 1'h0;
  assign wresp_io_banks_16_wdata_bits = 1'h0;
  assign wresp_io_banks_17_wdata_valid = 1'h0;
  assign wresp_io_banks_17_wdata_bits = 1'h0;
  assign wresp_io_banks_18_wdata_valid = 1'h0;
  assign wresp_io_banks_18_wdata_bits = 1'h0;
  assign wresp_io_banks_19_wdata_valid = 1'h0;
  assign wresp_io_banks_19_wdata_bits = 1'h0;
  assign wresp_io_banks_20_wdata_valid = 1'h0;
  assign wresp_io_banks_20_wdata_bits = 1'h0;
  assign wresp_io_banks_21_wdata_valid = 1'h0;
  assign wresp_io_banks_21_wdata_bits = 1'h0;
  assign wresp_io_banks_22_wdata_valid = 1'h0;
  assign wresp_io_banks_22_wdata_bits = 1'h0;
  assign wresp_io_banks_23_wdata_valid = 1'h0;
  assign wresp_io_banks_23_wdata_bits = 1'h0;
  assign wresp_io_banks_24_wdata_valid = 1'h0;
  assign wresp_io_banks_24_wdata_bits = 1'h0;
  assign wresp_io_banks_25_wdata_valid = 1'h0;
  assign wresp_io_banks_25_wdata_bits = 1'h0;
  assign wresp_io_banks_26_wdata_valid = 1'h0;
  assign wresp_io_banks_26_wdata_bits = 1'h0;
  assign wresp_io_banks_27_wdata_valid = 1'h0;
  assign wresp_io_banks_27_wdata_bits = 1'h0;
  assign wresp_io_banks_28_wdata_valid = 1'h0;
  assign wresp_io_banks_28_wdata_bits = 1'h0;
  assign wresp_io_banks_29_wdata_valid = 1'h0;
  assign wresp_io_banks_29_wdata_bits = 1'h0;
  assign wresp_io_banks_30_wdata_valid = 1'h0;
  assign wresp_io_banks_30_wdata_bits = 1'h0;
  assign wresp_io_banks_31_wdata_valid = 1'h0;
  assign wresp_io_banks_31_wdata_bits = 1'h0;
  assign wresp_io_banks_32_wdata_valid = 1'h0;
  assign wresp_io_banks_32_wdata_bits = 1'h0;
  assign wresp_io_banks_33_wdata_valid = 1'h0;
  assign wresp_io_banks_33_wdata_bits = 1'h0;
  assign wresp_io_banks_34_wdata_valid = 1'h0;
  assign wresp_io_banks_34_wdata_bits = 1'h0;
  assign wresp_io_banks_35_wdata_valid = 1'h0;
  assign wresp_io_banks_35_wdata_bits = 1'h0;
  assign wresp_io_banks_36_wdata_valid = 1'h0;
  assign wresp_io_banks_36_wdata_bits = 1'h0;
  assign wresp_io_banks_37_wdata_valid = 1'h0;
  assign wresp_io_banks_37_wdata_bits = 1'h0;
  assign wresp_io_banks_38_wdata_valid = 1'h0;
  assign wresp_io_banks_38_wdata_bits = 1'h0;
  assign wresp_io_banks_39_wdata_valid = 1'h0;
  assign wresp_io_banks_39_wdata_bits = 1'h0;
  assign wresp_io_banks_40_wdata_valid = 1'h0;
  assign wresp_io_banks_40_wdata_bits = 1'h0;
  assign wresp_io_banks_41_wdata_valid = 1'h0;
  assign wresp_io_banks_41_wdata_bits = 1'h0;
  assign wresp_io_banks_42_wdata_valid = 1'h0;
  assign wresp_io_banks_42_wdata_bits = 1'h0;
  assign wresp_io_banks_43_wdata_valid = 1'h0;
  assign wresp_io_banks_43_wdata_bits = 1'h0;
  assign wresp_io_banks_44_wdata_valid = 1'h0;
  assign wresp_io_banks_44_wdata_bits = 1'h0;
  assign wresp_io_banks_45_wdata_valid = 1'h0;
  assign wresp_io_banks_45_wdata_bits = 1'h0;
  assign wresp_io_banks_46_wdata_valid = 1'h0;
  assign wresp_io_banks_46_wdata_bits = 1'h0;
  assign wresp_io_banks_47_wdata_valid = 1'h0;
  assign wresp_io_banks_47_wdata_bits = 1'h0;
  assign wresp_io_banks_48_wdata_valid = 1'h0;
  assign wresp_io_banks_48_wdata_bits = 1'h0;
  assign wresp_io_banks_49_wdata_valid = 1'h0;
  assign wresp_io_banks_49_wdata_bits = 1'h0;
  assign wresp_io_banks_50_wdata_valid = 1'h0;
  assign wresp_io_banks_50_wdata_bits = 1'h0;
  assign wresp_io_banks_51_wdata_valid = 1'h0;
  assign wresp_io_banks_51_wdata_bits = 1'h0;
  assign wresp_io_banks_52_wdata_valid = 1'h0;
  assign wresp_io_banks_52_wdata_bits = 1'h0;
  assign wresp_io_banks_53_wdata_valid = 1'h0;
  assign wresp_io_banks_53_wdata_bits = 1'h0;
  assign wresp_io_banks_54_wdata_valid = 1'h0;
  assign wresp_io_banks_54_wdata_bits = 1'h0;
  assign wresp_io_banks_55_wdata_valid = 1'h0;
  assign wresp_io_banks_55_wdata_bits = 1'h0;
  assign wresp_io_banks_56_wdata_valid = 1'h0;
  assign wresp_io_banks_56_wdata_bits = 1'h0;
  assign wresp_io_banks_57_wdata_valid = 1'h0;
  assign wresp_io_banks_57_wdata_bits = 1'h0;
  assign wresp_io_banks_58_wdata_valid = 1'h0;
  assign wresp_io_banks_58_wdata_bits = 1'h0;
  assign wresp_io_banks_59_wdata_valid = 1'h0;
  assign wresp_io_banks_59_wdata_bits = 1'h0;
  assign wresp_io_banks_60_wdata_valid = 1'h0;
  assign wresp_io_banks_60_wdata_bits = 1'h0;
  assign wresp_io_banks_61_wdata_valid = 1'h0;
  assign wresp_io_banks_61_wdata_bits = 1'h0;
  assign wresp_io_banks_62_wdata_valid = 1'h0;
  assign wresp_io_banks_62_wdata_bits = 1'h0;
  assign wresp_io_banks_63_wdata_valid = 1'h0;
  assign wresp_io_banks_63_wdata_bits = 1'h0;
endmodule
module MuxPipe( // @[:@64816.2]
  output        io_in_ready, // @[:@64819.4]
  input         io_in_valid, // @[:@64819.4]
  input  [63:0] io_in_bits_0_addr, // @[:@64819.4]
  input  [31:0] io_in_bits_0_size, // @[:@64819.4]
  input         io_in_bits_0_isWr, // @[:@64819.4]
  input  [31:0] io_in_bits_0_tag, // @[:@64819.4]
  input         io_out_ready, // @[:@64819.4]
  output        io_out_valid, // @[:@64819.4]
  output [63:0] io_out_bits_addr, // @[:@64819.4]
  output [31:0] io_out_bits_size, // @[:@64819.4]
  output        io_out_bits_isWr, // @[:@64819.4]
  output [31:0] io_out_bits_tag // @[:@64819.4]
);
  wire  _T_42; // @[MuxN.scala 28:31:@64821.4]
  assign _T_42 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@64821.4]
  assign io_in_ready = io_out_ready | _T_42; // @[MuxN.scala 71:15:@64830.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@64829.4]
  assign io_out_bits_addr = io_in_bits_0_addr; // @[MuxN.scala 72:15:@64835.4]
  assign io_out_bits_size = io_in_bits_0_size; // @[MuxN.scala 72:15:@64834.4]
  assign io_out_bits_isWr = io_in_bits_0_isWr; // @[MuxN.scala 72:15:@64832.4]
  assign io_out_bits_tag = io_in_bits_0_tag; // @[MuxN.scala 72:15:@64831.4]
endmodule
module MuxPipe_1( // @[:@64837.2]
  output        io_in_ready, // @[:@64840.4]
  input         io_in_valid, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_0, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_1, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_2, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_3, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_4, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_5, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_6, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_7, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_8, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_9, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_10, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_11, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_12, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_13, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_14, // @[:@64840.4]
  input  [31:0] io_in_bits_0_wdata_15, // @[:@64840.4]
  input         io_in_bits_0_wstrb_0, // @[:@64840.4]
  input         io_in_bits_0_wstrb_1, // @[:@64840.4]
  input         io_in_bits_0_wstrb_2, // @[:@64840.4]
  input         io_in_bits_0_wstrb_3, // @[:@64840.4]
  input         io_in_bits_0_wstrb_4, // @[:@64840.4]
  input         io_in_bits_0_wstrb_5, // @[:@64840.4]
  input         io_in_bits_0_wstrb_6, // @[:@64840.4]
  input         io_in_bits_0_wstrb_7, // @[:@64840.4]
  input         io_in_bits_0_wstrb_8, // @[:@64840.4]
  input         io_in_bits_0_wstrb_9, // @[:@64840.4]
  input         io_in_bits_0_wstrb_10, // @[:@64840.4]
  input         io_in_bits_0_wstrb_11, // @[:@64840.4]
  input         io_in_bits_0_wstrb_12, // @[:@64840.4]
  input         io_in_bits_0_wstrb_13, // @[:@64840.4]
  input         io_in_bits_0_wstrb_14, // @[:@64840.4]
  input         io_in_bits_0_wstrb_15, // @[:@64840.4]
  input         io_in_bits_0_wstrb_16, // @[:@64840.4]
  input         io_in_bits_0_wstrb_17, // @[:@64840.4]
  input         io_in_bits_0_wstrb_18, // @[:@64840.4]
  input         io_in_bits_0_wstrb_19, // @[:@64840.4]
  input         io_in_bits_0_wstrb_20, // @[:@64840.4]
  input         io_in_bits_0_wstrb_21, // @[:@64840.4]
  input         io_in_bits_0_wstrb_22, // @[:@64840.4]
  input         io_in_bits_0_wstrb_23, // @[:@64840.4]
  input         io_in_bits_0_wstrb_24, // @[:@64840.4]
  input         io_in_bits_0_wstrb_25, // @[:@64840.4]
  input         io_in_bits_0_wstrb_26, // @[:@64840.4]
  input         io_in_bits_0_wstrb_27, // @[:@64840.4]
  input         io_in_bits_0_wstrb_28, // @[:@64840.4]
  input         io_in_bits_0_wstrb_29, // @[:@64840.4]
  input         io_in_bits_0_wstrb_30, // @[:@64840.4]
  input         io_in_bits_0_wstrb_31, // @[:@64840.4]
  input         io_in_bits_0_wstrb_32, // @[:@64840.4]
  input         io_in_bits_0_wstrb_33, // @[:@64840.4]
  input         io_in_bits_0_wstrb_34, // @[:@64840.4]
  input         io_in_bits_0_wstrb_35, // @[:@64840.4]
  input         io_in_bits_0_wstrb_36, // @[:@64840.4]
  input         io_in_bits_0_wstrb_37, // @[:@64840.4]
  input         io_in_bits_0_wstrb_38, // @[:@64840.4]
  input         io_in_bits_0_wstrb_39, // @[:@64840.4]
  input         io_in_bits_0_wstrb_40, // @[:@64840.4]
  input         io_in_bits_0_wstrb_41, // @[:@64840.4]
  input         io_in_bits_0_wstrb_42, // @[:@64840.4]
  input         io_in_bits_0_wstrb_43, // @[:@64840.4]
  input         io_in_bits_0_wstrb_44, // @[:@64840.4]
  input         io_in_bits_0_wstrb_45, // @[:@64840.4]
  input         io_in_bits_0_wstrb_46, // @[:@64840.4]
  input         io_in_bits_0_wstrb_47, // @[:@64840.4]
  input         io_in_bits_0_wstrb_48, // @[:@64840.4]
  input         io_in_bits_0_wstrb_49, // @[:@64840.4]
  input         io_in_bits_0_wstrb_50, // @[:@64840.4]
  input         io_in_bits_0_wstrb_51, // @[:@64840.4]
  input         io_in_bits_0_wstrb_52, // @[:@64840.4]
  input         io_in_bits_0_wstrb_53, // @[:@64840.4]
  input         io_in_bits_0_wstrb_54, // @[:@64840.4]
  input         io_in_bits_0_wstrb_55, // @[:@64840.4]
  input         io_in_bits_0_wstrb_56, // @[:@64840.4]
  input         io_in_bits_0_wstrb_57, // @[:@64840.4]
  input         io_in_bits_0_wstrb_58, // @[:@64840.4]
  input         io_in_bits_0_wstrb_59, // @[:@64840.4]
  input         io_in_bits_0_wstrb_60, // @[:@64840.4]
  input         io_in_bits_0_wstrb_61, // @[:@64840.4]
  input         io_in_bits_0_wstrb_62, // @[:@64840.4]
  input         io_in_bits_0_wstrb_63, // @[:@64840.4]
  input         io_out_ready, // @[:@64840.4]
  output        io_out_valid, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_0, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_1, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_2, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_3, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_4, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_5, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_6, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_7, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_8, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_9, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_10, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_11, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_12, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_13, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_14, // @[:@64840.4]
  output [31:0] io_out_bits_wdata_15, // @[:@64840.4]
  output        io_out_bits_wstrb_0, // @[:@64840.4]
  output        io_out_bits_wstrb_1, // @[:@64840.4]
  output        io_out_bits_wstrb_2, // @[:@64840.4]
  output        io_out_bits_wstrb_3, // @[:@64840.4]
  output        io_out_bits_wstrb_4, // @[:@64840.4]
  output        io_out_bits_wstrb_5, // @[:@64840.4]
  output        io_out_bits_wstrb_6, // @[:@64840.4]
  output        io_out_bits_wstrb_7, // @[:@64840.4]
  output        io_out_bits_wstrb_8, // @[:@64840.4]
  output        io_out_bits_wstrb_9, // @[:@64840.4]
  output        io_out_bits_wstrb_10, // @[:@64840.4]
  output        io_out_bits_wstrb_11, // @[:@64840.4]
  output        io_out_bits_wstrb_12, // @[:@64840.4]
  output        io_out_bits_wstrb_13, // @[:@64840.4]
  output        io_out_bits_wstrb_14, // @[:@64840.4]
  output        io_out_bits_wstrb_15, // @[:@64840.4]
  output        io_out_bits_wstrb_16, // @[:@64840.4]
  output        io_out_bits_wstrb_17, // @[:@64840.4]
  output        io_out_bits_wstrb_18, // @[:@64840.4]
  output        io_out_bits_wstrb_19, // @[:@64840.4]
  output        io_out_bits_wstrb_20, // @[:@64840.4]
  output        io_out_bits_wstrb_21, // @[:@64840.4]
  output        io_out_bits_wstrb_22, // @[:@64840.4]
  output        io_out_bits_wstrb_23, // @[:@64840.4]
  output        io_out_bits_wstrb_24, // @[:@64840.4]
  output        io_out_bits_wstrb_25, // @[:@64840.4]
  output        io_out_bits_wstrb_26, // @[:@64840.4]
  output        io_out_bits_wstrb_27, // @[:@64840.4]
  output        io_out_bits_wstrb_28, // @[:@64840.4]
  output        io_out_bits_wstrb_29, // @[:@64840.4]
  output        io_out_bits_wstrb_30, // @[:@64840.4]
  output        io_out_bits_wstrb_31, // @[:@64840.4]
  output        io_out_bits_wstrb_32, // @[:@64840.4]
  output        io_out_bits_wstrb_33, // @[:@64840.4]
  output        io_out_bits_wstrb_34, // @[:@64840.4]
  output        io_out_bits_wstrb_35, // @[:@64840.4]
  output        io_out_bits_wstrb_36, // @[:@64840.4]
  output        io_out_bits_wstrb_37, // @[:@64840.4]
  output        io_out_bits_wstrb_38, // @[:@64840.4]
  output        io_out_bits_wstrb_39, // @[:@64840.4]
  output        io_out_bits_wstrb_40, // @[:@64840.4]
  output        io_out_bits_wstrb_41, // @[:@64840.4]
  output        io_out_bits_wstrb_42, // @[:@64840.4]
  output        io_out_bits_wstrb_43, // @[:@64840.4]
  output        io_out_bits_wstrb_44, // @[:@64840.4]
  output        io_out_bits_wstrb_45, // @[:@64840.4]
  output        io_out_bits_wstrb_46, // @[:@64840.4]
  output        io_out_bits_wstrb_47, // @[:@64840.4]
  output        io_out_bits_wstrb_48, // @[:@64840.4]
  output        io_out_bits_wstrb_49, // @[:@64840.4]
  output        io_out_bits_wstrb_50, // @[:@64840.4]
  output        io_out_bits_wstrb_51, // @[:@64840.4]
  output        io_out_bits_wstrb_52, // @[:@64840.4]
  output        io_out_bits_wstrb_53, // @[:@64840.4]
  output        io_out_bits_wstrb_54, // @[:@64840.4]
  output        io_out_bits_wstrb_55, // @[:@64840.4]
  output        io_out_bits_wstrb_56, // @[:@64840.4]
  output        io_out_bits_wstrb_57, // @[:@64840.4]
  output        io_out_bits_wstrb_58, // @[:@64840.4]
  output        io_out_bits_wstrb_59, // @[:@64840.4]
  output        io_out_bits_wstrb_60, // @[:@64840.4]
  output        io_out_bits_wstrb_61, // @[:@64840.4]
  output        io_out_bits_wstrb_62, // @[:@64840.4]
  output        io_out_bits_wstrb_63 // @[:@64840.4]
);
  wire  _T_146; // @[MuxN.scala 28:31:@64842.4]
  assign _T_146 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@64842.4]
  assign io_in_ready = io_out_ready | _T_146; // @[MuxN.scala 71:15:@64927.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@64926.4]
  assign io_out_bits_wdata_0 = io_in_bits_0_wdata_0; // @[MuxN.scala 72:15:@64993.4]
  assign io_out_bits_wdata_1 = io_in_bits_0_wdata_1; // @[MuxN.scala 72:15:@64994.4]
  assign io_out_bits_wdata_2 = io_in_bits_0_wdata_2; // @[MuxN.scala 72:15:@64995.4]
  assign io_out_bits_wdata_3 = io_in_bits_0_wdata_3; // @[MuxN.scala 72:15:@64996.4]
  assign io_out_bits_wdata_4 = io_in_bits_0_wdata_4; // @[MuxN.scala 72:15:@64997.4]
  assign io_out_bits_wdata_5 = io_in_bits_0_wdata_5; // @[MuxN.scala 72:15:@64998.4]
  assign io_out_bits_wdata_6 = io_in_bits_0_wdata_6; // @[MuxN.scala 72:15:@64999.4]
  assign io_out_bits_wdata_7 = io_in_bits_0_wdata_7; // @[MuxN.scala 72:15:@65000.4]
  assign io_out_bits_wdata_8 = io_in_bits_0_wdata_8; // @[MuxN.scala 72:15:@65001.4]
  assign io_out_bits_wdata_9 = io_in_bits_0_wdata_9; // @[MuxN.scala 72:15:@65002.4]
  assign io_out_bits_wdata_10 = io_in_bits_0_wdata_10; // @[MuxN.scala 72:15:@65003.4]
  assign io_out_bits_wdata_11 = io_in_bits_0_wdata_11; // @[MuxN.scala 72:15:@65004.4]
  assign io_out_bits_wdata_12 = io_in_bits_0_wdata_12; // @[MuxN.scala 72:15:@65005.4]
  assign io_out_bits_wdata_13 = io_in_bits_0_wdata_13; // @[MuxN.scala 72:15:@65006.4]
  assign io_out_bits_wdata_14 = io_in_bits_0_wdata_14; // @[MuxN.scala 72:15:@65007.4]
  assign io_out_bits_wdata_15 = io_in_bits_0_wdata_15; // @[MuxN.scala 72:15:@65008.4]
  assign io_out_bits_wstrb_0 = io_in_bits_0_wstrb_0; // @[MuxN.scala 72:15:@64929.4]
  assign io_out_bits_wstrb_1 = io_in_bits_0_wstrb_1; // @[MuxN.scala 72:15:@64930.4]
  assign io_out_bits_wstrb_2 = io_in_bits_0_wstrb_2; // @[MuxN.scala 72:15:@64931.4]
  assign io_out_bits_wstrb_3 = io_in_bits_0_wstrb_3; // @[MuxN.scala 72:15:@64932.4]
  assign io_out_bits_wstrb_4 = io_in_bits_0_wstrb_4; // @[MuxN.scala 72:15:@64933.4]
  assign io_out_bits_wstrb_5 = io_in_bits_0_wstrb_5; // @[MuxN.scala 72:15:@64934.4]
  assign io_out_bits_wstrb_6 = io_in_bits_0_wstrb_6; // @[MuxN.scala 72:15:@64935.4]
  assign io_out_bits_wstrb_7 = io_in_bits_0_wstrb_7; // @[MuxN.scala 72:15:@64936.4]
  assign io_out_bits_wstrb_8 = io_in_bits_0_wstrb_8; // @[MuxN.scala 72:15:@64937.4]
  assign io_out_bits_wstrb_9 = io_in_bits_0_wstrb_9; // @[MuxN.scala 72:15:@64938.4]
  assign io_out_bits_wstrb_10 = io_in_bits_0_wstrb_10; // @[MuxN.scala 72:15:@64939.4]
  assign io_out_bits_wstrb_11 = io_in_bits_0_wstrb_11; // @[MuxN.scala 72:15:@64940.4]
  assign io_out_bits_wstrb_12 = io_in_bits_0_wstrb_12; // @[MuxN.scala 72:15:@64941.4]
  assign io_out_bits_wstrb_13 = io_in_bits_0_wstrb_13; // @[MuxN.scala 72:15:@64942.4]
  assign io_out_bits_wstrb_14 = io_in_bits_0_wstrb_14; // @[MuxN.scala 72:15:@64943.4]
  assign io_out_bits_wstrb_15 = io_in_bits_0_wstrb_15; // @[MuxN.scala 72:15:@64944.4]
  assign io_out_bits_wstrb_16 = io_in_bits_0_wstrb_16; // @[MuxN.scala 72:15:@64945.4]
  assign io_out_bits_wstrb_17 = io_in_bits_0_wstrb_17; // @[MuxN.scala 72:15:@64946.4]
  assign io_out_bits_wstrb_18 = io_in_bits_0_wstrb_18; // @[MuxN.scala 72:15:@64947.4]
  assign io_out_bits_wstrb_19 = io_in_bits_0_wstrb_19; // @[MuxN.scala 72:15:@64948.4]
  assign io_out_bits_wstrb_20 = io_in_bits_0_wstrb_20; // @[MuxN.scala 72:15:@64949.4]
  assign io_out_bits_wstrb_21 = io_in_bits_0_wstrb_21; // @[MuxN.scala 72:15:@64950.4]
  assign io_out_bits_wstrb_22 = io_in_bits_0_wstrb_22; // @[MuxN.scala 72:15:@64951.4]
  assign io_out_bits_wstrb_23 = io_in_bits_0_wstrb_23; // @[MuxN.scala 72:15:@64952.4]
  assign io_out_bits_wstrb_24 = io_in_bits_0_wstrb_24; // @[MuxN.scala 72:15:@64953.4]
  assign io_out_bits_wstrb_25 = io_in_bits_0_wstrb_25; // @[MuxN.scala 72:15:@64954.4]
  assign io_out_bits_wstrb_26 = io_in_bits_0_wstrb_26; // @[MuxN.scala 72:15:@64955.4]
  assign io_out_bits_wstrb_27 = io_in_bits_0_wstrb_27; // @[MuxN.scala 72:15:@64956.4]
  assign io_out_bits_wstrb_28 = io_in_bits_0_wstrb_28; // @[MuxN.scala 72:15:@64957.4]
  assign io_out_bits_wstrb_29 = io_in_bits_0_wstrb_29; // @[MuxN.scala 72:15:@64958.4]
  assign io_out_bits_wstrb_30 = io_in_bits_0_wstrb_30; // @[MuxN.scala 72:15:@64959.4]
  assign io_out_bits_wstrb_31 = io_in_bits_0_wstrb_31; // @[MuxN.scala 72:15:@64960.4]
  assign io_out_bits_wstrb_32 = io_in_bits_0_wstrb_32; // @[MuxN.scala 72:15:@64961.4]
  assign io_out_bits_wstrb_33 = io_in_bits_0_wstrb_33; // @[MuxN.scala 72:15:@64962.4]
  assign io_out_bits_wstrb_34 = io_in_bits_0_wstrb_34; // @[MuxN.scala 72:15:@64963.4]
  assign io_out_bits_wstrb_35 = io_in_bits_0_wstrb_35; // @[MuxN.scala 72:15:@64964.4]
  assign io_out_bits_wstrb_36 = io_in_bits_0_wstrb_36; // @[MuxN.scala 72:15:@64965.4]
  assign io_out_bits_wstrb_37 = io_in_bits_0_wstrb_37; // @[MuxN.scala 72:15:@64966.4]
  assign io_out_bits_wstrb_38 = io_in_bits_0_wstrb_38; // @[MuxN.scala 72:15:@64967.4]
  assign io_out_bits_wstrb_39 = io_in_bits_0_wstrb_39; // @[MuxN.scala 72:15:@64968.4]
  assign io_out_bits_wstrb_40 = io_in_bits_0_wstrb_40; // @[MuxN.scala 72:15:@64969.4]
  assign io_out_bits_wstrb_41 = io_in_bits_0_wstrb_41; // @[MuxN.scala 72:15:@64970.4]
  assign io_out_bits_wstrb_42 = io_in_bits_0_wstrb_42; // @[MuxN.scala 72:15:@64971.4]
  assign io_out_bits_wstrb_43 = io_in_bits_0_wstrb_43; // @[MuxN.scala 72:15:@64972.4]
  assign io_out_bits_wstrb_44 = io_in_bits_0_wstrb_44; // @[MuxN.scala 72:15:@64973.4]
  assign io_out_bits_wstrb_45 = io_in_bits_0_wstrb_45; // @[MuxN.scala 72:15:@64974.4]
  assign io_out_bits_wstrb_46 = io_in_bits_0_wstrb_46; // @[MuxN.scala 72:15:@64975.4]
  assign io_out_bits_wstrb_47 = io_in_bits_0_wstrb_47; // @[MuxN.scala 72:15:@64976.4]
  assign io_out_bits_wstrb_48 = io_in_bits_0_wstrb_48; // @[MuxN.scala 72:15:@64977.4]
  assign io_out_bits_wstrb_49 = io_in_bits_0_wstrb_49; // @[MuxN.scala 72:15:@64978.4]
  assign io_out_bits_wstrb_50 = io_in_bits_0_wstrb_50; // @[MuxN.scala 72:15:@64979.4]
  assign io_out_bits_wstrb_51 = io_in_bits_0_wstrb_51; // @[MuxN.scala 72:15:@64980.4]
  assign io_out_bits_wstrb_52 = io_in_bits_0_wstrb_52; // @[MuxN.scala 72:15:@64981.4]
  assign io_out_bits_wstrb_53 = io_in_bits_0_wstrb_53; // @[MuxN.scala 72:15:@64982.4]
  assign io_out_bits_wstrb_54 = io_in_bits_0_wstrb_54; // @[MuxN.scala 72:15:@64983.4]
  assign io_out_bits_wstrb_55 = io_in_bits_0_wstrb_55; // @[MuxN.scala 72:15:@64984.4]
  assign io_out_bits_wstrb_56 = io_in_bits_0_wstrb_56; // @[MuxN.scala 72:15:@64985.4]
  assign io_out_bits_wstrb_57 = io_in_bits_0_wstrb_57; // @[MuxN.scala 72:15:@64986.4]
  assign io_out_bits_wstrb_58 = io_in_bits_0_wstrb_58; // @[MuxN.scala 72:15:@64987.4]
  assign io_out_bits_wstrb_59 = io_in_bits_0_wstrb_59; // @[MuxN.scala 72:15:@64988.4]
  assign io_out_bits_wstrb_60 = io_in_bits_0_wstrb_60; // @[MuxN.scala 72:15:@64989.4]
  assign io_out_bits_wstrb_61 = io_in_bits_0_wstrb_61; // @[MuxN.scala 72:15:@64990.4]
  assign io_out_bits_wstrb_62 = io_in_bits_0_wstrb_62; // @[MuxN.scala 72:15:@64991.4]
  assign io_out_bits_wstrb_63 = io_in_bits_0_wstrb_63; // @[MuxN.scala 72:15:@64992.4]
endmodule
module ElementCounter( // @[:@65010.2]
  input         clock, // @[:@65011.4]
  input         reset, // @[:@65012.4]
  input         io_reset, // @[:@65013.4]
  input         io_enable, // @[:@65013.4]
  output [31:0] io_out // @[:@65013.4]
);
  reg [31:0] count; // @[Counter.scala 37:22:@65015.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_14; // @[Counter.scala 39:24:@65016.4]
  wire [31:0] newCount; // @[Counter.scala 39:24:@65017.4]
  wire [31:0] _GEN_0; // @[Counter.scala 43:26:@65022.6]
  wire [31:0] _GEN_1; // @[Counter.scala 41:18:@65018.4]
  assign _T_14 = count + 32'h1; // @[Counter.scala 39:24:@65016.4]
  assign newCount = count + 32'h1; // @[Counter.scala 39:24:@65017.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 43:26:@65022.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 41:18:@65018.4]
  assign io_out = count; // @[Counter.scala 47:10:@65025.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module StreamArbiter( // @[:@65027.2]
  input         clock, // @[:@65028.4]
  input         reset, // @[:@65029.4]
  output        io_app_0_cmd_ready, // @[:@65030.4]
  input         io_app_0_cmd_valid, // @[:@65030.4]
  input  [63:0] io_app_0_cmd_bits_addr, // @[:@65030.4]
  input  [31:0] io_app_0_cmd_bits_size, // @[:@65030.4]
  input         io_app_0_cmd_bits_isWr, // @[:@65030.4]
  input  [31:0] io_app_0_cmd_bits_tag, // @[:@65030.4]
  output        io_app_0_wdata_ready, // @[:@65030.4]
  input         io_app_0_wdata_valid, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_0, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_1, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_2, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_3, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_4, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_5, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_6, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_7, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_8, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_9, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_10, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_11, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_12, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_13, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_14, // @[:@65030.4]
  input  [31:0] io_app_0_wdata_bits_wdata_15, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_0, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_1, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_2, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_3, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_4, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_5, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_6, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_7, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_8, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_9, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_10, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_11, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_12, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_13, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_14, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_15, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_16, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_17, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_18, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_19, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_20, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_21, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_22, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_23, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_24, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_25, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_26, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_27, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_28, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_29, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_30, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_31, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_32, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_33, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_34, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_35, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_36, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_37, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_38, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_39, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_40, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_41, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_42, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_43, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_44, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_45, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_46, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_47, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_48, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_49, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_50, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_51, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_52, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_53, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_54, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_55, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_56, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_57, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_58, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_59, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_60, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_61, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_62, // @[:@65030.4]
  input         io_app_0_wdata_bits_wstrb_63, // @[:@65030.4]
  input         io_app_0_rresp_ready, // @[:@65030.4]
  input         io_app_0_wresp_ready, // @[:@65030.4]
  output        io_app_0_wresp_valid, // @[:@65030.4]
  input         io_dram_cmd_ready, // @[:@65030.4]
  output        io_dram_cmd_valid, // @[:@65030.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@65030.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@65030.4]
  output        io_dram_cmd_bits_isWr, // @[:@65030.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@65030.4]
  input         io_dram_wdata_ready, // @[:@65030.4]
  output        io_dram_wdata_valid, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@65030.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@65030.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@65030.4]
  output        io_dram_rresp_ready, // @[:@65030.4]
  output        io_dram_wresp_ready, // @[:@65030.4]
  input         io_dram_wresp_valid, // @[:@65030.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@65030.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@65259.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@65259.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@65259.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@65259.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@65259.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@65266.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@65266.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@65266.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@65266.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@65266.4]
  wire  cmdMux_io_in_ready; // @[StreamArbiter.scala 25:22:@65276.4]
  wire  cmdMux_io_in_valid; // @[StreamArbiter.scala 25:22:@65276.4]
  wire [63:0] cmdMux_io_in_bits_0_addr; // @[StreamArbiter.scala 25:22:@65276.4]
  wire [31:0] cmdMux_io_in_bits_0_size; // @[StreamArbiter.scala 25:22:@65276.4]
  wire  cmdMux_io_in_bits_0_isWr; // @[StreamArbiter.scala 25:22:@65276.4]
  wire [31:0] cmdMux_io_in_bits_0_tag; // @[StreamArbiter.scala 25:22:@65276.4]
  wire  cmdMux_io_out_ready; // @[StreamArbiter.scala 25:22:@65276.4]
  wire  cmdMux_io_out_valid; // @[StreamArbiter.scala 25:22:@65276.4]
  wire [63:0] cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 25:22:@65276.4]
  wire [31:0] cmdMux_io_out_bits_size; // @[StreamArbiter.scala 25:22:@65276.4]
  wire  cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 25:22:@65276.4]
  wire [31:0] cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 25:22:@65276.4]
  wire  wdataMux_io_in_ready; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_valid; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_0; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_1; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_2; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_3; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_4; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_5; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_6; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_7; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_8; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_9; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_10; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_11; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_12; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_13; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_14; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_15; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_0; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_1; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_2; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_3; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_4; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_5; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_6; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_7; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_8; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_9; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_10; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_11; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_12; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_13; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_14; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_15; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_16; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_17; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_18; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_19; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_20; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_21; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_22; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_23; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_24; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_25; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_26; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_27; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_28; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_29; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_30; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_31; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_32; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_33; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_34; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_35; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_36; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_37; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_38; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_39; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_40; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_41; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_42; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_43; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_44; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_45; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_46; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_47; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_48; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_49; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_50; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_51; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_52; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_53; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_54; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_55; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_56; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_57; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_58; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_59; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_60; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_61; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_62; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_in_bits_0_wstrb_63; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_ready; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_valid; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 35:24:@65299.4]
  wire [31:0] wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 35:24:@65299.4]
  wire  elementCtr_clock; // @[StreamArbiter.scala 36:26:@65302.4]
  wire  elementCtr_reset; // @[StreamArbiter.scala 36:26:@65302.4]
  wire  elementCtr_io_reset; // @[StreamArbiter.scala 36:26:@65302.4]
  wire  elementCtr_io_enable; // @[StreamArbiter.scala 36:26:@65302.4]
  wire [31:0] elementCtr_io_out; // @[StreamArbiter.scala 36:26:@65302.4]
  wire  _T_346; // @[package.scala 96:25:@65271.4 package.scala 96:25:@65272.4]
  wire  cmdIdx; // @[StreamArbiter.scala 21:16:@65273.4]
  wire [1:0] cmdInDecoder; // @[OneHot.scala 45:35:@65275.4]
  wire  _T_355; // @[FringeBundles.scala 114:28:@65291.4]
  wire [22:0] _T_356; // @[FringeBundles.scala 114:28:@65293.4]
  wire [23:0] _T_358; // @[FringeBundles.scala 115:37:@65296.4]
  wire  _T_360; // @[StreamArbiter.scala 37:49:@65305.4]
  wire [31:0] _T_365; // @[:@65309.4 :@65310.4]
  wire [7:0] _T_366; // @[FringeBundles.scala 114:28:@65311.4]
  wire [255:0] cmdOutDecoder; // @[OneHot.scala 45:35:@65317.4]
  wire  _T_379; // @[StreamArbiter.scala 42:78:@65320.4]
  wire  _T_380; // @[StreamArbiter.scala 42:121:@65321.4]
  wire [7:0] _T_395; // @[FringeBundles.scala 140:28:@65508.4]
  wire [255:0] wrespDecoder; // @[OneHot.scala 45:35:@65515.4]
  wire  _T_400; // @[StreamArbiter.scala 61:55:@65520.4]
  wire  _T_403; // @[StreamArbiter.scala 62:85:@65524.4]
  wire  _T_404; // @[StreamArbiter.scala 62:70:@65525.4]
  wire  _T_409; // @[StreamArbiter.scala 67:58:@65549.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@65259.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@65266.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  MuxPipe cmdMux ( // @[StreamArbiter.scala 25:22:@65276.4]
    .io_in_ready(cmdMux_io_in_ready),
    .io_in_valid(cmdMux_io_in_valid),
    .io_in_bits_0_addr(cmdMux_io_in_bits_0_addr),
    .io_in_bits_0_size(cmdMux_io_in_bits_0_size),
    .io_in_bits_0_isWr(cmdMux_io_in_bits_0_isWr),
    .io_in_bits_0_tag(cmdMux_io_in_bits_0_tag),
    .io_out_ready(cmdMux_io_out_ready),
    .io_out_valid(cmdMux_io_out_valid),
    .io_out_bits_addr(cmdMux_io_out_bits_addr),
    .io_out_bits_size(cmdMux_io_out_bits_size),
    .io_out_bits_isWr(cmdMux_io_out_bits_isWr),
    .io_out_bits_tag(cmdMux_io_out_bits_tag)
  );
  MuxPipe_1 wdataMux ( // @[StreamArbiter.scala 35:24:@65299.4]
    .io_in_ready(wdataMux_io_in_ready),
    .io_in_valid(wdataMux_io_in_valid),
    .io_in_bits_0_wdata_0(wdataMux_io_in_bits_0_wdata_0),
    .io_in_bits_0_wdata_1(wdataMux_io_in_bits_0_wdata_1),
    .io_in_bits_0_wdata_2(wdataMux_io_in_bits_0_wdata_2),
    .io_in_bits_0_wdata_3(wdataMux_io_in_bits_0_wdata_3),
    .io_in_bits_0_wdata_4(wdataMux_io_in_bits_0_wdata_4),
    .io_in_bits_0_wdata_5(wdataMux_io_in_bits_0_wdata_5),
    .io_in_bits_0_wdata_6(wdataMux_io_in_bits_0_wdata_6),
    .io_in_bits_0_wdata_7(wdataMux_io_in_bits_0_wdata_7),
    .io_in_bits_0_wdata_8(wdataMux_io_in_bits_0_wdata_8),
    .io_in_bits_0_wdata_9(wdataMux_io_in_bits_0_wdata_9),
    .io_in_bits_0_wdata_10(wdataMux_io_in_bits_0_wdata_10),
    .io_in_bits_0_wdata_11(wdataMux_io_in_bits_0_wdata_11),
    .io_in_bits_0_wdata_12(wdataMux_io_in_bits_0_wdata_12),
    .io_in_bits_0_wdata_13(wdataMux_io_in_bits_0_wdata_13),
    .io_in_bits_0_wdata_14(wdataMux_io_in_bits_0_wdata_14),
    .io_in_bits_0_wdata_15(wdataMux_io_in_bits_0_wdata_15),
    .io_in_bits_0_wstrb_0(wdataMux_io_in_bits_0_wstrb_0),
    .io_in_bits_0_wstrb_1(wdataMux_io_in_bits_0_wstrb_1),
    .io_in_bits_0_wstrb_2(wdataMux_io_in_bits_0_wstrb_2),
    .io_in_bits_0_wstrb_3(wdataMux_io_in_bits_0_wstrb_3),
    .io_in_bits_0_wstrb_4(wdataMux_io_in_bits_0_wstrb_4),
    .io_in_bits_0_wstrb_5(wdataMux_io_in_bits_0_wstrb_5),
    .io_in_bits_0_wstrb_6(wdataMux_io_in_bits_0_wstrb_6),
    .io_in_bits_0_wstrb_7(wdataMux_io_in_bits_0_wstrb_7),
    .io_in_bits_0_wstrb_8(wdataMux_io_in_bits_0_wstrb_8),
    .io_in_bits_0_wstrb_9(wdataMux_io_in_bits_0_wstrb_9),
    .io_in_bits_0_wstrb_10(wdataMux_io_in_bits_0_wstrb_10),
    .io_in_bits_0_wstrb_11(wdataMux_io_in_bits_0_wstrb_11),
    .io_in_bits_0_wstrb_12(wdataMux_io_in_bits_0_wstrb_12),
    .io_in_bits_0_wstrb_13(wdataMux_io_in_bits_0_wstrb_13),
    .io_in_bits_0_wstrb_14(wdataMux_io_in_bits_0_wstrb_14),
    .io_in_bits_0_wstrb_15(wdataMux_io_in_bits_0_wstrb_15),
    .io_in_bits_0_wstrb_16(wdataMux_io_in_bits_0_wstrb_16),
    .io_in_bits_0_wstrb_17(wdataMux_io_in_bits_0_wstrb_17),
    .io_in_bits_0_wstrb_18(wdataMux_io_in_bits_0_wstrb_18),
    .io_in_bits_0_wstrb_19(wdataMux_io_in_bits_0_wstrb_19),
    .io_in_bits_0_wstrb_20(wdataMux_io_in_bits_0_wstrb_20),
    .io_in_bits_0_wstrb_21(wdataMux_io_in_bits_0_wstrb_21),
    .io_in_bits_0_wstrb_22(wdataMux_io_in_bits_0_wstrb_22),
    .io_in_bits_0_wstrb_23(wdataMux_io_in_bits_0_wstrb_23),
    .io_in_bits_0_wstrb_24(wdataMux_io_in_bits_0_wstrb_24),
    .io_in_bits_0_wstrb_25(wdataMux_io_in_bits_0_wstrb_25),
    .io_in_bits_0_wstrb_26(wdataMux_io_in_bits_0_wstrb_26),
    .io_in_bits_0_wstrb_27(wdataMux_io_in_bits_0_wstrb_27),
    .io_in_bits_0_wstrb_28(wdataMux_io_in_bits_0_wstrb_28),
    .io_in_bits_0_wstrb_29(wdataMux_io_in_bits_0_wstrb_29),
    .io_in_bits_0_wstrb_30(wdataMux_io_in_bits_0_wstrb_30),
    .io_in_bits_0_wstrb_31(wdataMux_io_in_bits_0_wstrb_31),
    .io_in_bits_0_wstrb_32(wdataMux_io_in_bits_0_wstrb_32),
    .io_in_bits_0_wstrb_33(wdataMux_io_in_bits_0_wstrb_33),
    .io_in_bits_0_wstrb_34(wdataMux_io_in_bits_0_wstrb_34),
    .io_in_bits_0_wstrb_35(wdataMux_io_in_bits_0_wstrb_35),
    .io_in_bits_0_wstrb_36(wdataMux_io_in_bits_0_wstrb_36),
    .io_in_bits_0_wstrb_37(wdataMux_io_in_bits_0_wstrb_37),
    .io_in_bits_0_wstrb_38(wdataMux_io_in_bits_0_wstrb_38),
    .io_in_bits_0_wstrb_39(wdataMux_io_in_bits_0_wstrb_39),
    .io_in_bits_0_wstrb_40(wdataMux_io_in_bits_0_wstrb_40),
    .io_in_bits_0_wstrb_41(wdataMux_io_in_bits_0_wstrb_41),
    .io_in_bits_0_wstrb_42(wdataMux_io_in_bits_0_wstrb_42),
    .io_in_bits_0_wstrb_43(wdataMux_io_in_bits_0_wstrb_43),
    .io_in_bits_0_wstrb_44(wdataMux_io_in_bits_0_wstrb_44),
    .io_in_bits_0_wstrb_45(wdataMux_io_in_bits_0_wstrb_45),
    .io_in_bits_0_wstrb_46(wdataMux_io_in_bits_0_wstrb_46),
    .io_in_bits_0_wstrb_47(wdataMux_io_in_bits_0_wstrb_47),
    .io_in_bits_0_wstrb_48(wdataMux_io_in_bits_0_wstrb_48),
    .io_in_bits_0_wstrb_49(wdataMux_io_in_bits_0_wstrb_49),
    .io_in_bits_0_wstrb_50(wdataMux_io_in_bits_0_wstrb_50),
    .io_in_bits_0_wstrb_51(wdataMux_io_in_bits_0_wstrb_51),
    .io_in_bits_0_wstrb_52(wdataMux_io_in_bits_0_wstrb_52),
    .io_in_bits_0_wstrb_53(wdataMux_io_in_bits_0_wstrb_53),
    .io_in_bits_0_wstrb_54(wdataMux_io_in_bits_0_wstrb_54),
    .io_in_bits_0_wstrb_55(wdataMux_io_in_bits_0_wstrb_55),
    .io_in_bits_0_wstrb_56(wdataMux_io_in_bits_0_wstrb_56),
    .io_in_bits_0_wstrb_57(wdataMux_io_in_bits_0_wstrb_57),
    .io_in_bits_0_wstrb_58(wdataMux_io_in_bits_0_wstrb_58),
    .io_in_bits_0_wstrb_59(wdataMux_io_in_bits_0_wstrb_59),
    .io_in_bits_0_wstrb_60(wdataMux_io_in_bits_0_wstrb_60),
    .io_in_bits_0_wstrb_61(wdataMux_io_in_bits_0_wstrb_61),
    .io_in_bits_0_wstrb_62(wdataMux_io_in_bits_0_wstrb_62),
    .io_in_bits_0_wstrb_63(wdataMux_io_in_bits_0_wstrb_63),
    .io_out_ready(wdataMux_io_out_ready),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  ElementCounter elementCtr ( // @[StreamArbiter.scala 36:26:@65302.4]
    .clock(elementCtr_clock),
    .reset(elementCtr_reset),
    .io_reset(elementCtr_io_reset),
    .io_enable(elementCtr_io_enable),
    .io_out(elementCtr_io_out)
  );
  assign _T_346 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@65271.4 package.scala 96:25:@65272.4]
  assign cmdIdx = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[StreamArbiter.scala 21:16:@65273.4]
  assign cmdInDecoder = 2'h1 << cmdIdx; // @[OneHot.scala 45:35:@65275.4]
  assign _T_355 = io_app_0_cmd_bits_tag[8]; // @[FringeBundles.scala 114:28:@65291.4]
  assign _T_356 = io_app_0_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@65293.4]
  assign _T_358 = {_T_356,_T_355}; // @[FringeBundles.scala 115:37:@65296.4]
  assign _T_360 = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:49:@65305.4]
  assign _T_365 = cmdMux_io_out_bits_tag; // @[:@65309.4 :@65310.4]
  assign _T_366 = _T_365[7:0]; // @[FringeBundles.scala 114:28:@65311.4]
  assign cmdOutDecoder = 256'h1 << _T_366; // @[OneHot.scala 45:35:@65317.4]
  assign _T_379 = io_app_0_wdata_valid & cmdMux_io_out_valid; // @[StreamArbiter.scala 42:78:@65320.4]
  assign _T_380 = elementCtr_io_out < cmdMux_io_out_bits_size; // @[StreamArbiter.scala 42:121:@65321.4]
  assign _T_395 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@65508.4]
  assign wrespDecoder = 256'h1 << _T_395; // @[OneHot.scala 45:35:@65515.4]
  assign _T_400 = cmdInDecoder[0]; // @[StreamArbiter.scala 61:55:@65520.4]
  assign _T_403 = cmdOutDecoder[0]; // @[StreamArbiter.scala 62:85:@65524.4]
  assign _T_404 = _T_360 & _T_403; // @[StreamArbiter.scala 62:70:@65525.4]
  assign _T_409 = wrespDecoder[0]; // @[StreamArbiter.scala 67:58:@65549.4]
  assign io_app_0_cmd_ready = cmdMux_io_in_ready & _T_400; // @[StreamArbiter.scala 61:19:@65522.4]
  assign io_app_0_wdata_ready = _T_404 & _T_380; // @[StreamArbiter.scala 62:21:@65528.4]
  assign io_app_0_wresp_valid = io_dram_wresp_valid & _T_409; // @[StreamArbiter.scala 67:21:@65551.4]
  assign io_dram_cmd_valid = cmdMux_io_out_valid; // @[StreamArbiter.scala 46:15:@65411.4]
  assign io_dram_cmd_bits_addr = cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 46:15:@65410.4]
  assign io_dram_cmd_bits_size = cmdMux_io_out_bits_size; // @[StreamArbiter.scala 46:15:@65409.4]
  assign io_dram_cmd_bits_isWr = cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 46:15:@65407.4]
  assign io_dram_cmd_bits_tag = cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 46:15:@65406.4]
  assign io_dram_wdata_valid = wdataMux_io_out_valid; // @[StreamArbiter.scala 47:17:@65494.4]
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 47:17:@65478.4]
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 47:17:@65479.4]
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 47:17:@65480.4]
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 47:17:@65481.4]
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 47:17:@65482.4]
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 47:17:@65483.4]
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 47:17:@65484.4]
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 47:17:@65485.4]
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 47:17:@65486.4]
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 47:17:@65487.4]
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 47:17:@65488.4]
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 47:17:@65489.4]
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 47:17:@65490.4]
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 47:17:@65491.4]
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 47:17:@65492.4]
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 47:17:@65493.4]
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 47:17:@65414.4]
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 47:17:@65415.4]
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 47:17:@65416.4]
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 47:17:@65417.4]
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 47:17:@65418.4]
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 47:17:@65419.4]
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 47:17:@65420.4]
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 47:17:@65421.4]
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 47:17:@65422.4]
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 47:17:@65423.4]
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 47:17:@65424.4]
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 47:17:@65425.4]
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 47:17:@65426.4]
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 47:17:@65427.4]
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 47:17:@65428.4]
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 47:17:@65429.4]
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 47:17:@65430.4]
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 47:17:@65431.4]
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 47:17:@65432.4]
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 47:17:@65433.4]
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 47:17:@65434.4]
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 47:17:@65435.4]
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 47:17:@65436.4]
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 47:17:@65437.4]
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 47:17:@65438.4]
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 47:17:@65439.4]
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 47:17:@65440.4]
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 47:17:@65441.4]
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 47:17:@65442.4]
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 47:17:@65443.4]
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 47:17:@65444.4]
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 47:17:@65445.4]
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 47:17:@65446.4]
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 47:17:@65447.4]
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 47:17:@65448.4]
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 47:17:@65449.4]
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 47:17:@65450.4]
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 47:17:@65451.4]
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 47:17:@65452.4]
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 47:17:@65453.4]
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 47:17:@65454.4]
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 47:17:@65455.4]
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 47:17:@65456.4]
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 47:17:@65457.4]
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 47:17:@65458.4]
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 47:17:@65459.4]
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 47:17:@65460.4]
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 47:17:@65461.4]
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 47:17:@65462.4]
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 47:17:@65463.4]
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 47:17:@65464.4]
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 47:17:@65465.4]
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 47:17:@65466.4]
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 47:17:@65467.4]
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 47:17:@65468.4]
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 47:17:@65469.4]
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 47:17:@65470.4]
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 47:17:@65471.4]
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 47:17:@65472.4]
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 47:17:@65473.4]
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 47:17:@65474.4]
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 47:17:@65475.4]
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 47:17:@65476.4]
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 47:17:@65477.4]
  assign io_dram_rresp_ready = io_app_0_rresp_ready; // @[StreamArbiter.scala 72:23:@65555.4]
  assign io_dram_wresp_ready = io_app_0_wresp_ready; // @[StreamArbiter.scala 73:23:@65558.4]
  assign RetimeWrapper_clock = clock; // @[:@65260.4]
  assign RetimeWrapper_reset = reset; // @[:@65261.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@65263.4]
  assign RetimeWrapper_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@65262.4]
  assign RetimeWrapper_1_clock = clock; // @[:@65267.4]
  assign RetimeWrapper_1_reset = reset; // @[:@65268.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@65270.4]
  assign RetimeWrapper_1_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@65269.4]
  assign cmdMux_io_in_valid = io_app_0_cmd_valid; // @[StreamArbiter.scala 26:22:@65279.4]
  assign cmdMux_io_in_bits_0_addr = io_app_0_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@65285.4]
  assign cmdMux_io_in_bits_0_size = io_app_0_cmd_bits_size; // @[StreamArbiter.scala 29:9:@65284.4]
  assign cmdMux_io_in_bits_0_isWr = io_app_0_cmd_bits_isWr; // @[StreamArbiter.scala 29:9:@65282.4]
  assign cmdMux_io_in_bits_0_tag = {_T_358,8'h0}; // @[StreamArbiter.scala 29:9:@65281.4 FringeBundles.scala 115:32:@65298.4]
  assign cmdMux_io_out_ready = io_dram_cmd_valid & io_dram_cmd_ready; // @[StreamArbiter.scala 46:15:@65412.4 StreamArbiter.scala 57:23:@65518.4]
  assign wdataMux_io_in_valid = _T_379 & _T_380; // @[StreamArbiter.scala 42:24:@65323.4]
  assign wdataMux_io_in_bits_0_wdata_0 = io_app_0_wdata_bits_wdata_0; // @[StreamArbiter.scala 44:23:@65390.4]
  assign wdataMux_io_in_bits_0_wdata_1 = io_app_0_wdata_bits_wdata_1; // @[StreamArbiter.scala 44:23:@65391.4]
  assign wdataMux_io_in_bits_0_wdata_2 = io_app_0_wdata_bits_wdata_2; // @[StreamArbiter.scala 44:23:@65392.4]
  assign wdataMux_io_in_bits_0_wdata_3 = io_app_0_wdata_bits_wdata_3; // @[StreamArbiter.scala 44:23:@65393.4]
  assign wdataMux_io_in_bits_0_wdata_4 = io_app_0_wdata_bits_wdata_4; // @[StreamArbiter.scala 44:23:@65394.4]
  assign wdataMux_io_in_bits_0_wdata_5 = io_app_0_wdata_bits_wdata_5; // @[StreamArbiter.scala 44:23:@65395.4]
  assign wdataMux_io_in_bits_0_wdata_6 = io_app_0_wdata_bits_wdata_6; // @[StreamArbiter.scala 44:23:@65396.4]
  assign wdataMux_io_in_bits_0_wdata_7 = io_app_0_wdata_bits_wdata_7; // @[StreamArbiter.scala 44:23:@65397.4]
  assign wdataMux_io_in_bits_0_wdata_8 = io_app_0_wdata_bits_wdata_8; // @[StreamArbiter.scala 44:23:@65398.4]
  assign wdataMux_io_in_bits_0_wdata_9 = io_app_0_wdata_bits_wdata_9; // @[StreamArbiter.scala 44:23:@65399.4]
  assign wdataMux_io_in_bits_0_wdata_10 = io_app_0_wdata_bits_wdata_10; // @[StreamArbiter.scala 44:23:@65400.4]
  assign wdataMux_io_in_bits_0_wdata_11 = io_app_0_wdata_bits_wdata_11; // @[StreamArbiter.scala 44:23:@65401.4]
  assign wdataMux_io_in_bits_0_wdata_12 = io_app_0_wdata_bits_wdata_12; // @[StreamArbiter.scala 44:23:@65402.4]
  assign wdataMux_io_in_bits_0_wdata_13 = io_app_0_wdata_bits_wdata_13; // @[StreamArbiter.scala 44:23:@65403.4]
  assign wdataMux_io_in_bits_0_wdata_14 = io_app_0_wdata_bits_wdata_14; // @[StreamArbiter.scala 44:23:@65404.4]
  assign wdataMux_io_in_bits_0_wdata_15 = io_app_0_wdata_bits_wdata_15; // @[StreamArbiter.scala 44:23:@65405.4]
  assign wdataMux_io_in_bits_0_wstrb_0 = io_app_0_wdata_bits_wstrb_0; // @[StreamArbiter.scala 44:23:@65326.4]
  assign wdataMux_io_in_bits_0_wstrb_1 = io_app_0_wdata_bits_wstrb_1; // @[StreamArbiter.scala 44:23:@65327.4]
  assign wdataMux_io_in_bits_0_wstrb_2 = io_app_0_wdata_bits_wstrb_2; // @[StreamArbiter.scala 44:23:@65328.4]
  assign wdataMux_io_in_bits_0_wstrb_3 = io_app_0_wdata_bits_wstrb_3; // @[StreamArbiter.scala 44:23:@65329.4]
  assign wdataMux_io_in_bits_0_wstrb_4 = io_app_0_wdata_bits_wstrb_4; // @[StreamArbiter.scala 44:23:@65330.4]
  assign wdataMux_io_in_bits_0_wstrb_5 = io_app_0_wdata_bits_wstrb_5; // @[StreamArbiter.scala 44:23:@65331.4]
  assign wdataMux_io_in_bits_0_wstrb_6 = io_app_0_wdata_bits_wstrb_6; // @[StreamArbiter.scala 44:23:@65332.4]
  assign wdataMux_io_in_bits_0_wstrb_7 = io_app_0_wdata_bits_wstrb_7; // @[StreamArbiter.scala 44:23:@65333.4]
  assign wdataMux_io_in_bits_0_wstrb_8 = io_app_0_wdata_bits_wstrb_8; // @[StreamArbiter.scala 44:23:@65334.4]
  assign wdataMux_io_in_bits_0_wstrb_9 = io_app_0_wdata_bits_wstrb_9; // @[StreamArbiter.scala 44:23:@65335.4]
  assign wdataMux_io_in_bits_0_wstrb_10 = io_app_0_wdata_bits_wstrb_10; // @[StreamArbiter.scala 44:23:@65336.4]
  assign wdataMux_io_in_bits_0_wstrb_11 = io_app_0_wdata_bits_wstrb_11; // @[StreamArbiter.scala 44:23:@65337.4]
  assign wdataMux_io_in_bits_0_wstrb_12 = io_app_0_wdata_bits_wstrb_12; // @[StreamArbiter.scala 44:23:@65338.4]
  assign wdataMux_io_in_bits_0_wstrb_13 = io_app_0_wdata_bits_wstrb_13; // @[StreamArbiter.scala 44:23:@65339.4]
  assign wdataMux_io_in_bits_0_wstrb_14 = io_app_0_wdata_bits_wstrb_14; // @[StreamArbiter.scala 44:23:@65340.4]
  assign wdataMux_io_in_bits_0_wstrb_15 = io_app_0_wdata_bits_wstrb_15; // @[StreamArbiter.scala 44:23:@65341.4]
  assign wdataMux_io_in_bits_0_wstrb_16 = io_app_0_wdata_bits_wstrb_16; // @[StreamArbiter.scala 44:23:@65342.4]
  assign wdataMux_io_in_bits_0_wstrb_17 = io_app_0_wdata_bits_wstrb_17; // @[StreamArbiter.scala 44:23:@65343.4]
  assign wdataMux_io_in_bits_0_wstrb_18 = io_app_0_wdata_bits_wstrb_18; // @[StreamArbiter.scala 44:23:@65344.4]
  assign wdataMux_io_in_bits_0_wstrb_19 = io_app_0_wdata_bits_wstrb_19; // @[StreamArbiter.scala 44:23:@65345.4]
  assign wdataMux_io_in_bits_0_wstrb_20 = io_app_0_wdata_bits_wstrb_20; // @[StreamArbiter.scala 44:23:@65346.4]
  assign wdataMux_io_in_bits_0_wstrb_21 = io_app_0_wdata_bits_wstrb_21; // @[StreamArbiter.scala 44:23:@65347.4]
  assign wdataMux_io_in_bits_0_wstrb_22 = io_app_0_wdata_bits_wstrb_22; // @[StreamArbiter.scala 44:23:@65348.4]
  assign wdataMux_io_in_bits_0_wstrb_23 = io_app_0_wdata_bits_wstrb_23; // @[StreamArbiter.scala 44:23:@65349.4]
  assign wdataMux_io_in_bits_0_wstrb_24 = io_app_0_wdata_bits_wstrb_24; // @[StreamArbiter.scala 44:23:@65350.4]
  assign wdataMux_io_in_bits_0_wstrb_25 = io_app_0_wdata_bits_wstrb_25; // @[StreamArbiter.scala 44:23:@65351.4]
  assign wdataMux_io_in_bits_0_wstrb_26 = io_app_0_wdata_bits_wstrb_26; // @[StreamArbiter.scala 44:23:@65352.4]
  assign wdataMux_io_in_bits_0_wstrb_27 = io_app_0_wdata_bits_wstrb_27; // @[StreamArbiter.scala 44:23:@65353.4]
  assign wdataMux_io_in_bits_0_wstrb_28 = io_app_0_wdata_bits_wstrb_28; // @[StreamArbiter.scala 44:23:@65354.4]
  assign wdataMux_io_in_bits_0_wstrb_29 = io_app_0_wdata_bits_wstrb_29; // @[StreamArbiter.scala 44:23:@65355.4]
  assign wdataMux_io_in_bits_0_wstrb_30 = io_app_0_wdata_bits_wstrb_30; // @[StreamArbiter.scala 44:23:@65356.4]
  assign wdataMux_io_in_bits_0_wstrb_31 = io_app_0_wdata_bits_wstrb_31; // @[StreamArbiter.scala 44:23:@65357.4]
  assign wdataMux_io_in_bits_0_wstrb_32 = io_app_0_wdata_bits_wstrb_32; // @[StreamArbiter.scala 44:23:@65358.4]
  assign wdataMux_io_in_bits_0_wstrb_33 = io_app_0_wdata_bits_wstrb_33; // @[StreamArbiter.scala 44:23:@65359.4]
  assign wdataMux_io_in_bits_0_wstrb_34 = io_app_0_wdata_bits_wstrb_34; // @[StreamArbiter.scala 44:23:@65360.4]
  assign wdataMux_io_in_bits_0_wstrb_35 = io_app_0_wdata_bits_wstrb_35; // @[StreamArbiter.scala 44:23:@65361.4]
  assign wdataMux_io_in_bits_0_wstrb_36 = io_app_0_wdata_bits_wstrb_36; // @[StreamArbiter.scala 44:23:@65362.4]
  assign wdataMux_io_in_bits_0_wstrb_37 = io_app_0_wdata_bits_wstrb_37; // @[StreamArbiter.scala 44:23:@65363.4]
  assign wdataMux_io_in_bits_0_wstrb_38 = io_app_0_wdata_bits_wstrb_38; // @[StreamArbiter.scala 44:23:@65364.4]
  assign wdataMux_io_in_bits_0_wstrb_39 = io_app_0_wdata_bits_wstrb_39; // @[StreamArbiter.scala 44:23:@65365.4]
  assign wdataMux_io_in_bits_0_wstrb_40 = io_app_0_wdata_bits_wstrb_40; // @[StreamArbiter.scala 44:23:@65366.4]
  assign wdataMux_io_in_bits_0_wstrb_41 = io_app_0_wdata_bits_wstrb_41; // @[StreamArbiter.scala 44:23:@65367.4]
  assign wdataMux_io_in_bits_0_wstrb_42 = io_app_0_wdata_bits_wstrb_42; // @[StreamArbiter.scala 44:23:@65368.4]
  assign wdataMux_io_in_bits_0_wstrb_43 = io_app_0_wdata_bits_wstrb_43; // @[StreamArbiter.scala 44:23:@65369.4]
  assign wdataMux_io_in_bits_0_wstrb_44 = io_app_0_wdata_bits_wstrb_44; // @[StreamArbiter.scala 44:23:@65370.4]
  assign wdataMux_io_in_bits_0_wstrb_45 = io_app_0_wdata_bits_wstrb_45; // @[StreamArbiter.scala 44:23:@65371.4]
  assign wdataMux_io_in_bits_0_wstrb_46 = io_app_0_wdata_bits_wstrb_46; // @[StreamArbiter.scala 44:23:@65372.4]
  assign wdataMux_io_in_bits_0_wstrb_47 = io_app_0_wdata_bits_wstrb_47; // @[StreamArbiter.scala 44:23:@65373.4]
  assign wdataMux_io_in_bits_0_wstrb_48 = io_app_0_wdata_bits_wstrb_48; // @[StreamArbiter.scala 44:23:@65374.4]
  assign wdataMux_io_in_bits_0_wstrb_49 = io_app_0_wdata_bits_wstrb_49; // @[StreamArbiter.scala 44:23:@65375.4]
  assign wdataMux_io_in_bits_0_wstrb_50 = io_app_0_wdata_bits_wstrb_50; // @[StreamArbiter.scala 44:23:@65376.4]
  assign wdataMux_io_in_bits_0_wstrb_51 = io_app_0_wdata_bits_wstrb_51; // @[StreamArbiter.scala 44:23:@65377.4]
  assign wdataMux_io_in_bits_0_wstrb_52 = io_app_0_wdata_bits_wstrb_52; // @[StreamArbiter.scala 44:23:@65378.4]
  assign wdataMux_io_in_bits_0_wstrb_53 = io_app_0_wdata_bits_wstrb_53; // @[StreamArbiter.scala 44:23:@65379.4]
  assign wdataMux_io_in_bits_0_wstrb_54 = io_app_0_wdata_bits_wstrb_54; // @[StreamArbiter.scala 44:23:@65380.4]
  assign wdataMux_io_in_bits_0_wstrb_55 = io_app_0_wdata_bits_wstrb_55; // @[StreamArbiter.scala 44:23:@65381.4]
  assign wdataMux_io_in_bits_0_wstrb_56 = io_app_0_wdata_bits_wstrb_56; // @[StreamArbiter.scala 44:23:@65382.4]
  assign wdataMux_io_in_bits_0_wstrb_57 = io_app_0_wdata_bits_wstrb_57; // @[StreamArbiter.scala 44:23:@65383.4]
  assign wdataMux_io_in_bits_0_wstrb_58 = io_app_0_wdata_bits_wstrb_58; // @[StreamArbiter.scala 44:23:@65384.4]
  assign wdataMux_io_in_bits_0_wstrb_59 = io_app_0_wdata_bits_wstrb_59; // @[StreamArbiter.scala 44:23:@65385.4]
  assign wdataMux_io_in_bits_0_wstrb_60 = io_app_0_wdata_bits_wstrb_60; // @[StreamArbiter.scala 44:23:@65386.4]
  assign wdataMux_io_in_bits_0_wstrb_61 = io_app_0_wdata_bits_wstrb_61; // @[StreamArbiter.scala 44:23:@65387.4]
  assign wdataMux_io_in_bits_0_wstrb_62 = io_app_0_wdata_bits_wstrb_62; // @[StreamArbiter.scala 44:23:@65388.4]
  assign wdataMux_io_in_bits_0_wstrb_63 = io_app_0_wdata_bits_wstrb_63; // @[StreamArbiter.scala 44:23:@65389.4]
  assign wdataMux_io_out_ready = io_dram_wdata_valid & io_dram_wdata_ready; // @[StreamArbiter.scala 47:17:@65495.4 StreamArbiter.scala 58:25:@65519.4]
  assign elementCtr_clock = clock; // @[:@65303.4]
  assign elementCtr_reset = reset; // @[:@65304.4]
  assign elementCtr_io_reset = cmdMux_io_out_ready; // @[StreamArbiter.scala 38:23:@65307.4]
  assign elementCtr_io_enable = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:24:@65306.4]
endmodule
module Counter_72( // @[:@65560.2]
  input         clock, // @[:@65561.4]
  input         reset, // @[:@65562.4]
  input         io_reset, // @[:@65563.4]
  input         io_enable, // @[:@65563.4]
  input  [31:0] io_stride, // @[:@65563.4]
  output [31:0] io_out, // @[:@65563.4]
  output [31:0] io_next // @[:@65563.4]
);
  reg [31:0] count; // @[Counter.scala 15:22:@65565.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_17; // @[Counter.scala 17:24:@65566.4]
  wire [31:0] newCount; // @[Counter.scala 17:24:@65567.4]
  wire [31:0] _GEN_0; // @[Counter.scala 21:26:@65572.6]
  wire [31:0] _GEN_1; // @[Counter.scala 19:18:@65568.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@65566.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@65567.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@65572.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 19:18:@65568.4]
  assign io_out = count; // @[Counter.scala 25:10:@65575.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@65576.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module AXICmdSplit( // @[:@65578.2]
  input         clock, // @[:@65579.4]
  input         reset, // @[:@65580.4]
  output        io_in_cmd_ready, // @[:@65581.4]
  input         io_in_cmd_valid, // @[:@65581.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@65581.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@65581.4]
  input         io_in_cmd_bits_isWr, // @[:@65581.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@65581.4]
  output        io_in_wdata_ready, // @[:@65581.4]
  input         io_in_wdata_valid, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@65581.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@65581.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@65581.4]
  input         io_in_rresp_ready, // @[:@65581.4]
  input         io_in_wresp_ready, // @[:@65581.4]
  output        io_in_wresp_valid, // @[:@65581.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@65581.4]
  input         io_out_cmd_ready, // @[:@65581.4]
  output        io_out_cmd_valid, // @[:@65581.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@65581.4]
  output [31:0] io_out_cmd_bits_size, // @[:@65581.4]
  output        io_out_cmd_bits_isWr, // @[:@65581.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@65581.4]
  input         io_out_wdata_ready, // @[:@65581.4]
  output        io_out_wdata_valid, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@65581.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@65581.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@65581.4]
  output        io_out_rresp_ready, // @[:@65581.4]
  output        io_out_wresp_ready, // @[:@65581.4]
  input         io_out_wresp_valid, // @[:@65581.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@65581.4]
);
  wire  cmdSizeCounter_clock; // @[AXIProtocol.scala 18:30:@65695.4]
  wire  cmdSizeCounter_reset; // @[AXIProtocol.scala 18:30:@65695.4]
  wire  cmdSizeCounter_io_reset; // @[AXIProtocol.scala 18:30:@65695.4]
  wire  cmdSizeCounter_io_enable; // @[AXIProtocol.scala 18:30:@65695.4]
  wire [31:0] cmdSizeCounter_io_stride; // @[AXIProtocol.scala 18:30:@65695.4]
  wire [31:0] cmdSizeCounter_io_out; // @[AXIProtocol.scala 18:30:@65695.4]
  wire [31:0] cmdSizeCounter_io_next; // @[AXIProtocol.scala 18:30:@65695.4]
  wire [32:0] _T_199; // @[AXIProtocol.scala 20:46:@65698.4]
  wire [32:0] _T_200; // @[AXIProtocol.scala 20:46:@65699.4]
  wire [31:0] cmdSizeRemaining; // @[AXIProtocol.scala 20:46:@65700.4]
  wire  lastCmd; // @[AXIProtocol.scala 23:35:@65701.4]
  wire [37:0] _GEN_0; // @[AXIProtocol.scala 27:47:@65704.4]
  wire [37:0] addrOffsetBytes; // @[AXIProtocol.scala 27:47:@65704.4]
  wire [63:0] _GEN_1; // @[AXIProtocol.scala 28:49:@65705.4]
  wire [64:0] _T_201; // @[AXIProtocol.scala 28:49:@65705.4]
  wire [63:0] cmdAddr_bits; // @[AXIProtocol.scala 28:49:@65706.4]
  wire [57:0] _T_204; // @[FringeBundles.scala 158:22:@65709.4]
  wire [7:0] cmdTag_streamID; // @[FringeBundles.scala 114:28:@65716.4]
  wire [22:0] cmdTag_uid; // @[FringeBundles.scala 114:28:@65720.4]
  wire [23:0] _T_214; // @[FringeBundles.scala 115:37:@65723.4]
  wire  cmdIssue; // @[AXIProtocol.scala 36:35:@65726.4]
  wire  _T_223; // @[FringeBundles.scala 140:28:@65737.4]
  Counter_72 cmdSizeCounter ( // @[AXIProtocol.scala 18:30:@65695.4]
    .clock(cmdSizeCounter_clock),
    .reset(cmdSizeCounter_reset),
    .io_reset(cmdSizeCounter_io_reset),
    .io_enable(cmdSizeCounter_io_enable),
    .io_stride(cmdSizeCounter_io_stride),
    .io_out(cmdSizeCounter_io_out),
    .io_next(cmdSizeCounter_io_next)
  );
  assign _T_199 = io_in_cmd_bits_size - cmdSizeCounter_io_out; // @[AXIProtocol.scala 20:46:@65698.4]
  assign _T_200 = $unsigned(_T_199); // @[AXIProtocol.scala 20:46:@65699.4]
  assign cmdSizeRemaining = _T_200[31:0]; // @[AXIProtocol.scala 20:46:@65700.4]
  assign lastCmd = cmdSizeRemaining <= 32'h100; // @[AXIProtocol.scala 23:35:@65701.4]
  assign _GEN_0 = {{6'd0}, cmdSizeCounter_io_out}; // @[AXIProtocol.scala 27:47:@65704.4]
  assign addrOffsetBytes = _GEN_0 << 6; // @[AXIProtocol.scala 27:47:@65704.4]
  assign _GEN_1 = {{26'd0}, addrOffsetBytes}; // @[AXIProtocol.scala 28:49:@65705.4]
  assign _T_201 = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@65705.4]
  assign cmdAddr_bits = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@65706.4]
  assign _T_204 = cmdAddr_bits[63:6]; // @[FringeBundles.scala 158:22:@65709.4]
  assign cmdTag_streamID = io_in_cmd_bits_tag[7:0]; // @[FringeBundles.scala 114:28:@65716.4]
  assign cmdTag_uid = io_in_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@65720.4]
  assign _T_214 = {cmdTag_uid,lastCmd}; // @[FringeBundles.scala 115:37:@65723.4]
  assign cmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 36:35:@65726.4]
  assign _T_223 = io_out_wresp_bits_tag[8]; // @[FringeBundles.scala 140:28:@65737.4]
  assign io_in_cmd_ready = lastCmd & cmdIssue; // @[AXIProtocol.scala 15:10:@65694.4 AXIProtocol.scala 38:19:@65728.4]
  assign io_in_wdata_ready = io_out_wdata_ready; // @[AXIProtocol.scala 15:10:@65687.4]
  assign io_in_wresp_valid = io_out_wresp_valid & _T_223; // @[AXIProtocol.scala 15:10:@65584.4 AXIProtocol.scala 46:21:@65742.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 15:10:@65583.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 15:10:@65693.4]
  assign io_out_cmd_bits_addr = {_T_204,6'h0}; // @[AXIProtocol.scala 15:10:@65692.4 AXIProtocol.scala 29:24:@65711.4]
  assign io_out_cmd_bits_size = lastCmd ? cmdSizeRemaining : 32'h100; // @[AXIProtocol.scala 15:10:@65691.4 AXIProtocol.scala 25:24:@65703.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 15:10:@65689.4]
  assign io_out_cmd_bits_tag = {_T_214,cmdTag_streamID}; // @[AXIProtocol.scala 15:10:@65688.4 FringeBundles.scala 115:32:@65725.4]
  assign io_out_wdata_valid = io_in_wdata_valid; // @[AXIProtocol.scala 15:10:@65686.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 15:10:@65670.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 15:10:@65671.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 15:10:@65672.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 15:10:@65673.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 15:10:@65674.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 15:10:@65675.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 15:10:@65676.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 15:10:@65677.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 15:10:@65678.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 15:10:@65679.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 15:10:@65680.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 15:10:@65681.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 15:10:@65682.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 15:10:@65683.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 15:10:@65684.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 15:10:@65685.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 15:10:@65606.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 15:10:@65607.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 15:10:@65608.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 15:10:@65609.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 15:10:@65610.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 15:10:@65611.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 15:10:@65612.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 15:10:@65613.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 15:10:@65614.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 15:10:@65615.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 15:10:@65616.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 15:10:@65617.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 15:10:@65618.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 15:10:@65619.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 15:10:@65620.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 15:10:@65621.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 15:10:@65622.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 15:10:@65623.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 15:10:@65624.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 15:10:@65625.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 15:10:@65626.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 15:10:@65627.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 15:10:@65628.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 15:10:@65629.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 15:10:@65630.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 15:10:@65631.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 15:10:@65632.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 15:10:@65633.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 15:10:@65634.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 15:10:@65635.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 15:10:@65636.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 15:10:@65637.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 15:10:@65638.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 15:10:@65639.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 15:10:@65640.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 15:10:@65641.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 15:10:@65642.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 15:10:@65643.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 15:10:@65644.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 15:10:@65645.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 15:10:@65646.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 15:10:@65647.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 15:10:@65648.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 15:10:@65649.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 15:10:@65650.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 15:10:@65651.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 15:10:@65652.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 15:10:@65653.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 15:10:@65654.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 15:10:@65655.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 15:10:@65656.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 15:10:@65657.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 15:10:@65658.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 15:10:@65659.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 15:10:@65660.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 15:10:@65661.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 15:10:@65662.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 15:10:@65663.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 15:10:@65664.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 15:10:@65665.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 15:10:@65666.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 15:10:@65667.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 15:10:@65668.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 15:10:@65669.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 15:10:@65604.4]
  assign io_out_wresp_ready = _T_223 ? io_in_wresp_ready : 1'h1; // @[AXIProtocol.scala 15:10:@65585.4 AXIProtocol.scala 47:22:@65744.4]
  assign cmdSizeCounter_clock = clock; // @[:@65696.4]
  assign cmdSizeCounter_reset = reset; // @[:@65697.4]
  assign cmdSizeCounter_io_reset = lastCmd & cmdIssue; // @[AXIProtocol.scala 40:27:@65729.4]
  assign cmdSizeCounter_io_enable = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 41:28:@65730.4]
  assign cmdSizeCounter_io_stride = 32'h100; // @[AXIProtocol.scala 42:28:@65731.4]
endmodule
module AXICmdIssue( // @[:@65764.2]
  input         clock, // @[:@65765.4]
  input         reset, // @[:@65766.4]
  output        io_in_cmd_ready, // @[:@65767.4]
  input         io_in_cmd_valid, // @[:@65767.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@65767.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@65767.4]
  input         io_in_cmd_bits_isWr, // @[:@65767.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@65767.4]
  output        io_in_wdata_ready, // @[:@65767.4]
  input         io_in_wdata_valid, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@65767.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@65767.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@65767.4]
  input         io_in_rresp_ready, // @[:@65767.4]
  input         io_in_wresp_ready, // @[:@65767.4]
  output        io_in_wresp_valid, // @[:@65767.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@65767.4]
  input         io_out_cmd_ready, // @[:@65767.4]
  output        io_out_cmd_valid, // @[:@65767.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@65767.4]
  output [31:0] io_out_cmd_bits_size, // @[:@65767.4]
  output        io_out_cmd_bits_isWr, // @[:@65767.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@65767.4]
  input         io_out_wdata_ready, // @[:@65767.4]
  output        io_out_wdata_valid, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@65767.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@65767.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@65767.4]
  output        io_out_wdata_bits_wlast, // @[:@65767.4]
  output        io_out_rresp_ready, // @[:@65767.4]
  output        io_out_wresp_ready, // @[:@65767.4]
  input         io_out_wresp_valid, // @[:@65767.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@65767.4]
);
  wire  wdataCounter_clock; // @[AXIProtocol.scala 59:28:@65881.4]
  wire  wdataCounter_reset; // @[AXIProtocol.scala 59:28:@65881.4]
  wire  wdataCounter_io_reset; // @[AXIProtocol.scala 59:28:@65881.4]
  wire  wdataCounter_io_enable; // @[AXIProtocol.scala 59:28:@65881.4]
  wire [31:0] wdataCounter_io_stride; // @[AXIProtocol.scala 59:28:@65881.4]
  wire [31:0] wdataCounter_io_out; // @[AXIProtocol.scala 59:28:@65881.4]
  wire [31:0] wdataCounter_io_next; // @[AXIProtocol.scala 59:28:@65881.4]
  reg  writeIssued; // @[AXIProtocol.scala 61:28:@65884.4]
  reg [31:0] _RAND_0;
  wire  dramCmdIssue; // @[AXIProtocol.scala 63:39:@65885.4]
  wire  dramWriteIssue; // @[AXIProtocol.scala 64:43:@65886.4]
  wire  _T_201; // @[AXIProtocol.scala 68:54:@65887.4]
  wire  wlast; // @[AXIProtocol.scala 68:30:@65888.4]
  wire  _T_203; // @[AXIProtocol.scala 72:28:@65894.6]
  wire  _GEN_0; // @[AXIProtocol.scala 72:40:@65895.6]
  wire  _GEN_1; // @[AXIProtocol.scala 70:15:@65890.4]
  wire  _T_208; // @[AXIProtocol.scala 84:55:@65904.4]
  wire  _T_210; // @[AXIProtocol.scala 84:44:@65905.4]
  Counter_72 wdataCounter ( // @[AXIProtocol.scala 59:28:@65881.4]
    .clock(wdataCounter_clock),
    .reset(wdataCounter_reset),
    .io_reset(wdataCounter_io_reset),
    .io_enable(wdataCounter_io_enable),
    .io_stride(wdataCounter_io_stride),
    .io_out(wdataCounter_io_out),
    .io_next(wdataCounter_io_next)
  );
  assign dramCmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 63:39:@65885.4]
  assign dramWriteIssue = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 64:43:@65886.4]
  assign _T_201 = wdataCounter_io_next == io_in_cmd_bits_size; // @[AXIProtocol.scala 68:54:@65887.4]
  assign wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 68:30:@65888.4]
  assign _T_203 = dramCmdIssue & io_in_cmd_bits_isWr; // @[AXIProtocol.scala 72:28:@65894.6]
  assign _GEN_0 = _T_203 ? 1'h1 : writeIssued; // @[AXIProtocol.scala 72:40:@65895.6]
  assign _GEN_1 = wlast ? 1'h0 : _GEN_0; // @[AXIProtocol.scala 70:15:@65890.4]
  assign _T_208 = writeIssued == 1'h0; // @[AXIProtocol.scala 84:55:@65904.4]
  assign _T_210 = io_in_cmd_bits_isWr ? _T_208 : 1'h1; // @[AXIProtocol.scala 84:44:@65905.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? wlast : dramCmdIssue; // @[AXIProtocol.scala 56:10:@65880.4 AXIProtocol.scala 81:19:@65902.4]
  assign io_in_wdata_ready = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 56:10:@65873.4 AXIProtocol.scala 82:21:@65903.4]
  assign io_in_wresp_valid = io_out_wresp_valid; // @[AXIProtocol.scala 56:10:@65770.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 56:10:@65769.4]
  assign io_out_cmd_valid = io_in_cmd_valid & _T_210; // @[AXIProtocol.scala 56:10:@65879.4 AXIProtocol.scala 84:20:@65907.4]
  assign io_out_cmd_bits_addr = io_in_cmd_bits_addr; // @[AXIProtocol.scala 56:10:@65878.4]
  assign io_out_cmd_bits_size = io_in_cmd_bits_size; // @[AXIProtocol.scala 56:10:@65877.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 56:10:@65875.4]
  assign io_out_cmd_bits_tag = io_in_cmd_bits_tag; // @[AXIProtocol.scala 56:10:@65874.4]
  assign io_out_wdata_valid = io_in_wdata_valid & writeIssued; // @[AXIProtocol.scala 56:10:@65872.4 AXIProtocol.scala 86:22:@65909.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 56:10:@65856.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 56:10:@65857.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 56:10:@65858.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 56:10:@65859.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 56:10:@65860.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 56:10:@65861.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 56:10:@65862.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 56:10:@65863.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 56:10:@65864.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 56:10:@65865.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 56:10:@65866.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 56:10:@65867.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 56:10:@65868.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 56:10:@65869.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 56:10:@65870.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 56:10:@65871.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 56:10:@65792.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 56:10:@65793.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 56:10:@65794.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 56:10:@65795.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 56:10:@65796.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 56:10:@65797.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 56:10:@65798.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 56:10:@65799.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 56:10:@65800.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 56:10:@65801.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 56:10:@65802.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 56:10:@65803.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 56:10:@65804.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 56:10:@65805.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 56:10:@65806.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 56:10:@65807.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 56:10:@65808.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 56:10:@65809.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 56:10:@65810.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 56:10:@65811.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 56:10:@65812.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 56:10:@65813.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 56:10:@65814.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 56:10:@65815.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 56:10:@65816.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 56:10:@65817.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 56:10:@65818.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 56:10:@65819.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 56:10:@65820.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 56:10:@65821.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 56:10:@65822.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 56:10:@65823.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 56:10:@65824.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 56:10:@65825.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 56:10:@65826.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 56:10:@65827.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 56:10:@65828.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 56:10:@65829.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 56:10:@65830.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 56:10:@65831.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 56:10:@65832.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 56:10:@65833.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 56:10:@65834.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 56:10:@65835.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 56:10:@65836.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 56:10:@65837.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 56:10:@65838.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 56:10:@65839.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 56:10:@65840.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 56:10:@65841.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 56:10:@65842.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 56:10:@65843.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 56:10:@65844.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 56:10:@65845.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 56:10:@65846.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 56:10:@65847.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 56:10:@65848.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 56:10:@65849.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 56:10:@65850.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 56:10:@65851.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 56:10:@65852.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 56:10:@65853.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 56:10:@65854.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 56:10:@65855.4]
  assign io_out_wdata_bits_wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 56:10:@65791.4 AXIProtocol.scala 87:27:@65910.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 56:10:@65790.4]
  assign io_out_wresp_ready = io_in_wresp_ready; // @[AXIProtocol.scala 56:10:@65771.4]
  assign wdataCounter_clock = clock; // @[:@65882.4]
  assign wdataCounter_reset = reset; // @[:@65883.4]
  assign wdataCounter_io_reset = dramWriteIssue & _T_201; // @[AXIProtocol.scala 76:25:@65898.4]
  assign wdataCounter_io_enable = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 77:26:@65899.4]
  assign wdataCounter_io_stride = 32'h1; // @[AXIProtocol.scala 78:26:@65900.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeIssued = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      writeIssued <= 1'h0;
    end else begin
      if (wlast) begin
        writeIssued <= 1'h0;
      end else begin
        if (_T_203) begin
          writeIssued <= 1'h1;
        end
      end
    end
  end
endmodule
module DRAMArbiter( // @[:@65912.2]
  input         clock, // @[:@65913.4]
  input         reset, // @[:@65914.4]
  input         io_enable, // @[:@65915.4]
  output        io_app_stores_0_cmd_ready, // @[:@65915.4]
  input         io_app_stores_0_cmd_valid, // @[:@65915.4]
  input  [63:0] io_app_stores_0_cmd_bits_addr, // @[:@65915.4]
  input  [31:0] io_app_stores_0_cmd_bits_size, // @[:@65915.4]
  output        io_app_stores_0_data_ready, // @[:@65915.4]
  input         io_app_stores_0_data_valid, // @[:@65915.4]
  input  [31:0] io_app_stores_0_data_bits_wdata_0, // @[:@65915.4]
  input         io_app_stores_0_data_bits_wstrb, // @[:@65915.4]
  input         io_app_stores_0_wresp_ready, // @[:@65915.4]
  output        io_app_stores_0_wresp_valid, // @[:@65915.4]
  output        io_app_stores_0_wresp_bits, // @[:@65915.4]
  input         io_dram_cmd_ready, // @[:@65915.4]
  output        io_dram_cmd_valid, // @[:@65915.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@65915.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@65915.4]
  output        io_dram_cmd_bits_isWr, // @[:@65915.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@65915.4]
  input         io_dram_wdata_ready, // @[:@65915.4]
  output        io_dram_wdata_valid, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@65915.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@65915.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@65915.4]
  output        io_dram_wdata_bits_wlast, // @[:@65915.4]
  output        io_dram_rresp_ready, // @[:@65915.4]
  output        io_dram_wresp_ready, // @[:@65915.4]
  input         io_dram_wresp_valid, // @[:@65915.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@65915.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@66801.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@66815.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@67043.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@67158.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@67158.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@66801.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@66815.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@67043.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@67158.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_app_stores_0_cmd_ready = StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 68:18:@66814.4]
  assign io_app_stores_0_data_ready = StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 68:18:@66810.4]
  assign io_app_stores_0_wresp_valid = StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 68:18:@66805.4]
  assign io_app_stores_0_wresp_bits = StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 68:18:@66804.4]
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@67383.4 DRAMArbiter.scala 100:23:@67386.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@67382.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@67381.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@67379.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@67378.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@67376.4 DRAMArbiter.scala 101:25:@67388.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@67360.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@67361.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@67362.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@67363.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@67364.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@67365.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@67366.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@67367.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@67368.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@67369.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@67370.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@67371.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@67372.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@67373.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@67374.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@67375.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@67296.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@67297.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@67298.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@67299.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@67300.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@67301.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@67302.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@67303.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@67304.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@67305.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@67306.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@67307.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@67308.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@67309.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@67310.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@67311.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@67312.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@67313.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@67314.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@67315.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@67316.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@67317.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@67318.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@67319.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@67320.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@67321.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@67322.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@67323.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@67324.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@67325.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@67326.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@67327.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@67328.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@67329.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@67330.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@67331.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@67332.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@67333.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@67334.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@67335.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@67336.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@67337.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@67338.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@67339.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@67340.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@67341.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@67342.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@67343.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@67344.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@67345.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@67346.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@67347.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@67348.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@67349.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@67350.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@67351.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@67352.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@67353.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@67354.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@67355.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@67356.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@67357.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@67358.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@67359.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@67295.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@67294.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@67275.4]
  assign StreamControllerStore_clock = clock; // @[:@66802.4]
  assign StreamControllerStore_reset = reset; // @[:@66803.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@66930.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@66923.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@66820.4]
  assign StreamControllerStore_io_store_cmd_valid = io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 68:18:@66813.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = io_app_stores_0_cmd_bits_addr; // @[DRAMArbiter.scala 68:18:@66812.4]
  assign StreamControllerStore_io_store_cmd_bits_size = io_app_stores_0_cmd_bits_size; // @[DRAMArbiter.scala 68:18:@66811.4]
  assign StreamControllerStore_io_store_data_valid = io_app_stores_0_data_valid; // @[DRAMArbiter.scala 68:18:@66809.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = io_app_stores_0_data_bits_wdata_0; // @[DRAMArbiter.scala 68:18:@66808.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = io_app_stores_0_data_bits_wstrb; // @[DRAMArbiter.scala 68:18:@66807.4]
  assign StreamControllerStore_io_store_wresp_ready = io_app_stores_0_wresp_ready; // @[DRAMArbiter.scala 68:18:@66806.4]
  assign StreamArbiter_clock = clock; // @[:@66816.4]
  assign StreamArbiter_reset = reset; // @[:@66817.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@67041.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@67040.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@67039.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@67037.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@67036.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@67034.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@67018.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@67019.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@67020.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@67021.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@67022.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@67023.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@67024.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@67025.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@67026.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@67027.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@67028.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@67029.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@67030.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@67031.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@67032.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@67033.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@66954.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@66955.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@66956.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@66957.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@66958.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@66959.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@66960.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@66961.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@66962.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@66963.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@66964.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@66965.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@66966.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@66967.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@66968.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@66969.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@66970.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@66971.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@66972.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@66973.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@66974.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@66975.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@66976.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@66977.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@66978.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@66979.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@66980.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@66981.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@66982.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@66983.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@66984.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@66985.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@66986.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@66987.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@66988.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@66989.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@66990.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@66991.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@66992.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@66993.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@66994.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@66995.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@66996.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@66997.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@66998.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@66999.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@67000.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@67001.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@67002.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@67003.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@67004.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@67005.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@67006.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@67007.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@67008.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@67009.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@67010.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@67011.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@67012.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@67013.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@67014.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@67015.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@67016.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@67017.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@66952.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@66933.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@67157.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@67150.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@67047.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@67046.4]
  assign AXICmdSplit_clock = clock; // @[:@67044.4]
  assign AXICmdSplit_reset = reset; // @[:@67045.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@67156.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@67155.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@67154.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@67152.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@67151.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@67149.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@67133.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@67134.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@67135.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@67136.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@67137.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@67138.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@67139.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@67140.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@67141.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@67142.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@67143.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@67144.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@67145.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@67146.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@67147.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@67148.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@67069.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@67070.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@67071.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@67072.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@67073.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@67074.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@67075.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@67076.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@67077.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@67078.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@67079.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@67080.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@67081.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@67082.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@67083.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@67084.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@67085.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@67086.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@67087.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@67088.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@67089.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@67090.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@67091.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@67092.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@67093.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@67094.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@67095.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@67096.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@67097.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@67098.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@67099.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@67100.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@67101.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@67102.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@67103.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@67104.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@67105.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@67106.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@67107.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@67108.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@67109.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@67110.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@67111.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@67112.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@67113.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@67114.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@67115.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@67116.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@67117.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@67118.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@67119.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@67120.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@67121.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@67122.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@67123.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@67124.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@67125.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@67126.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@67127.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@67128.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@67129.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@67130.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@67131.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@67132.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@67067.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@67048.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@67272.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@67265.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@67162.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@67161.4]
  assign AXICmdIssue_clock = clock; // @[:@67159.4]
  assign AXICmdIssue_reset = reset; // @[:@67160.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@67271.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@67270.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@67269.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@67267.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@67266.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@67264.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@67248.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@67249.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@67250.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@67251.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@67252.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@67253.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@67254.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@67255.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@67256.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@67257.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@67258.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@67259.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@67260.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@67261.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@67262.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@67263.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@67184.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@67185.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@67186.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@67187.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@67188.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@67189.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@67190.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@67191.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@67192.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@67193.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@67194.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@67195.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@67196.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@67197.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@67198.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@67199.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@67200.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@67201.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@67202.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@67203.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@67204.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@67205.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@67206.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@67207.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@67208.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@67209.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@67210.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@67211.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@67212.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@67213.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@67214.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@67215.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@67216.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@67217.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@67218.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@67219.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@67220.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@67221.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@67222.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@67223.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@67224.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@67225.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@67226.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@67227.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@67228.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@67229.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@67230.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@67231.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@67232.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@67233.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@67234.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@67235.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@67236.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@67237.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@67238.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@67239.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@67240.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@67241.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@67242.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@67243.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@67244.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@67245.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@67246.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@67247.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@67182.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@67163.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@67384.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@67377.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@67274.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@67273.4]
endmodule
module DRAMArbiter_1( // @[:@81613.2]
  input         clock, // @[:@81614.4]
  input         reset, // @[:@81615.4]
  input         io_enable, // @[:@81616.4]
  input         io_dram_cmd_ready, // @[:@81616.4]
  output        io_dram_cmd_valid, // @[:@81616.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@81616.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@81616.4]
  output        io_dram_cmd_bits_isWr, // @[:@81616.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@81616.4]
  input         io_dram_wdata_ready, // @[:@81616.4]
  output        io_dram_wdata_valid, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@81616.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@81616.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@81616.4]
  output        io_dram_wdata_bits_wlast, // @[:@81616.4]
  output        io_dram_rresp_ready, // @[:@81616.4]
  output        io_dram_wresp_ready, // @[:@81616.4]
  input         io_dram_wresp_valid, // @[:@81616.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@81616.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@82502.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@82516.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@82744.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@82859.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@82859.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@82502.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@82516.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@82744.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@82859.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@83084.4 DRAMArbiter.scala 100:23:@83087.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@83083.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@83082.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@83080.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@83079.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@83077.4 DRAMArbiter.scala 101:25:@83089.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@83061.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@83062.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@83063.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@83064.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@83065.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@83066.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@83067.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@83068.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@83069.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@83070.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@83071.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@83072.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@83073.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@83074.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@83075.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@83076.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@82997.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@82998.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@82999.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@83000.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@83001.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@83002.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@83003.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@83004.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@83005.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@83006.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@83007.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@83008.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@83009.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@83010.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@83011.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@83012.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@83013.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@83014.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@83015.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@83016.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@83017.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@83018.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@83019.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@83020.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@83021.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@83022.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@83023.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@83024.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@83025.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@83026.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@83027.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@83028.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@83029.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@83030.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@83031.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@83032.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@83033.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@83034.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@83035.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@83036.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@83037.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@83038.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@83039.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@83040.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@83041.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@83042.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@83043.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@83044.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@83045.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@83046.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@83047.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@83048.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@83049.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@83050.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@83051.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@83052.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@83053.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@83054.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@83055.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@83056.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@83057.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@83058.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@83059.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@83060.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@82996.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@82995.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@82976.4]
  assign StreamControllerStore_clock = clock; // @[:@82503.4]
  assign StreamControllerStore_reset = reset; // @[:@82504.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@82631.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@82624.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@82521.4]
  assign StreamControllerStore_io_store_cmd_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@82514.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = 64'h0; // @[DRAMArbiter.scala 68:18:@82513.4]
  assign StreamControllerStore_io_store_cmd_bits_size = 32'h0; // @[DRAMArbiter.scala 68:18:@82512.4]
  assign StreamControllerStore_io_store_data_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@82510.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = 32'h0; // @[DRAMArbiter.scala 68:18:@82509.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = 1'h0; // @[DRAMArbiter.scala 68:18:@82508.4]
  assign StreamControllerStore_io_store_wresp_ready = 1'h0; // @[DRAMArbiter.scala 68:18:@82507.4]
  assign StreamArbiter_clock = clock; // @[:@82517.4]
  assign StreamArbiter_reset = reset; // @[:@82518.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@82742.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@82741.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@82740.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@82738.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@82737.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@82735.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@82719.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@82720.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@82721.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@82722.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@82723.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@82724.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@82725.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@82726.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@82727.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@82728.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@82729.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@82730.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@82731.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@82732.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@82733.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@82734.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@82655.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@82656.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@82657.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@82658.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@82659.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@82660.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@82661.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@82662.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@82663.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@82664.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@82665.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@82666.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@82667.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@82668.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@82669.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@82670.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@82671.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@82672.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@82673.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@82674.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@82675.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@82676.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@82677.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@82678.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@82679.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@82680.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@82681.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@82682.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@82683.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@82684.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@82685.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@82686.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@82687.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@82688.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@82689.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@82690.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@82691.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@82692.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@82693.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@82694.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@82695.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@82696.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@82697.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@82698.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@82699.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@82700.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@82701.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@82702.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@82703.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@82704.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@82705.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@82706.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@82707.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@82708.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@82709.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@82710.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@82711.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@82712.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@82713.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@82714.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@82715.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@82716.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@82717.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@82718.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@82653.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@82634.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@82858.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@82851.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@82748.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@82747.4]
  assign AXICmdSplit_clock = clock; // @[:@82745.4]
  assign AXICmdSplit_reset = reset; // @[:@82746.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@82857.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@82856.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@82855.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@82853.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@82852.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@82850.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@82834.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@82835.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@82836.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@82837.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@82838.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@82839.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@82840.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@82841.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@82842.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@82843.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@82844.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@82845.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@82846.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@82847.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@82848.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@82849.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@82770.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@82771.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@82772.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@82773.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@82774.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@82775.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@82776.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@82777.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@82778.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@82779.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@82780.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@82781.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@82782.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@82783.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@82784.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@82785.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@82786.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@82787.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@82788.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@82789.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@82790.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@82791.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@82792.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@82793.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@82794.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@82795.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@82796.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@82797.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@82798.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@82799.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@82800.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@82801.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@82802.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@82803.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@82804.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@82805.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@82806.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@82807.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@82808.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@82809.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@82810.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@82811.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@82812.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@82813.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@82814.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@82815.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@82816.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@82817.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@82818.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@82819.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@82820.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@82821.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@82822.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@82823.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@82824.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@82825.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@82826.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@82827.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@82828.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@82829.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@82830.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@82831.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@82832.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@82833.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@82768.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@82749.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@82973.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@82966.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@82863.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@82862.4]
  assign AXICmdIssue_clock = clock; // @[:@82860.4]
  assign AXICmdIssue_reset = reset; // @[:@82861.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@82972.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@82971.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@82970.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@82968.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@82967.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@82965.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@82949.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@82950.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@82951.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@82952.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@82953.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@82954.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@82955.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@82956.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@82957.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@82958.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@82959.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@82960.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@82961.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@82962.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@82963.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@82964.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@82885.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@82886.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@82887.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@82888.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@82889.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@82890.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@82891.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@82892.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@82893.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@82894.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@82895.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@82896.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@82897.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@82898.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@82899.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@82900.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@82901.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@82902.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@82903.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@82904.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@82905.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@82906.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@82907.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@82908.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@82909.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@82910.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@82911.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@82912.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@82913.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@82914.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@82915.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@82916.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@82917.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@82918.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@82919.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@82920.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@82921.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@82922.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@82923.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@82924.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@82925.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@82926.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@82927.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@82928.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@82929.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@82930.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@82931.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@82932.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@82933.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@82934.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@82935.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@82936.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@82937.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@82938.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@82939.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@82940.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@82941.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@82942.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@82943.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@82944.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@82945.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@82946.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@82947.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@82948.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@82883.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@82864.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@83085.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@83078.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@82975.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@82974.4]
endmodule
module DRAMHeap( // @[:@113721.2]
  input         io_accel_0_req_valid, // @[:@113724.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@113724.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@113724.4]
  output        io_accel_0_resp_valid, // @[:@113724.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@113724.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@113724.4]
  output        io_host_0_req_valid, // @[:@113724.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@113724.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@113724.4]
  input         io_host_0_resp_valid, // @[:@113724.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@113724.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@113724.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@113731.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@113733.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@113732.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@113728.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@113727.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@113726.4]
endmodule
module RetimeWrapper_509( // @[:@113747.2]
  input         clock, // @[:@113748.4]
  input         reset, // @[:@113749.4]
  input         io_flow, // @[:@113750.4]
  input  [63:0] io_in, // @[:@113750.4]
  output [63:0] io_out // @[:@113750.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@113752.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@113752.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@113752.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@113752.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@113752.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@113752.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@113752.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@113765.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@113764.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@113763.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@113762.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@113761.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@113759.4]
endmodule
module FringeFF( // @[:@113767.2]
  input         clock, // @[:@113768.4]
  input         reset, // @[:@113769.4]
  input  [63:0] io_in, // @[:@113770.4]
  input         io_reset, // @[:@113770.4]
  output [63:0] io_out, // @[:@113770.4]
  input         io_enable // @[:@113770.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@113773.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@113773.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@113773.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@113773.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@113773.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@113778.4 package.scala 96:25:@113779.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@113784.6]
  RetimeWrapper_509 RetimeWrapper ( // @[package.scala 93:22:@113773.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@113778.4 package.scala 96:25:@113779.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@113784.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@113790.4]
  assign RetimeWrapper_clock = clock; // @[:@113774.4]
  assign RetimeWrapper_reset = reset; // @[:@113775.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@113777.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@113776.4]
endmodule
module MuxN( // @[:@142406.2]
  input  [63:0] io_ins_0, // @[:@142409.4]
  input  [63:0] io_ins_1, // @[:@142409.4]
  input  [63:0] io_ins_2, // @[:@142409.4]
  input  [63:0] io_ins_3, // @[:@142409.4]
  input  [63:0] io_ins_4, // @[:@142409.4]
  input  [63:0] io_ins_5, // @[:@142409.4]
  input  [63:0] io_ins_6, // @[:@142409.4]
  input  [63:0] io_ins_7, // @[:@142409.4]
  input  [63:0] io_ins_8, // @[:@142409.4]
  input  [63:0] io_ins_9, // @[:@142409.4]
  input  [63:0] io_ins_10, // @[:@142409.4]
  input  [63:0] io_ins_11, // @[:@142409.4]
  input  [63:0] io_ins_12, // @[:@142409.4]
  input  [63:0] io_ins_13, // @[:@142409.4]
  input  [63:0] io_ins_14, // @[:@142409.4]
  input  [63:0] io_ins_15, // @[:@142409.4]
  input  [63:0] io_ins_16, // @[:@142409.4]
  input  [63:0] io_ins_17, // @[:@142409.4]
  input  [63:0] io_ins_18, // @[:@142409.4]
  input  [63:0] io_ins_19, // @[:@142409.4]
  input  [63:0] io_ins_20, // @[:@142409.4]
  input  [63:0] io_ins_21, // @[:@142409.4]
  input  [63:0] io_ins_22, // @[:@142409.4]
  input  [63:0] io_ins_23, // @[:@142409.4]
  input  [63:0] io_ins_24, // @[:@142409.4]
  input  [63:0] io_ins_25, // @[:@142409.4]
  input  [63:0] io_ins_26, // @[:@142409.4]
  input  [63:0] io_ins_27, // @[:@142409.4]
  input  [63:0] io_ins_28, // @[:@142409.4]
  input  [63:0] io_ins_29, // @[:@142409.4]
  input  [63:0] io_ins_30, // @[:@142409.4]
  input  [63:0] io_ins_31, // @[:@142409.4]
  input  [63:0] io_ins_32, // @[:@142409.4]
  input  [63:0] io_ins_33, // @[:@142409.4]
  input  [63:0] io_ins_34, // @[:@142409.4]
  input  [63:0] io_ins_35, // @[:@142409.4]
  input  [63:0] io_ins_36, // @[:@142409.4]
  input  [63:0] io_ins_37, // @[:@142409.4]
  input  [63:0] io_ins_38, // @[:@142409.4]
  input  [63:0] io_ins_39, // @[:@142409.4]
  input  [63:0] io_ins_40, // @[:@142409.4]
  input  [63:0] io_ins_41, // @[:@142409.4]
  input  [63:0] io_ins_42, // @[:@142409.4]
  input  [63:0] io_ins_43, // @[:@142409.4]
  input  [63:0] io_ins_44, // @[:@142409.4]
  input  [63:0] io_ins_45, // @[:@142409.4]
  input  [63:0] io_ins_46, // @[:@142409.4]
  input  [63:0] io_ins_47, // @[:@142409.4]
  input  [63:0] io_ins_48, // @[:@142409.4]
  input  [63:0] io_ins_49, // @[:@142409.4]
  input  [63:0] io_ins_50, // @[:@142409.4]
  input  [63:0] io_ins_51, // @[:@142409.4]
  input  [63:0] io_ins_52, // @[:@142409.4]
  input  [63:0] io_ins_53, // @[:@142409.4]
  input  [63:0] io_ins_54, // @[:@142409.4]
  input  [63:0] io_ins_55, // @[:@142409.4]
  input  [63:0] io_ins_56, // @[:@142409.4]
  input  [63:0] io_ins_57, // @[:@142409.4]
  input  [63:0] io_ins_58, // @[:@142409.4]
  input  [63:0] io_ins_59, // @[:@142409.4]
  input  [63:0] io_ins_60, // @[:@142409.4]
  input  [63:0] io_ins_61, // @[:@142409.4]
  input  [63:0] io_ins_62, // @[:@142409.4]
  input  [63:0] io_ins_63, // @[:@142409.4]
  input  [63:0] io_ins_64, // @[:@142409.4]
  input  [63:0] io_ins_65, // @[:@142409.4]
  input  [63:0] io_ins_66, // @[:@142409.4]
  input  [63:0] io_ins_67, // @[:@142409.4]
  input  [63:0] io_ins_68, // @[:@142409.4]
  input  [63:0] io_ins_69, // @[:@142409.4]
  input  [63:0] io_ins_70, // @[:@142409.4]
  input  [63:0] io_ins_71, // @[:@142409.4]
  input  [63:0] io_ins_72, // @[:@142409.4]
  input  [63:0] io_ins_73, // @[:@142409.4]
  input  [63:0] io_ins_74, // @[:@142409.4]
  input  [63:0] io_ins_75, // @[:@142409.4]
  input  [63:0] io_ins_76, // @[:@142409.4]
  input  [63:0] io_ins_77, // @[:@142409.4]
  input  [63:0] io_ins_78, // @[:@142409.4]
  input  [63:0] io_ins_79, // @[:@142409.4]
  input  [63:0] io_ins_80, // @[:@142409.4]
  input  [63:0] io_ins_81, // @[:@142409.4]
  input  [63:0] io_ins_82, // @[:@142409.4]
  input  [63:0] io_ins_83, // @[:@142409.4]
  input  [63:0] io_ins_84, // @[:@142409.4]
  input  [63:0] io_ins_85, // @[:@142409.4]
  input  [63:0] io_ins_86, // @[:@142409.4]
  input  [63:0] io_ins_87, // @[:@142409.4]
  input  [63:0] io_ins_88, // @[:@142409.4]
  input  [63:0] io_ins_89, // @[:@142409.4]
  input  [63:0] io_ins_90, // @[:@142409.4]
  input  [63:0] io_ins_91, // @[:@142409.4]
  input  [63:0] io_ins_92, // @[:@142409.4]
  input  [63:0] io_ins_93, // @[:@142409.4]
  input  [63:0] io_ins_94, // @[:@142409.4]
  input  [63:0] io_ins_95, // @[:@142409.4]
  input  [63:0] io_ins_96, // @[:@142409.4]
  input  [63:0] io_ins_97, // @[:@142409.4]
  input  [63:0] io_ins_98, // @[:@142409.4]
  input  [63:0] io_ins_99, // @[:@142409.4]
  input  [63:0] io_ins_100, // @[:@142409.4]
  input  [63:0] io_ins_101, // @[:@142409.4]
  input  [63:0] io_ins_102, // @[:@142409.4]
  input  [63:0] io_ins_103, // @[:@142409.4]
  input  [63:0] io_ins_104, // @[:@142409.4]
  input  [63:0] io_ins_105, // @[:@142409.4]
  input  [63:0] io_ins_106, // @[:@142409.4]
  input  [63:0] io_ins_107, // @[:@142409.4]
  input  [63:0] io_ins_108, // @[:@142409.4]
  input  [63:0] io_ins_109, // @[:@142409.4]
  input  [63:0] io_ins_110, // @[:@142409.4]
  input  [63:0] io_ins_111, // @[:@142409.4]
  input  [63:0] io_ins_112, // @[:@142409.4]
  input  [63:0] io_ins_113, // @[:@142409.4]
  input  [63:0] io_ins_114, // @[:@142409.4]
  input  [63:0] io_ins_115, // @[:@142409.4]
  input  [63:0] io_ins_116, // @[:@142409.4]
  input  [63:0] io_ins_117, // @[:@142409.4]
  input  [63:0] io_ins_118, // @[:@142409.4]
  input  [63:0] io_ins_119, // @[:@142409.4]
  input  [63:0] io_ins_120, // @[:@142409.4]
  input  [63:0] io_ins_121, // @[:@142409.4]
  input  [63:0] io_ins_122, // @[:@142409.4]
  input  [63:0] io_ins_123, // @[:@142409.4]
  input  [63:0] io_ins_124, // @[:@142409.4]
  input  [63:0] io_ins_125, // @[:@142409.4]
  input  [63:0] io_ins_126, // @[:@142409.4]
  input  [63:0] io_ins_127, // @[:@142409.4]
  input  [63:0] io_ins_128, // @[:@142409.4]
  input  [63:0] io_ins_129, // @[:@142409.4]
  input  [63:0] io_ins_130, // @[:@142409.4]
  input  [63:0] io_ins_131, // @[:@142409.4]
  input  [63:0] io_ins_132, // @[:@142409.4]
  input  [63:0] io_ins_133, // @[:@142409.4]
  input  [63:0] io_ins_134, // @[:@142409.4]
  input  [63:0] io_ins_135, // @[:@142409.4]
  input  [63:0] io_ins_136, // @[:@142409.4]
  input  [63:0] io_ins_137, // @[:@142409.4]
  input  [63:0] io_ins_138, // @[:@142409.4]
  input  [63:0] io_ins_139, // @[:@142409.4]
  input  [63:0] io_ins_140, // @[:@142409.4]
  input  [63:0] io_ins_141, // @[:@142409.4]
  input  [63:0] io_ins_142, // @[:@142409.4]
  input  [63:0] io_ins_143, // @[:@142409.4]
  input  [63:0] io_ins_144, // @[:@142409.4]
  input  [63:0] io_ins_145, // @[:@142409.4]
  input  [63:0] io_ins_146, // @[:@142409.4]
  input  [63:0] io_ins_147, // @[:@142409.4]
  input  [63:0] io_ins_148, // @[:@142409.4]
  input  [63:0] io_ins_149, // @[:@142409.4]
  input  [63:0] io_ins_150, // @[:@142409.4]
  input  [63:0] io_ins_151, // @[:@142409.4]
  input  [63:0] io_ins_152, // @[:@142409.4]
  input  [63:0] io_ins_153, // @[:@142409.4]
  input  [63:0] io_ins_154, // @[:@142409.4]
  input  [63:0] io_ins_155, // @[:@142409.4]
  input  [63:0] io_ins_156, // @[:@142409.4]
  input  [63:0] io_ins_157, // @[:@142409.4]
  input  [63:0] io_ins_158, // @[:@142409.4]
  input  [63:0] io_ins_159, // @[:@142409.4]
  input  [63:0] io_ins_160, // @[:@142409.4]
  input  [63:0] io_ins_161, // @[:@142409.4]
  input  [63:0] io_ins_162, // @[:@142409.4]
  input  [63:0] io_ins_163, // @[:@142409.4]
  input  [63:0] io_ins_164, // @[:@142409.4]
  input  [63:0] io_ins_165, // @[:@142409.4]
  input  [63:0] io_ins_166, // @[:@142409.4]
  input  [63:0] io_ins_167, // @[:@142409.4]
  input  [63:0] io_ins_168, // @[:@142409.4]
  input  [63:0] io_ins_169, // @[:@142409.4]
  input  [63:0] io_ins_170, // @[:@142409.4]
  input  [63:0] io_ins_171, // @[:@142409.4]
  input  [63:0] io_ins_172, // @[:@142409.4]
  input  [63:0] io_ins_173, // @[:@142409.4]
  input  [63:0] io_ins_174, // @[:@142409.4]
  input  [63:0] io_ins_175, // @[:@142409.4]
  input  [63:0] io_ins_176, // @[:@142409.4]
  input  [63:0] io_ins_177, // @[:@142409.4]
  input  [63:0] io_ins_178, // @[:@142409.4]
  input  [63:0] io_ins_179, // @[:@142409.4]
  input  [63:0] io_ins_180, // @[:@142409.4]
  input  [63:0] io_ins_181, // @[:@142409.4]
  input  [63:0] io_ins_182, // @[:@142409.4]
  input  [63:0] io_ins_183, // @[:@142409.4]
  input  [63:0] io_ins_184, // @[:@142409.4]
  input  [63:0] io_ins_185, // @[:@142409.4]
  input  [63:0] io_ins_186, // @[:@142409.4]
  input  [63:0] io_ins_187, // @[:@142409.4]
  input  [63:0] io_ins_188, // @[:@142409.4]
  input  [63:0] io_ins_189, // @[:@142409.4]
  input  [63:0] io_ins_190, // @[:@142409.4]
  input  [63:0] io_ins_191, // @[:@142409.4]
  input  [63:0] io_ins_192, // @[:@142409.4]
  input  [63:0] io_ins_193, // @[:@142409.4]
  input  [63:0] io_ins_194, // @[:@142409.4]
  input  [63:0] io_ins_195, // @[:@142409.4]
  input  [63:0] io_ins_196, // @[:@142409.4]
  input  [63:0] io_ins_197, // @[:@142409.4]
  input  [63:0] io_ins_198, // @[:@142409.4]
  input  [63:0] io_ins_199, // @[:@142409.4]
  input  [63:0] io_ins_200, // @[:@142409.4]
  input  [63:0] io_ins_201, // @[:@142409.4]
  input  [63:0] io_ins_202, // @[:@142409.4]
  input  [63:0] io_ins_203, // @[:@142409.4]
  input  [63:0] io_ins_204, // @[:@142409.4]
  input  [63:0] io_ins_205, // @[:@142409.4]
  input  [63:0] io_ins_206, // @[:@142409.4]
  input  [63:0] io_ins_207, // @[:@142409.4]
  input  [63:0] io_ins_208, // @[:@142409.4]
  input  [63:0] io_ins_209, // @[:@142409.4]
  input  [63:0] io_ins_210, // @[:@142409.4]
  input  [63:0] io_ins_211, // @[:@142409.4]
  input  [63:0] io_ins_212, // @[:@142409.4]
  input  [63:0] io_ins_213, // @[:@142409.4]
  input  [63:0] io_ins_214, // @[:@142409.4]
  input  [63:0] io_ins_215, // @[:@142409.4]
  input  [63:0] io_ins_216, // @[:@142409.4]
  input  [63:0] io_ins_217, // @[:@142409.4]
  input  [63:0] io_ins_218, // @[:@142409.4]
  input  [63:0] io_ins_219, // @[:@142409.4]
  input  [63:0] io_ins_220, // @[:@142409.4]
  input  [63:0] io_ins_221, // @[:@142409.4]
  input  [63:0] io_ins_222, // @[:@142409.4]
  input  [63:0] io_ins_223, // @[:@142409.4]
  input  [63:0] io_ins_224, // @[:@142409.4]
  input  [63:0] io_ins_225, // @[:@142409.4]
  input  [63:0] io_ins_226, // @[:@142409.4]
  input  [63:0] io_ins_227, // @[:@142409.4]
  input  [63:0] io_ins_228, // @[:@142409.4]
  input  [63:0] io_ins_229, // @[:@142409.4]
  input  [63:0] io_ins_230, // @[:@142409.4]
  input  [63:0] io_ins_231, // @[:@142409.4]
  input  [63:0] io_ins_232, // @[:@142409.4]
  input  [63:0] io_ins_233, // @[:@142409.4]
  input  [63:0] io_ins_234, // @[:@142409.4]
  input  [63:0] io_ins_235, // @[:@142409.4]
  input  [63:0] io_ins_236, // @[:@142409.4]
  input  [63:0] io_ins_237, // @[:@142409.4]
  input  [63:0] io_ins_238, // @[:@142409.4]
  input  [63:0] io_ins_239, // @[:@142409.4]
  input  [63:0] io_ins_240, // @[:@142409.4]
  input  [63:0] io_ins_241, // @[:@142409.4]
  input  [63:0] io_ins_242, // @[:@142409.4]
  input  [63:0] io_ins_243, // @[:@142409.4]
  input  [63:0] io_ins_244, // @[:@142409.4]
  input  [63:0] io_ins_245, // @[:@142409.4]
  input  [63:0] io_ins_246, // @[:@142409.4]
  input  [63:0] io_ins_247, // @[:@142409.4]
  input  [63:0] io_ins_248, // @[:@142409.4]
  input  [63:0] io_ins_249, // @[:@142409.4]
  input  [63:0] io_ins_250, // @[:@142409.4]
  input  [63:0] io_ins_251, // @[:@142409.4]
  input  [63:0] io_ins_252, // @[:@142409.4]
  input  [63:0] io_ins_253, // @[:@142409.4]
  input  [63:0] io_ins_254, // @[:@142409.4]
  input  [63:0] io_ins_255, // @[:@142409.4]
  input  [63:0] io_ins_256, // @[:@142409.4]
  input  [63:0] io_ins_257, // @[:@142409.4]
  input  [63:0] io_ins_258, // @[:@142409.4]
  input  [63:0] io_ins_259, // @[:@142409.4]
  input  [63:0] io_ins_260, // @[:@142409.4]
  input  [63:0] io_ins_261, // @[:@142409.4]
  input  [63:0] io_ins_262, // @[:@142409.4]
  input  [63:0] io_ins_263, // @[:@142409.4]
  input  [63:0] io_ins_264, // @[:@142409.4]
  input  [63:0] io_ins_265, // @[:@142409.4]
  input  [63:0] io_ins_266, // @[:@142409.4]
  input  [63:0] io_ins_267, // @[:@142409.4]
  input  [63:0] io_ins_268, // @[:@142409.4]
  input  [63:0] io_ins_269, // @[:@142409.4]
  input  [63:0] io_ins_270, // @[:@142409.4]
  input  [63:0] io_ins_271, // @[:@142409.4]
  input  [63:0] io_ins_272, // @[:@142409.4]
  input  [63:0] io_ins_273, // @[:@142409.4]
  input  [63:0] io_ins_274, // @[:@142409.4]
  input  [63:0] io_ins_275, // @[:@142409.4]
  input  [63:0] io_ins_276, // @[:@142409.4]
  input  [63:0] io_ins_277, // @[:@142409.4]
  input  [63:0] io_ins_278, // @[:@142409.4]
  input  [63:0] io_ins_279, // @[:@142409.4]
  input  [63:0] io_ins_280, // @[:@142409.4]
  input  [63:0] io_ins_281, // @[:@142409.4]
  input  [63:0] io_ins_282, // @[:@142409.4]
  input  [63:0] io_ins_283, // @[:@142409.4]
  input  [63:0] io_ins_284, // @[:@142409.4]
  input  [63:0] io_ins_285, // @[:@142409.4]
  input  [63:0] io_ins_286, // @[:@142409.4]
  input  [63:0] io_ins_287, // @[:@142409.4]
  input  [63:0] io_ins_288, // @[:@142409.4]
  input  [63:0] io_ins_289, // @[:@142409.4]
  input  [63:0] io_ins_290, // @[:@142409.4]
  input  [63:0] io_ins_291, // @[:@142409.4]
  input  [63:0] io_ins_292, // @[:@142409.4]
  input  [63:0] io_ins_293, // @[:@142409.4]
  input  [63:0] io_ins_294, // @[:@142409.4]
  input  [63:0] io_ins_295, // @[:@142409.4]
  input  [63:0] io_ins_296, // @[:@142409.4]
  input  [63:0] io_ins_297, // @[:@142409.4]
  input  [63:0] io_ins_298, // @[:@142409.4]
  input  [63:0] io_ins_299, // @[:@142409.4]
  input  [63:0] io_ins_300, // @[:@142409.4]
  input  [63:0] io_ins_301, // @[:@142409.4]
  input  [63:0] io_ins_302, // @[:@142409.4]
  input  [63:0] io_ins_303, // @[:@142409.4]
  input  [63:0] io_ins_304, // @[:@142409.4]
  input  [63:0] io_ins_305, // @[:@142409.4]
  input  [63:0] io_ins_306, // @[:@142409.4]
  input  [63:0] io_ins_307, // @[:@142409.4]
  input  [63:0] io_ins_308, // @[:@142409.4]
  input  [63:0] io_ins_309, // @[:@142409.4]
  input  [63:0] io_ins_310, // @[:@142409.4]
  input  [63:0] io_ins_311, // @[:@142409.4]
  input  [63:0] io_ins_312, // @[:@142409.4]
  input  [63:0] io_ins_313, // @[:@142409.4]
  input  [63:0] io_ins_314, // @[:@142409.4]
  input  [63:0] io_ins_315, // @[:@142409.4]
  input  [63:0] io_ins_316, // @[:@142409.4]
  input  [63:0] io_ins_317, // @[:@142409.4]
  input  [63:0] io_ins_318, // @[:@142409.4]
  input  [63:0] io_ins_319, // @[:@142409.4]
  input  [63:0] io_ins_320, // @[:@142409.4]
  input  [63:0] io_ins_321, // @[:@142409.4]
  input  [63:0] io_ins_322, // @[:@142409.4]
  input  [63:0] io_ins_323, // @[:@142409.4]
  input  [63:0] io_ins_324, // @[:@142409.4]
  input  [63:0] io_ins_325, // @[:@142409.4]
  input  [63:0] io_ins_326, // @[:@142409.4]
  input  [63:0] io_ins_327, // @[:@142409.4]
  input  [63:0] io_ins_328, // @[:@142409.4]
  input  [63:0] io_ins_329, // @[:@142409.4]
  input  [63:0] io_ins_330, // @[:@142409.4]
  input  [63:0] io_ins_331, // @[:@142409.4]
  input  [63:0] io_ins_332, // @[:@142409.4]
  input  [63:0] io_ins_333, // @[:@142409.4]
  input  [63:0] io_ins_334, // @[:@142409.4]
  input  [63:0] io_ins_335, // @[:@142409.4]
  input  [63:0] io_ins_336, // @[:@142409.4]
  input  [63:0] io_ins_337, // @[:@142409.4]
  input  [63:0] io_ins_338, // @[:@142409.4]
  input  [63:0] io_ins_339, // @[:@142409.4]
  input  [63:0] io_ins_340, // @[:@142409.4]
  input  [63:0] io_ins_341, // @[:@142409.4]
  input  [63:0] io_ins_342, // @[:@142409.4]
  input  [63:0] io_ins_343, // @[:@142409.4]
  input  [63:0] io_ins_344, // @[:@142409.4]
  input  [63:0] io_ins_345, // @[:@142409.4]
  input  [63:0] io_ins_346, // @[:@142409.4]
  input  [63:0] io_ins_347, // @[:@142409.4]
  input  [63:0] io_ins_348, // @[:@142409.4]
  input  [63:0] io_ins_349, // @[:@142409.4]
  input  [63:0] io_ins_350, // @[:@142409.4]
  input  [63:0] io_ins_351, // @[:@142409.4]
  input  [63:0] io_ins_352, // @[:@142409.4]
  input  [63:0] io_ins_353, // @[:@142409.4]
  input  [63:0] io_ins_354, // @[:@142409.4]
  input  [63:0] io_ins_355, // @[:@142409.4]
  input  [63:0] io_ins_356, // @[:@142409.4]
  input  [63:0] io_ins_357, // @[:@142409.4]
  input  [63:0] io_ins_358, // @[:@142409.4]
  input  [63:0] io_ins_359, // @[:@142409.4]
  input  [63:0] io_ins_360, // @[:@142409.4]
  input  [63:0] io_ins_361, // @[:@142409.4]
  input  [63:0] io_ins_362, // @[:@142409.4]
  input  [63:0] io_ins_363, // @[:@142409.4]
  input  [63:0] io_ins_364, // @[:@142409.4]
  input  [63:0] io_ins_365, // @[:@142409.4]
  input  [63:0] io_ins_366, // @[:@142409.4]
  input  [63:0] io_ins_367, // @[:@142409.4]
  input  [63:0] io_ins_368, // @[:@142409.4]
  input  [63:0] io_ins_369, // @[:@142409.4]
  input  [63:0] io_ins_370, // @[:@142409.4]
  input  [63:0] io_ins_371, // @[:@142409.4]
  input  [63:0] io_ins_372, // @[:@142409.4]
  input  [63:0] io_ins_373, // @[:@142409.4]
  input  [63:0] io_ins_374, // @[:@142409.4]
  input  [63:0] io_ins_375, // @[:@142409.4]
  input  [63:0] io_ins_376, // @[:@142409.4]
  input  [63:0] io_ins_377, // @[:@142409.4]
  input  [63:0] io_ins_378, // @[:@142409.4]
  input  [63:0] io_ins_379, // @[:@142409.4]
  input  [63:0] io_ins_380, // @[:@142409.4]
  input  [63:0] io_ins_381, // @[:@142409.4]
  input  [63:0] io_ins_382, // @[:@142409.4]
  input  [63:0] io_ins_383, // @[:@142409.4]
  input  [63:0] io_ins_384, // @[:@142409.4]
  input  [63:0] io_ins_385, // @[:@142409.4]
  input  [63:0] io_ins_386, // @[:@142409.4]
  input  [63:0] io_ins_387, // @[:@142409.4]
  input  [63:0] io_ins_388, // @[:@142409.4]
  input  [63:0] io_ins_389, // @[:@142409.4]
  input  [63:0] io_ins_390, // @[:@142409.4]
  input  [63:0] io_ins_391, // @[:@142409.4]
  input  [63:0] io_ins_392, // @[:@142409.4]
  input  [63:0] io_ins_393, // @[:@142409.4]
  input  [63:0] io_ins_394, // @[:@142409.4]
  input  [63:0] io_ins_395, // @[:@142409.4]
  input  [63:0] io_ins_396, // @[:@142409.4]
  input  [63:0] io_ins_397, // @[:@142409.4]
  input  [63:0] io_ins_398, // @[:@142409.4]
  input  [63:0] io_ins_399, // @[:@142409.4]
  input  [63:0] io_ins_400, // @[:@142409.4]
  input  [63:0] io_ins_401, // @[:@142409.4]
  input  [63:0] io_ins_402, // @[:@142409.4]
  input  [63:0] io_ins_403, // @[:@142409.4]
  input  [63:0] io_ins_404, // @[:@142409.4]
  input  [63:0] io_ins_405, // @[:@142409.4]
  input  [63:0] io_ins_406, // @[:@142409.4]
  input  [63:0] io_ins_407, // @[:@142409.4]
  input  [63:0] io_ins_408, // @[:@142409.4]
  input  [63:0] io_ins_409, // @[:@142409.4]
  input  [63:0] io_ins_410, // @[:@142409.4]
  input  [63:0] io_ins_411, // @[:@142409.4]
  input  [63:0] io_ins_412, // @[:@142409.4]
  input  [63:0] io_ins_413, // @[:@142409.4]
  input  [63:0] io_ins_414, // @[:@142409.4]
  input  [63:0] io_ins_415, // @[:@142409.4]
  input  [63:0] io_ins_416, // @[:@142409.4]
  input  [63:0] io_ins_417, // @[:@142409.4]
  input  [63:0] io_ins_418, // @[:@142409.4]
  input  [63:0] io_ins_419, // @[:@142409.4]
  input  [63:0] io_ins_420, // @[:@142409.4]
  input  [63:0] io_ins_421, // @[:@142409.4]
  input  [63:0] io_ins_422, // @[:@142409.4]
  input  [63:0] io_ins_423, // @[:@142409.4]
  input  [63:0] io_ins_424, // @[:@142409.4]
  input  [63:0] io_ins_425, // @[:@142409.4]
  input  [63:0] io_ins_426, // @[:@142409.4]
  input  [63:0] io_ins_427, // @[:@142409.4]
  input  [63:0] io_ins_428, // @[:@142409.4]
  input  [63:0] io_ins_429, // @[:@142409.4]
  input  [63:0] io_ins_430, // @[:@142409.4]
  input  [63:0] io_ins_431, // @[:@142409.4]
  input  [63:0] io_ins_432, // @[:@142409.4]
  input  [63:0] io_ins_433, // @[:@142409.4]
  input  [63:0] io_ins_434, // @[:@142409.4]
  input  [63:0] io_ins_435, // @[:@142409.4]
  input  [63:0] io_ins_436, // @[:@142409.4]
  input  [63:0] io_ins_437, // @[:@142409.4]
  input  [63:0] io_ins_438, // @[:@142409.4]
  input  [63:0] io_ins_439, // @[:@142409.4]
  input  [63:0] io_ins_440, // @[:@142409.4]
  input  [63:0] io_ins_441, // @[:@142409.4]
  input  [63:0] io_ins_442, // @[:@142409.4]
  input  [63:0] io_ins_443, // @[:@142409.4]
  input  [63:0] io_ins_444, // @[:@142409.4]
  input  [63:0] io_ins_445, // @[:@142409.4]
  input  [63:0] io_ins_446, // @[:@142409.4]
  input  [63:0] io_ins_447, // @[:@142409.4]
  input  [63:0] io_ins_448, // @[:@142409.4]
  input  [63:0] io_ins_449, // @[:@142409.4]
  input  [63:0] io_ins_450, // @[:@142409.4]
  input  [63:0] io_ins_451, // @[:@142409.4]
  input  [63:0] io_ins_452, // @[:@142409.4]
  input  [63:0] io_ins_453, // @[:@142409.4]
  input  [63:0] io_ins_454, // @[:@142409.4]
  input  [63:0] io_ins_455, // @[:@142409.4]
  input  [63:0] io_ins_456, // @[:@142409.4]
  input  [63:0] io_ins_457, // @[:@142409.4]
  input  [63:0] io_ins_458, // @[:@142409.4]
  input  [63:0] io_ins_459, // @[:@142409.4]
  input  [63:0] io_ins_460, // @[:@142409.4]
  input  [63:0] io_ins_461, // @[:@142409.4]
  input  [63:0] io_ins_462, // @[:@142409.4]
  input  [63:0] io_ins_463, // @[:@142409.4]
  input  [63:0] io_ins_464, // @[:@142409.4]
  input  [63:0] io_ins_465, // @[:@142409.4]
  input  [63:0] io_ins_466, // @[:@142409.4]
  input  [63:0] io_ins_467, // @[:@142409.4]
  input  [63:0] io_ins_468, // @[:@142409.4]
  input  [63:0] io_ins_469, // @[:@142409.4]
  input  [63:0] io_ins_470, // @[:@142409.4]
  input  [63:0] io_ins_471, // @[:@142409.4]
  input  [63:0] io_ins_472, // @[:@142409.4]
  input  [63:0] io_ins_473, // @[:@142409.4]
  input  [63:0] io_ins_474, // @[:@142409.4]
  input  [63:0] io_ins_475, // @[:@142409.4]
  input  [63:0] io_ins_476, // @[:@142409.4]
  input  [63:0] io_ins_477, // @[:@142409.4]
  input  [63:0] io_ins_478, // @[:@142409.4]
  input  [63:0] io_ins_479, // @[:@142409.4]
  input  [63:0] io_ins_480, // @[:@142409.4]
  input  [63:0] io_ins_481, // @[:@142409.4]
  input  [63:0] io_ins_482, // @[:@142409.4]
  input  [63:0] io_ins_483, // @[:@142409.4]
  input  [63:0] io_ins_484, // @[:@142409.4]
  input  [63:0] io_ins_485, // @[:@142409.4]
  input  [63:0] io_ins_486, // @[:@142409.4]
  input  [63:0] io_ins_487, // @[:@142409.4]
  input  [63:0] io_ins_488, // @[:@142409.4]
  input  [63:0] io_ins_489, // @[:@142409.4]
  input  [63:0] io_ins_490, // @[:@142409.4]
  input  [63:0] io_ins_491, // @[:@142409.4]
  input  [63:0] io_ins_492, // @[:@142409.4]
  input  [63:0] io_ins_493, // @[:@142409.4]
  input  [63:0] io_ins_494, // @[:@142409.4]
  input  [63:0] io_ins_495, // @[:@142409.4]
  input  [63:0] io_ins_496, // @[:@142409.4]
  input  [63:0] io_ins_497, // @[:@142409.4]
  input  [63:0] io_ins_498, // @[:@142409.4]
  input  [63:0] io_ins_499, // @[:@142409.4]
  input  [63:0] io_ins_500, // @[:@142409.4]
  input  [63:0] io_ins_501, // @[:@142409.4]
  input  [63:0] io_ins_502, // @[:@142409.4]
  input  [8:0]  io_sel, // @[:@142409.4]
  output [63:0] io_out // @[:@142409.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@142411.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@142411.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@142411.4]
  assign io_out = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@142411.4]
endmodule
module RegFile( // @[:@142413.2]
  input         clock, // @[:@142414.4]
  input         reset, // @[:@142415.4]
  input  [31:0] io_raddr, // @[:@142416.4]
  input         io_wen, // @[:@142416.4]
  input  [31:0] io_waddr, // @[:@142416.4]
  input  [63:0] io_wdata, // @[:@142416.4]
  output [63:0] io_rdata, // @[:@142416.4]
  input         io_reset, // @[:@142416.4]
  output [63:0] io_argIns_0, // @[:@142416.4]
  output [63:0] io_argIns_1, // @[:@142416.4]
  output [63:0] io_argIns_2, // @[:@142416.4]
  output [63:0] io_argIns_3, // @[:@142416.4]
  input         io_argOuts_0_valid, // @[:@142416.4]
  input  [63:0] io_argOuts_0_bits, // @[:@142416.4]
  input         io_argOuts_1_valid, // @[:@142416.4]
  input  [63:0] io_argOuts_1_bits // @[:@142416.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@144426.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@144426.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@144426.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@144426.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@144426.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@144426.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@144438.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@144438.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@144438.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@144438.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@144438.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@144438.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@144457.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@144457.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@144457.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@144457.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@144457.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@144457.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@144469.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@144469.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@144469.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@144469.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@144469.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@144469.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@144481.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@144481.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@144481.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@144481.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@144481.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@144481.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@144495.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@144495.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@144495.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@144495.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@144495.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@144495.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@144509.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@144509.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@144509.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@144509.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@144509.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@144509.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@144523.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@144523.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@144523.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@144523.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@144523.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@144523.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@144537.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@144537.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@144537.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@144537.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@144537.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@144537.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@144551.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@144551.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@144551.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@144551.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@144551.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@144551.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@144565.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@144565.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@144565.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@144565.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@144565.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@144565.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@144579.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@144579.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@144579.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@144579.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@144579.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@144579.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@144593.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@144593.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@144593.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@144593.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@144593.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@144593.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@144607.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@144607.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@144607.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@144607.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@144607.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@144607.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@144621.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@144621.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@144621.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@144621.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@144621.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@144621.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@144635.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@144635.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@144635.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@144635.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@144635.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@144635.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@144649.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@144649.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@144649.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@144649.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@144649.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@144649.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@144663.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@144663.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@144663.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@144663.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@144663.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@144663.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@144677.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@144677.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@144677.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@144677.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@144677.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@144677.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@144691.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@144691.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@144691.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@144691.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@144691.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@144691.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@144705.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@144705.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@144705.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@144705.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@144705.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@144705.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@144719.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@144719.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@144719.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@144719.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@144719.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@144719.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@144733.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@144733.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@144733.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@144733.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@144733.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@144733.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@144747.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@144747.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@144747.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@144747.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@144747.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@144747.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@144761.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@144761.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@144761.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@144761.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@144761.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@144761.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@144775.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@144775.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@144775.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@144775.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@144775.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@144775.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@144789.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@144789.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@144789.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@144789.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@144789.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@144789.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@144803.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@144803.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@144803.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@144803.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@144803.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@144803.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@144817.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@144817.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@144817.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@144817.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@144817.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@144817.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@144831.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@144831.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@144831.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@144831.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@144831.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@144831.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@144845.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@144845.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@144845.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@144845.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@144845.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@144845.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@144859.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@144859.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@144859.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@144859.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@144859.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@144859.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@144873.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@144873.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@144873.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@144873.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@144873.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@144873.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@144887.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@144887.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@144887.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@144887.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@144887.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@144887.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@144901.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@144901.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@144901.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@144901.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@144901.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@144901.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@144915.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@144915.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@144915.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@144915.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@144915.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@144915.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@144929.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@144929.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@144929.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@144929.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@144929.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@144929.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@144943.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@144943.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@144943.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@144943.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@144943.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@144943.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@144957.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@144957.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@144957.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@144957.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@144957.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@144957.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@144971.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@144971.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@144971.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@144971.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@144971.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@144971.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@144985.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@144985.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@144985.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@144985.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@144985.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@144985.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@144999.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@144999.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@144999.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@144999.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@144999.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@144999.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@145013.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@145013.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@145013.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@145013.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@145013.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@145013.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@145027.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@145027.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@145027.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@145027.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@145027.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@145027.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@145041.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@145041.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@145041.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@145041.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@145041.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@145041.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@145055.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@145055.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@145055.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@145055.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@145055.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@145055.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@145069.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@145069.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@145069.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@145069.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@145069.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@145069.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@145083.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@145083.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@145083.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@145083.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@145083.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@145083.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@145097.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@145097.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@145097.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@145097.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@145097.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@145097.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@145111.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@145111.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@145111.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@145111.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@145111.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@145111.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@145125.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@145125.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@145125.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@145125.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@145125.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@145125.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@145139.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@145139.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@145139.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@145139.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@145139.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@145139.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@145153.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@145153.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@145153.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@145153.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@145153.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@145153.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@145167.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@145167.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@145167.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@145167.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@145167.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@145167.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@145181.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@145181.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@145181.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@145181.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@145181.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@145181.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@145195.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@145195.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@145195.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@145195.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@145195.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@145195.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@145209.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@145209.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@145209.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@145209.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@145209.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@145209.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@145223.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@145223.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@145223.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@145223.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@145223.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@145223.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@145237.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@145237.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@145237.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@145237.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@145237.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@145237.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@145251.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@145251.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@145251.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@145251.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@145251.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@145251.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@145265.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@145265.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@145265.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@145265.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@145265.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@145265.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@145279.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@145279.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@145279.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@145279.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@145279.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@145279.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@145293.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@145293.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@145293.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@145293.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@145293.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@145293.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@145307.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@145307.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@145307.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@145307.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@145307.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@145307.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@145321.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@145321.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@145321.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@145321.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@145321.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@145321.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@145335.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@145335.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@145335.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@145335.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@145335.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@145335.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@145349.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@145349.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@145349.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@145349.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@145349.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@145349.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@145363.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@145363.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@145363.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@145363.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@145363.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@145363.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@145377.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@145377.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@145377.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@145377.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@145377.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@145377.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@145391.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@145391.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@145391.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@145391.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@145391.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@145391.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@145405.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@145405.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@145405.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@145405.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@145405.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@145405.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@145419.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@145419.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@145419.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@145419.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@145419.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@145419.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@145433.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@145433.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@145433.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@145433.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@145433.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@145433.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@145447.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@145447.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@145447.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@145447.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@145447.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@145447.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@145461.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@145461.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@145461.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@145461.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@145461.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@145461.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@145475.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@145475.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@145475.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@145475.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@145475.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@145475.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@145489.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@145489.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@145489.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@145489.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@145489.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@145489.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@145503.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@145503.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@145503.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@145503.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@145503.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@145503.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@145517.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@145517.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@145517.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@145517.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@145517.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@145517.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@145531.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@145531.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@145531.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@145531.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@145531.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@145531.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@145545.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@145545.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@145545.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@145545.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@145545.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@145545.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@145559.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@145559.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@145559.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@145559.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@145559.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@145559.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@145573.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@145573.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@145573.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@145573.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@145573.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@145573.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@145587.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@145587.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@145587.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@145587.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@145587.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@145587.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@145601.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@145601.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@145601.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@145601.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@145601.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@145601.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@145615.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@145615.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@145615.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@145615.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@145615.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@145615.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@145629.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@145629.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@145629.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@145629.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@145629.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@145629.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@145643.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@145643.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@145643.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@145643.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@145643.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@145643.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@145657.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@145657.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@145657.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@145657.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@145657.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@145657.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@145671.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@145671.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@145671.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@145671.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@145671.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@145671.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@145685.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@145685.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@145685.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@145685.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@145685.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@145685.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@145699.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@145699.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@145699.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@145699.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@145699.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@145699.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@145713.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@145713.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@145713.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@145713.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@145713.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@145713.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@145727.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@145727.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@145727.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@145727.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@145727.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@145727.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@145741.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@145741.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@145741.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@145741.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@145741.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@145741.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@145755.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@145755.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@145755.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@145755.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@145755.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@145755.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@145769.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@145769.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@145769.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@145769.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@145769.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@145769.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@145783.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@145783.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@145783.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@145783.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@145783.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@145783.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@145797.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@145797.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@145797.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@145797.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@145797.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@145797.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@145811.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@145811.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@145811.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@145811.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@145811.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@145811.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@145825.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@145825.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@145825.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@145825.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@145825.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@145825.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@145839.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@145839.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@145839.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@145839.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@145839.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@145839.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@145853.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@145853.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@145853.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@145853.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@145853.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@145853.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@145867.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@145867.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@145867.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@145867.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@145867.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@145867.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@145881.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@145881.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@145881.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@145881.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@145881.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@145881.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@145895.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@145895.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@145895.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@145895.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@145895.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@145895.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@145909.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@145909.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@145909.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@145909.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@145909.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@145909.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@145923.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@145923.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@145923.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@145923.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@145923.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@145923.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@145937.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@145937.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@145937.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@145937.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@145937.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@145937.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@145951.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@145951.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@145951.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@145951.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@145951.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@145951.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@145965.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@145965.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@145965.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@145965.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@145965.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@145965.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@145979.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@145979.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@145979.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@145979.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@145979.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@145979.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@145993.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@145993.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@145993.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@145993.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@145993.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@145993.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@146007.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@146007.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@146007.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@146007.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@146007.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@146007.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@146021.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@146021.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@146021.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@146021.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@146021.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@146021.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@146035.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@146035.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@146035.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@146035.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@146035.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@146035.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@146049.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@146049.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@146049.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@146049.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@146049.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@146049.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@146063.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@146063.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@146063.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@146063.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@146063.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@146063.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@146077.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@146077.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@146077.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@146077.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@146077.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@146077.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@146091.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@146091.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@146091.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@146091.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@146091.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@146091.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@146105.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@146105.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@146105.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@146105.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@146105.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@146105.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@146119.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@146119.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@146119.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@146119.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@146119.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@146119.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@146133.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@146133.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@146133.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@146133.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@146133.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@146133.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@146147.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@146147.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@146147.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@146147.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@146147.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@146147.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@146161.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@146161.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@146161.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@146161.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@146161.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@146161.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@146175.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@146175.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@146175.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@146175.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@146175.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@146175.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@146189.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@146189.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@146189.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@146189.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@146189.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@146189.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@146203.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@146203.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@146203.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@146203.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@146203.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@146203.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@146217.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@146217.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@146217.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@146217.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@146217.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@146217.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@146231.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@146231.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@146231.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@146231.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@146231.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@146231.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@146245.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@146245.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@146245.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@146245.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@146245.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@146245.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@146259.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@146259.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@146259.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@146259.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@146259.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@146259.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@146273.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@146273.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@146273.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@146273.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@146273.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@146273.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@146287.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@146287.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@146287.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@146287.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@146287.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@146287.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@146301.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@146301.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@146301.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@146301.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@146301.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@146301.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@146315.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@146315.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@146315.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@146315.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@146315.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@146315.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@146329.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@146329.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@146329.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@146329.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@146329.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@146329.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@146343.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@146343.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@146343.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@146343.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@146343.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@146343.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@146357.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@146357.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@146357.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@146357.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@146357.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@146357.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@146371.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@146371.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@146371.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@146371.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@146371.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@146371.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@146385.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@146385.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@146385.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@146385.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@146385.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@146385.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@146399.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@146399.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@146399.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@146399.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@146399.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@146399.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@146413.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@146413.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@146413.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@146413.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@146413.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@146413.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@146427.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@146427.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@146427.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@146427.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@146427.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@146427.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@146441.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@146441.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@146441.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@146441.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@146441.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@146441.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@146455.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@146455.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@146455.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@146455.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@146455.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@146455.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@146469.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@146469.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@146469.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@146469.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@146469.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@146469.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@146483.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@146483.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@146483.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@146483.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@146483.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@146483.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@146497.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@146497.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@146497.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@146497.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@146497.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@146497.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@146511.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@146511.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@146511.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@146511.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@146511.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@146511.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@146525.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@146525.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@146525.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@146525.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@146525.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@146525.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@146539.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@146539.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@146539.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@146539.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@146539.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@146539.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@146553.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@146553.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@146553.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@146553.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@146553.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@146553.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@146567.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@146567.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@146567.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@146567.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@146567.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@146567.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@146581.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@146581.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@146581.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@146581.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@146581.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@146581.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@146595.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@146595.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@146595.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@146595.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@146595.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@146595.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@146609.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@146609.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@146609.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@146609.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@146609.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@146609.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@146623.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@146623.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@146623.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@146623.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@146623.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@146623.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@146637.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@146637.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@146637.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@146637.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@146637.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@146637.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@146651.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@146651.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@146651.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@146651.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@146651.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@146651.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@146665.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@146665.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@146665.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@146665.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@146665.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@146665.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@146679.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@146679.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@146679.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@146679.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@146679.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@146679.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@146693.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@146693.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@146693.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@146693.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@146693.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@146693.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@146707.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@146707.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@146707.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@146707.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@146707.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@146707.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@146721.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@146721.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@146721.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@146721.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@146721.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@146721.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@146735.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@146735.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@146735.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@146735.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@146735.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@146735.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@146749.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@146749.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@146749.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@146749.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@146749.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@146749.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@146763.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@146763.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@146763.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@146763.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@146763.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@146763.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@146777.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@146777.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@146777.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@146777.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@146777.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@146777.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@146791.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@146791.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@146791.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@146791.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@146791.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@146791.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@146805.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@146805.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@146805.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@146805.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@146805.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@146805.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@146819.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@146819.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@146819.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@146819.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@146819.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@146819.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@146833.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@146833.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@146833.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@146833.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@146833.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@146833.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@146847.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@146847.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@146847.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@146847.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@146847.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@146847.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@146861.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@146861.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@146861.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@146861.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@146861.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@146861.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@146875.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@146875.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@146875.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@146875.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@146875.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@146875.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@146889.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@146889.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@146889.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@146889.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@146889.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@146889.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@146903.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@146903.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@146903.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@146903.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@146903.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@146903.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@146917.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@146917.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@146917.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@146917.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@146917.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@146917.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@146931.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@146931.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@146931.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@146931.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@146931.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@146931.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@146945.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@146945.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@146945.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@146945.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@146945.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@146945.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@146959.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@146959.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@146959.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@146959.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@146959.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@146959.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@146973.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@146973.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@146973.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@146973.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@146973.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@146973.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@146987.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@146987.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@146987.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@146987.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@146987.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@146987.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@147001.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@147001.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@147001.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@147001.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@147001.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@147001.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@147015.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@147015.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@147015.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@147015.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@147015.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@147015.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@147029.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@147029.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@147029.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@147029.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@147029.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@147029.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@147043.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@147043.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@147043.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@147043.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@147043.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@147043.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@147057.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@147057.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@147057.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@147057.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@147057.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@147057.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@147071.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@147071.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@147071.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@147071.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@147071.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@147071.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@147085.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@147085.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@147085.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@147085.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@147085.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@147085.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@147099.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@147099.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@147099.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@147099.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@147099.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@147099.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@147113.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@147113.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@147113.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@147113.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@147113.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@147113.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@147127.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@147127.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@147127.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@147127.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@147127.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@147127.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@147141.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@147141.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@147141.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@147141.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@147141.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@147141.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@147155.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@147155.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@147155.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@147155.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@147155.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@147155.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@147169.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@147169.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@147169.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@147169.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@147169.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@147169.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@147183.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@147183.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@147183.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@147183.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@147183.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@147183.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@147197.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@147197.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@147197.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@147197.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@147197.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@147197.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@147211.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@147211.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@147211.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@147211.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@147211.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@147211.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@147225.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@147225.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@147225.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@147225.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@147225.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@147225.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@147239.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@147239.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@147239.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@147239.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@147239.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@147239.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@147253.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@147253.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@147253.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@147253.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@147253.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@147253.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@147267.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@147267.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@147267.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@147267.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@147267.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@147267.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@147281.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@147281.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@147281.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@147281.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@147281.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@147281.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@147295.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@147295.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@147295.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@147295.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@147295.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@147295.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@147309.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@147309.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@147309.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@147309.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@147309.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@147309.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@147323.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@147323.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@147323.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@147323.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@147323.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@147323.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@147337.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@147337.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@147337.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@147337.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@147337.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@147337.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@147351.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@147351.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@147351.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@147351.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@147351.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@147351.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@147365.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@147365.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@147365.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@147365.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@147365.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@147365.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@147379.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@147379.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@147379.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@147379.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@147379.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@147379.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@147393.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@147393.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@147393.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@147393.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@147393.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@147393.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@147407.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@147407.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@147407.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@147407.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@147407.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@147407.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@147421.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@147421.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@147421.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@147421.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@147421.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@147421.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@147435.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@147435.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@147435.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@147435.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@147435.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@147435.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@147449.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@147449.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@147449.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@147449.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@147449.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@147449.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@147463.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@147463.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@147463.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@147463.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@147463.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@147463.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@147477.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@147477.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@147477.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@147477.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@147477.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@147477.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@147491.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@147491.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@147491.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@147491.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@147491.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@147491.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@147505.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@147505.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@147505.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@147505.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@147505.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@147505.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@147519.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@147519.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@147519.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@147519.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@147519.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@147519.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@147533.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@147533.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@147533.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@147533.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@147533.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@147533.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@147547.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@147547.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@147547.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@147547.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@147547.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@147547.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@147561.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@147561.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@147561.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@147561.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@147561.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@147561.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@147575.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@147575.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@147575.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@147575.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@147575.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@147575.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@147589.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@147589.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@147589.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@147589.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@147589.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@147589.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@147603.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@147603.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@147603.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@147603.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@147603.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@147603.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@147617.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@147617.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@147617.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@147617.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@147617.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@147617.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@147631.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@147631.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@147631.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@147631.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@147631.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@147631.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@147645.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@147645.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@147645.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@147645.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@147645.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@147645.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@147659.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@147659.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@147659.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@147659.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@147659.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@147659.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@147673.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@147673.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@147673.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@147673.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@147673.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@147673.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@147687.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@147687.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@147687.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@147687.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@147687.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@147687.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@147701.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@147701.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@147701.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@147701.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@147701.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@147701.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@147715.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@147715.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@147715.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@147715.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@147715.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@147715.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@147729.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@147729.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@147729.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@147729.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@147729.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@147729.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@147743.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@147743.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@147743.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@147743.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@147743.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@147743.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@147757.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@147757.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@147757.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@147757.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@147757.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@147757.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@147771.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@147771.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@147771.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@147771.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@147771.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@147771.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@147785.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@147785.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@147785.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@147785.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@147785.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@147785.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@147799.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@147799.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@147799.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@147799.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@147799.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@147799.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@147813.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@147813.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@147813.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@147813.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@147813.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@147813.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@147827.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@147827.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@147827.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@147827.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@147827.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@147827.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@147841.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@147841.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@147841.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@147841.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@147841.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@147841.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@147855.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@147855.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@147855.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@147855.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@147855.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@147855.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@147869.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@147869.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@147869.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@147869.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@147869.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@147869.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@147883.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@147883.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@147883.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@147883.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@147883.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@147883.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@147897.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@147897.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@147897.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@147897.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@147897.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@147897.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@147911.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@147911.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@147911.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@147911.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@147911.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@147911.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@147925.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@147925.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@147925.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@147925.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@147925.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@147925.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@147939.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@147939.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@147939.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@147939.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@147939.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@147939.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@147953.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@147953.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@147953.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@147953.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@147953.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@147953.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@147967.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@147967.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@147967.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@147967.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@147967.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@147967.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@147981.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@147981.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@147981.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@147981.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@147981.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@147981.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@147995.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@147995.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@147995.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@147995.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@147995.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@147995.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@148009.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@148009.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@148009.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@148009.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@148009.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@148009.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@148023.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@148023.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@148023.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@148023.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@148023.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@148023.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@148037.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@148037.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@148037.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@148037.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@148037.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@148037.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@148051.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@148051.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@148051.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@148051.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@148051.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@148051.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@148065.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@148065.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@148065.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@148065.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@148065.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@148065.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@148079.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@148079.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@148079.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@148079.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@148079.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@148079.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@148093.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@148093.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@148093.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@148093.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@148093.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@148093.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@148107.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@148107.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@148107.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@148107.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@148107.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@148107.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@148121.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@148121.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@148121.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@148121.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@148121.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@148121.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@148135.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@148135.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@148135.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@148135.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@148135.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@148135.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@148149.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@148149.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@148149.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@148149.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@148149.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@148149.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@148163.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@148163.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@148163.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@148163.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@148163.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@148163.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@148177.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@148177.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@148177.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@148177.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@148177.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@148177.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@148191.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@148191.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@148191.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@148191.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@148191.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@148191.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@148205.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@148205.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@148205.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@148205.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@148205.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@148205.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@148219.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@148219.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@148219.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@148219.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@148219.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@148219.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@148233.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@148233.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@148233.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@148233.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@148233.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@148233.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@148247.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@148247.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@148247.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@148247.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@148247.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@148247.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@148261.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@148261.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@148261.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@148261.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@148261.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@148261.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@148275.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@148275.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@148275.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@148275.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@148275.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@148275.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@148289.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@148289.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@148289.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@148289.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@148289.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@148289.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@148303.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@148303.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@148303.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@148303.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@148303.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@148303.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@148317.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@148317.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@148317.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@148317.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@148317.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@148317.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@148331.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@148331.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@148331.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@148331.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@148331.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@148331.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@148345.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@148345.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@148345.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@148345.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@148345.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@148345.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@148359.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@148359.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@148359.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@148359.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@148359.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@148359.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@148373.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@148373.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@148373.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@148373.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@148373.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@148373.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@148387.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@148387.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@148387.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@148387.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@148387.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@148387.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@148401.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@148401.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@148401.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@148401.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@148401.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@148401.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@148415.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@148415.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@148415.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@148415.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@148415.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@148415.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@148429.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@148429.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@148429.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@148429.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@148429.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@148429.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@148443.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@148443.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@148443.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@148443.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@148443.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@148443.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@148457.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@148457.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@148457.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@148457.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@148457.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@148457.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@148471.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@148471.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@148471.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@148471.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@148471.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@148471.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@148485.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@148485.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@148485.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@148485.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@148485.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@148485.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@148499.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@148499.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@148499.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@148499.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@148499.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@148499.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@148513.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@148513.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@148513.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@148513.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@148513.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@148513.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@148527.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@148527.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@148527.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@148527.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@148527.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@148527.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@148541.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@148541.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@148541.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@148541.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@148541.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@148541.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@148555.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@148555.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@148555.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@148555.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@148555.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@148555.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@148569.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@148569.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@148569.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@148569.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@148569.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@148569.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@148583.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@148583.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@148583.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@148583.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@148583.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@148583.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@148597.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@148597.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@148597.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@148597.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@148597.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@148597.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@148611.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@148611.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@148611.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@148611.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@148611.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@148611.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@148625.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@148625.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@148625.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@148625.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@148625.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@148625.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@148639.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@148639.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@148639.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@148639.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@148639.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@148639.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@148653.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@148653.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@148653.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@148653.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@148653.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@148653.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@148667.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@148667.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@148667.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@148667.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@148667.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@148667.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@148681.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@148681.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@148681.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@148681.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@148681.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@148681.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@148695.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@148695.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@148695.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@148695.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@148695.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@148695.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@148709.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@148709.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@148709.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@148709.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@148709.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@148709.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@148723.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@148723.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@148723.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@148723.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@148723.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@148723.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@148737.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@148737.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@148737.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@148737.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@148737.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@148737.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@148751.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@148751.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@148751.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@148751.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@148751.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@148751.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@148765.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@148765.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@148765.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@148765.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@148765.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@148765.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@148779.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@148779.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@148779.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@148779.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@148779.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@148779.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@148793.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@148793.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@148793.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@148793.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@148793.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@148793.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@148807.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@148807.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@148807.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@148807.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@148807.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@148807.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@148821.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@148821.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@148821.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@148821.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@148821.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@148821.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@148835.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@148835.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@148835.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@148835.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@148835.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@148835.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@148849.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@148849.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@148849.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@148849.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@148849.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@148849.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@148863.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@148863.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@148863.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@148863.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@148863.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@148863.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@148877.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@148877.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@148877.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@148877.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@148877.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@148877.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@148891.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@148891.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@148891.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@148891.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@148891.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@148891.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@148905.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@148905.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@148905.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@148905.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@148905.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@148905.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@148919.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@148919.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@148919.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@148919.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@148919.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@148919.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@148933.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@148933.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@148933.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@148933.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@148933.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@148933.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@148947.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@148947.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@148947.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@148947.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@148947.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@148947.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@148961.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@148961.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@148961.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@148961.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@148961.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@148961.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@148975.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@148975.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@148975.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@148975.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@148975.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@148975.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@148989.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@148989.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@148989.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@148989.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@148989.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@148989.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@149003.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@149003.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@149003.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@149003.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@149003.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@149003.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@149017.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@149017.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@149017.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@149017.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@149017.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@149017.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@149031.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@149031.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@149031.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@149031.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@149031.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@149031.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@149045.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@149045.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@149045.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@149045.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@149045.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@149045.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@149059.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@149059.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@149059.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@149059.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@149059.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@149059.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@149073.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@149073.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@149073.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@149073.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@149073.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@149073.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@149087.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@149087.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@149087.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@149087.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@149087.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@149087.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@149101.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@149101.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@149101.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@149101.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@149101.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@149101.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@149115.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@149115.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@149115.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@149115.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@149115.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@149115.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@149129.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@149129.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@149129.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@149129.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@149129.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@149129.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@149143.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@149143.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@149143.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@149143.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@149143.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@149143.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@149157.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@149157.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@149157.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@149157.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@149157.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@149157.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@149171.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@149171.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@149171.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@149171.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@149171.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@149171.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@149185.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@149185.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@149185.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@149185.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@149185.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@149185.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@149199.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@149199.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@149199.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@149199.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@149199.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@149199.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@149213.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@149213.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@149213.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@149213.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@149213.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@149213.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@149227.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@149227.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@149227.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@149227.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@149227.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@149227.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@149241.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@149241.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@149241.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@149241.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@149241.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@149241.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@149255.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@149255.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@149255.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@149255.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@149255.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@149255.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@149269.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@149269.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@149269.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@149269.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@149269.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@149269.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@149283.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@149283.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@149283.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@149283.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@149283.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@149283.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@149297.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@149297.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@149297.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@149297.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@149297.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@149297.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@149311.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@149311.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@149311.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@149311.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@149311.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@149311.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@149325.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@149325.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@149325.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@149325.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@149325.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@149325.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@149339.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@149339.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@149339.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@149339.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@149339.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@149339.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@149353.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@149353.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@149353.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@149353.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@149353.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@149353.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@149367.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@149367.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@149367.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@149367.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@149367.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@149367.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@149381.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@149381.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@149381.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@149381.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@149381.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@149381.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@149395.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@149395.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@149395.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@149395.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@149395.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@149395.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@149409.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@149409.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@149409.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@149409.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@149409.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@149409.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@149423.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@149423.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@149423.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@149423.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@149423.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@149423.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@149437.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@149437.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@149437.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@149437.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@149437.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@149437.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@149451.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@149451.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@149451.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@149451.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@149451.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@149451.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@149465.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@149465.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@149465.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@149465.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@149465.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@149465.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@149479.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@149479.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@149479.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@149479.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@149479.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@149479.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@149493.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@149493.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@149493.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@149493.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@149493.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@149493.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@149507.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@149507.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@149507.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@149507.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@149507.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@149507.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@149521.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@149521.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@149521.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@149521.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@149521.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@149521.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@149535.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@149535.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@149535.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@149535.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@149535.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@149535.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@149549.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@149549.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@149549.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@149549.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@149549.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@149549.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@149563.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@149563.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@149563.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@149563.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@149563.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@149563.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@149577.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@149577.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@149577.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@149577.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@149577.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@149577.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@149591.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@149591.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@149591.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@149591.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@149591.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@149591.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@149605.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@149605.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@149605.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@149605.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@149605.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@149605.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@149619.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@149619.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@149619.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@149619.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@149619.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@149619.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@149633.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@149633.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@149633.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@149633.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@149633.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@149633.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@149647.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@149647.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@149647.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@149647.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@149647.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@149647.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@149661.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@149661.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@149661.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@149661.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@149661.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@149661.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@149675.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@149675.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@149675.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@149675.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@149675.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@149675.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@149689.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@149689.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@149689.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@149689.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@149689.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@149689.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@149703.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@149703.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@149703.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@149703.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@149703.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@149703.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@149717.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@149717.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@149717.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@149717.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@149717.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@149717.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@149731.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@149731.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@149731.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@149731.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@149731.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@149731.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@149745.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@149745.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@149745.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@149745.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@149745.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@149745.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@149759.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@149759.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@149759.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@149759.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@149759.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@149759.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@149773.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@149773.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@149773.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@149773.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@149773.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@149773.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@149787.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@149787.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@149787.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@149787.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@149787.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@149787.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@149801.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@149801.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@149801.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@149801.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@149801.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@149801.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@149815.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@149815.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@149815.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@149815.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@149815.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@149815.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@149829.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@149829.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@149829.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@149829.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@149829.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@149829.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@149843.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@149843.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@149843.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@149843.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@149843.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@149843.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@149857.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@149857.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@149857.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@149857.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@149857.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@149857.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@149871.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@149871.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@149871.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@149871.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@149871.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@149871.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@149885.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@149885.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@149885.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@149885.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@149885.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@149885.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@149899.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@149899.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@149899.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@149899.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@149899.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@149899.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@149913.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@149913.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@149913.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@149913.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@149913.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@149913.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@149927.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@149927.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@149927.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@149927.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@149927.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@149927.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@149941.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@149941.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@149941.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@149941.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@149941.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@149941.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@149955.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@149955.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@149955.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@149955.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@149955.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@149955.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@149969.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@149969.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@149969.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@149969.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@149969.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@149969.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@149983.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@149983.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@149983.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@149983.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@149983.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@149983.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@149997.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@149997.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@149997.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@149997.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@149997.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@149997.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@150011.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@150011.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@150011.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@150011.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@150011.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@150011.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@150025.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@150025.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@150025.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@150025.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@150025.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@150025.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@150039.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@150039.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@150039.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@150039.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@150039.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@150039.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@150053.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@150053.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@150053.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@150053.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@150053.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@150053.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@150067.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@150067.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@150067.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@150067.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@150067.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@150067.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@150081.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@150081.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@150081.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@150081.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@150081.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@150081.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@150095.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@150095.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@150095.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@150095.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@150095.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@150095.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@150109.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@150109.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@150109.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@150109.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@150109.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@150109.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@150123.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@150123.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@150123.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@150123.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@150123.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@150123.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@150137.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@150137.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@150137.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@150137.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@150137.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@150137.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@150151.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@150151.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@150151.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@150151.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@150151.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@150151.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@150165.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@150165.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@150165.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@150165.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@150165.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@150165.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@150179.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@150179.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@150179.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@150179.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@150179.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@150179.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@150193.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@150193.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@150193.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@150193.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@150193.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@150193.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@150207.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@150207.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@150207.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@150207.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@150207.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@150207.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@150221.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@150221.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@150221.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@150221.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@150221.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@150221.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@150235.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@150235.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@150235.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@150235.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@150235.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@150235.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@150249.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@150249.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@150249.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@150249.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@150249.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@150249.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@150263.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@150263.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@150263.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@150263.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@150263.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@150263.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@150277.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@150277.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@150277.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@150277.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@150277.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@150277.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@150291.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@150291.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@150291.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@150291.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@150291.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@150291.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@150305.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@150305.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@150305.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@150305.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@150305.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@150305.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@150319.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@150319.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@150319.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@150319.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@150319.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@150319.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@150333.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@150333.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@150333.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@150333.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@150333.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@150333.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@150347.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@150347.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@150347.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@150347.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@150347.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@150347.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@150361.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@150361.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@150361.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@150361.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@150361.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@150361.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@150375.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@150375.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@150375.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@150375.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@150375.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@150375.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@150389.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@150389.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@150389.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@150389.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@150389.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@150389.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@150403.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@150403.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@150403.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@150403.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@150403.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@150403.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@150417.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@150417.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@150417.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@150417.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@150417.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@150417.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@150431.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@150431.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@150431.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@150431.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@150431.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@150431.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@150445.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@150445.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@150445.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@150445.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@150445.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@150445.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@150459.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@150459.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@150459.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@150459.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@150459.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@150459.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@150473.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@150473.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@150473.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@150473.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@150473.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@150473.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@150487.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@150487.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@150487.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@150487.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@150487.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@150487.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@150501.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@150501.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@150501.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@150501.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@150501.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@150501.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@150515.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@150515.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@150515.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@150515.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@150515.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@150515.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@150529.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@150529.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@150529.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@150529.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@150529.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@150529.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@150543.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@150543.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@150543.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@150543.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@150543.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@150543.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@150557.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@150557.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@150557.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@150557.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@150557.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@150557.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@150571.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@150571.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@150571.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@150571.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@150571.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@150571.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@150585.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@150585.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@150585.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@150585.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@150585.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@150585.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@150599.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@150599.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@150599.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@150599.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@150599.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@150599.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@150613.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@150613.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@150613.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@150613.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@150613.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@150613.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@150627.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@150627.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@150627.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@150627.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@150627.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@150627.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@150641.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@150641.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@150641.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@150641.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@150641.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@150641.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@150655.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@150655.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@150655.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@150655.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@150655.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@150655.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@150669.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@150669.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@150669.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@150669.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@150669.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@150669.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@150683.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@150683.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@150683.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@150683.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@150683.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@150683.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@150697.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@150697.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@150697.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@150697.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@150697.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@150697.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@150711.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@150711.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@150711.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@150711.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@150711.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@150711.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@150725.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@150725.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@150725.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@150725.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@150725.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@150725.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@150739.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@150739.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@150739.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@150739.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@150739.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@150739.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@150753.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@150753.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@150753.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@150753.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@150753.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@150753.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@150767.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@150767.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@150767.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@150767.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@150767.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@150767.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@150781.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@150781.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@150781.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@150781.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@150781.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@150781.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@150795.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@150795.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@150795.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@150795.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@150795.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@150795.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@150809.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@150809.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@150809.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@150809.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@150809.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@150809.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@150823.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@150823.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@150823.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@150823.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@150823.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@150823.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@150837.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@150837.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@150837.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@150837.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@150837.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@150837.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@150851.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@150851.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@150851.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@150851.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@150851.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@150851.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@150865.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@150865.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@150865.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@150865.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@150865.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@150865.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@150879.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@150879.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@150879.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@150879.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@150879.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@150879.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@150893.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@150893.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@150893.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@150893.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@150893.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@150893.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@150907.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@150907.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@150907.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@150907.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@150907.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@150907.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@150921.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@150921.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@150921.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@150921.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@150921.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@150921.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@150935.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@150935.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@150935.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@150935.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@150935.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@150935.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@150949.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@150949.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@150949.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@150949.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@150949.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@150949.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@150963.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@150963.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@150963.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@150963.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@150963.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@150963.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@150977.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@150977.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@150977.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@150977.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@150977.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@150977.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@150991.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@150991.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@150991.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@150991.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@150991.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@150991.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@151005.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@151005.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@151005.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@151005.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@151005.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@151005.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@151019.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@151019.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@151019.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@151019.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@151019.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@151019.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@151033.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@151033.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@151033.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@151033.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@151033.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@151033.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@151047.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@151047.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@151047.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@151047.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@151047.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@151047.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@151061.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@151061.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@151061.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@151061.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@151061.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@151061.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@151075.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@151075.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@151075.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@151075.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@151075.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@151075.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@151089.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@151089.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@151089.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@151089.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@151089.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@151089.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@151103.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@151103.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@151103.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@151103.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@151103.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@151103.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@151117.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@151117.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@151117.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@151117.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@151117.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@151117.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@151131.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@151131.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@151131.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@151131.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@151131.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@151131.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@151145.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@151145.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@151145.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@151145.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@151145.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@151145.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@151159.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@151159.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@151159.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@151159.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@151159.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@151159.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@151173.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@151173.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@151173.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@151173.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@151173.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@151173.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@151187.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@151187.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@151187.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@151187.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@151187.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@151187.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@151201.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@151201.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@151201.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@151201.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@151201.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@151201.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@151215.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@151215.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@151215.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@151215.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@151215.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@151215.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@151229.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@151229.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@151229.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@151229.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@151229.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@151229.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@151243.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@151243.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@151243.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@151243.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@151243.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@151243.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@151257.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@151257.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@151257.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@151257.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@151257.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@151257.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@151271.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@151271.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@151271.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@151271.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@151271.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@151271.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@151285.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@151285.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@151285.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@151285.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@151285.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@151285.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@151299.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@151299.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@151299.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@151299.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@151299.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@151299.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@151313.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@151313.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@151313.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@151313.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@151313.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@151313.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@151327.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@151327.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@151327.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@151327.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@151327.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@151327.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@151341.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@151341.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@151341.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@151341.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@151341.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@151341.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@151355.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@151355.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@151355.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@151355.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@151355.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@151355.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@151369.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@151369.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@151369.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@151369.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@151369.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@151369.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@151383.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@151383.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@151383.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@151383.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@151383.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@151383.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@151397.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@151397.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@151397.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@151397.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@151397.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@151397.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@151411.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@151411.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@151411.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@151411.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@151411.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@151411.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@151425.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@151425.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@151425.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@151425.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@151425.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@151425.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@151439.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@151439.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@151439.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@151439.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@151439.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@151439.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@151453.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@151453.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@151453.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@151453.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@151453.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@151453.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@151467.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@151467.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@151467.4]
  wire  _T_3078; // @[RegFile.scala 80:42:@144429.4]
  wire  _T_3084; // @[RegFile.scala 68:46:@144441.4]
  wire  _T_3085; // @[RegFile.scala 68:34:@144442.4]
  wire  _T_3098; // @[RegFile.scala 80:42:@144460.4]
  wire  _T_3104; // @[RegFile.scala 80:42:@144472.4]
  wire  _T_3110; // @[RegFile.scala 74:80:@144484.4]
  wire  _T_3111; // @[RegFile.scala 74:68:@144485.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@144426.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@144438.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@144457.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@144469.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@144481.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@144495.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@144509.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@144523.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@144537.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@144551.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@144565.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@144579.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@144593.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@144607.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@144621.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@144635.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@144649.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@144663.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@144677.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@144691.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@144705.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@144719.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@144733.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@144747.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@144761.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@144775.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@144789.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@144803.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@144817.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@144831.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@144845.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@144859.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@144873.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@144887.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@144901.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@144915.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@144929.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@144943.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@144957.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@144971.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@144985.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@144999.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@145013.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@145027.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@145041.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@145055.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@145069.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@145083.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@145097.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@145111.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@145125.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@145139.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@145153.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@145167.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@145181.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@145195.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@145209.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@145223.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@145237.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@145251.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@145265.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@145279.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@145293.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@145307.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@145321.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@145335.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@145349.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@145363.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@145377.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@145391.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@145405.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@145419.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@145433.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@145447.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@145461.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@145475.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@145489.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@145503.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@145517.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@145531.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@145545.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@145559.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@145573.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@145587.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@145601.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@145615.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@145629.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@145643.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@145657.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@145671.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@145685.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@145699.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@145713.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@145727.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@145741.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@145755.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@145769.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@145783.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@145797.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@145811.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@145825.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@145839.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@145853.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@145867.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@145881.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@145895.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@145909.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@145923.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@145937.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@145951.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@145965.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@145979.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@145993.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@146007.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@146021.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@146035.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@146049.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@146063.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@146077.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@146091.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@146105.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@146119.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@146133.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@146147.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@146161.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@146175.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@146189.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@146203.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@146217.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@146231.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@146245.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@146259.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@146273.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@146287.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@146301.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@146315.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@146329.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@146343.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@146357.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@146371.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@146385.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@146399.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@146413.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@146427.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@146441.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@146455.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@146469.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@146483.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@146497.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@146511.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@146525.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@146539.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@146553.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@146567.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@146581.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@146595.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@146609.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@146623.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@146637.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@146651.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@146665.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@146679.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@146693.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@146707.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@146721.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@146735.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@146749.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@146763.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@146777.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@146791.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@146805.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@146819.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@146833.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@146847.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@146861.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@146875.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@146889.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@146903.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@146917.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@146931.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@146945.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@146959.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@146973.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@146987.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@147001.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@147015.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@147029.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@147043.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@147057.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@147071.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@147085.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@147099.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@147113.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@147127.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@147141.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@147155.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@147169.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@147183.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@147197.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@147211.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@147225.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@147239.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@147253.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@147267.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@147281.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@147295.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@147309.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@147323.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@147337.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@147351.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@147365.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@147379.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@147393.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@147407.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@147421.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@147435.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@147449.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@147463.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@147477.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@147491.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@147505.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@147519.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@147533.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@147547.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@147561.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@147575.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@147589.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@147603.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@147617.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@147631.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@147645.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@147659.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@147673.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@147687.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@147701.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@147715.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@147729.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@147743.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@147757.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@147771.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@147785.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@147799.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@147813.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@147827.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@147841.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@147855.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@147869.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@147883.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@147897.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@147911.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@147925.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@147939.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@147953.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@147967.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@147981.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@147995.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@148009.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@148023.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@148037.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@148051.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@148065.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@148079.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@148093.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@148107.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@148121.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@148135.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@148149.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@148163.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@148177.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@148191.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@148205.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@148219.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@148233.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@148247.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@148261.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@148275.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@148289.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@148303.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@148317.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@148331.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@148345.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@148359.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@148373.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@148387.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@148401.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@148415.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@148429.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@148443.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@148457.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@148471.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@148485.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@148499.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@148513.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@148527.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@148541.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@148555.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@148569.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@148583.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@148597.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@148611.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@148625.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@148639.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@148653.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@148667.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@148681.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@148695.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@148709.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@148723.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@148737.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@148751.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@148765.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@148779.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@148793.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@148807.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@148821.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@148835.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@148849.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@148863.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@148877.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@148891.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@148905.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@148919.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@148933.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@148947.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@148961.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@148975.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@148989.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@149003.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@149017.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@149031.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@149045.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@149059.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@149073.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@149087.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@149101.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@149115.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@149129.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@149143.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@149157.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@149171.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@149185.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@149199.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@149213.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@149227.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@149241.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@149255.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@149269.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@149283.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@149297.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@149311.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@149325.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@149339.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@149353.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@149367.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@149381.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@149395.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@149409.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@149423.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@149437.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@149451.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@149465.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@149479.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@149493.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@149507.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@149521.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@149535.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@149549.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@149563.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@149577.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@149591.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@149605.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@149619.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@149633.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@149647.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@149661.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@149675.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@149689.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@149703.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@149717.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@149731.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@149745.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@149759.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@149773.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@149787.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@149801.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@149815.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@149829.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@149843.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@149857.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@149871.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@149885.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@149899.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@149913.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@149927.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@149941.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@149955.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@149969.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@149983.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@149997.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@150011.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@150025.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@150039.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@150053.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@150067.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@150081.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@150095.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@150109.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@150123.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@150137.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@150151.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@150165.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@150179.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@150193.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@150207.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@150221.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@150235.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@150249.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@150263.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@150277.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@150291.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@150305.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@150319.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@150333.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@150347.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@150361.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@150375.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@150389.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@150403.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@150417.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@150431.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@150445.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@150459.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@150473.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@150487.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@150501.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@150515.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@150529.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@150543.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@150557.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@150571.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@150585.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@150599.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@150613.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@150627.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@150641.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@150655.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@150669.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@150683.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@150697.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@150711.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@150725.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@150739.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@150753.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@150767.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@150781.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@150795.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@150809.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@150823.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@150837.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@150851.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@150865.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@150879.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@150893.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@150907.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@150921.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@150935.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@150949.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@150963.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@150977.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@150991.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@151005.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@151019.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@151033.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@151047.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@151061.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@151075.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@151089.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@151103.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@151117.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@151131.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@151145.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@151159.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@151173.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@151187.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@151201.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@151215.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@151229.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@151243.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@151257.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@151271.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@151285.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@151299.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@151313.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@151327.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@151341.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@151355.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@151369.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@151383.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@151397.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@151411.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@151425.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@151439.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@151453.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@151467.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3078 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@144429.4]
  assign _T_3084 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@144441.4]
  assign _T_3085 = io_wen & _T_3084; // @[RegFile.scala 68:34:@144442.4]
  assign _T_3098 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@144460.4]
  assign _T_3104 = io_waddr == 32'h3; // @[RegFile.scala 80:42:@144472.4]
  assign _T_3110 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@144484.4]
  assign _T_3111 = io_wen & _T_3110; // @[RegFile.scala 74:68:@144485.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@152478.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@152484.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@152485.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@152486.4]
  assign io_argIns_3 = regs_3_io_out; // @[RegFile.scala 111:13:@152487.4]
  assign regs_0_clock = clock; // @[:@144427.4]
  assign regs_0_reset = reset; // @[:@144428.4 RegFile.scala 82:16:@144434.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@144432.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@144436.4]
  assign regs_0_io_enable = io_wen & _T_3078; // @[RegFile.scala 80:20:@144431.4]
  assign regs_1_clock = clock; // @[:@144439.4]
  assign regs_1_reset = reset; // @[:@144440.4 RegFile.scala 70:16:@144452.4]
  assign regs_1_io_in = _T_3085 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@144450.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@144455.4]
  assign regs_1_io_enable = _T_3085 ? _T_3085 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@144446.4]
  assign regs_2_clock = clock; // @[:@144458.4]
  assign regs_2_reset = reset; // @[:@144459.4 RegFile.scala 82:16:@144465.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@144463.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@144467.4]
  assign regs_2_io_enable = io_wen & _T_3098; // @[RegFile.scala 80:20:@144462.4]
  assign regs_3_clock = clock; // @[:@144470.4]
  assign regs_3_reset = reset; // @[:@144471.4 RegFile.scala 82:16:@144477.4]
  assign regs_3_io_in = io_wdata; // @[RegFile.scala 81:16:@144475.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 83:19:@144479.4]
  assign regs_3_io_enable = io_wen & _T_3104; // @[RegFile.scala 80:20:@144474.4]
  assign regs_4_clock = clock; // @[:@144482.4]
  assign regs_4_reset = io_reset; // @[:@144483.4 RegFile.scala 76:16:@144490.4]
  assign regs_4_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@144489.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@144493.4]
  assign regs_4_io_enable = io_argOuts_1_valid | _T_3111; // @[RegFile.scala 74:20:@144487.4]
  assign regs_5_clock = clock; // @[:@144496.4]
  assign regs_5_reset = io_reset; // @[:@144497.4 RegFile.scala 76:16:@144504.4]
  assign regs_5_io_in = 64'h0; // @[RegFile.scala 75:16:@144503.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@144507.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 74:20:@144501.4]
  assign regs_6_clock = clock; // @[:@144510.4]
  assign regs_6_reset = io_reset; // @[:@144511.4 RegFile.scala 76:16:@144518.4]
  assign regs_6_io_in = 64'h0; // @[RegFile.scala 75:16:@144517.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@144521.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 74:20:@144515.4]
  assign regs_7_clock = clock; // @[:@144524.4]
  assign regs_7_reset = io_reset; // @[:@144525.4 RegFile.scala 76:16:@144532.4]
  assign regs_7_io_in = 64'h0; // @[RegFile.scala 75:16:@144531.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@144535.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 74:20:@144529.4]
  assign regs_8_clock = clock; // @[:@144538.4]
  assign regs_8_reset = io_reset; // @[:@144539.4 RegFile.scala 76:16:@144546.4]
  assign regs_8_io_in = 64'h0; // @[RegFile.scala 75:16:@144545.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@144549.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 74:20:@144543.4]
  assign regs_9_clock = clock; // @[:@144552.4]
  assign regs_9_reset = io_reset; // @[:@144553.4 RegFile.scala 76:16:@144560.4]
  assign regs_9_io_in = 64'h0; // @[RegFile.scala 75:16:@144559.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@144563.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 74:20:@144557.4]
  assign regs_10_clock = clock; // @[:@144566.4]
  assign regs_10_reset = io_reset; // @[:@144567.4 RegFile.scala 76:16:@144574.4]
  assign regs_10_io_in = 64'h0; // @[RegFile.scala 75:16:@144573.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@144577.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 74:20:@144571.4]
  assign regs_11_clock = clock; // @[:@144580.4]
  assign regs_11_reset = io_reset; // @[:@144581.4 RegFile.scala 76:16:@144588.4]
  assign regs_11_io_in = 64'h0; // @[RegFile.scala 75:16:@144587.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@144591.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 74:20:@144585.4]
  assign regs_12_clock = clock; // @[:@144594.4]
  assign regs_12_reset = io_reset; // @[:@144595.4 RegFile.scala 76:16:@144602.4]
  assign regs_12_io_in = 64'h0; // @[RegFile.scala 75:16:@144601.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@144605.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 74:20:@144599.4]
  assign regs_13_clock = clock; // @[:@144608.4]
  assign regs_13_reset = io_reset; // @[:@144609.4 RegFile.scala 76:16:@144616.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 75:16:@144615.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@144619.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@144613.4]
  assign regs_14_clock = clock; // @[:@144622.4]
  assign regs_14_reset = io_reset; // @[:@144623.4 RegFile.scala 76:16:@144630.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 75:16:@144629.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@144633.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@144627.4]
  assign regs_15_clock = clock; // @[:@144636.4]
  assign regs_15_reset = io_reset; // @[:@144637.4 RegFile.scala 76:16:@144644.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 75:16:@144643.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@144647.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@144641.4]
  assign regs_16_clock = clock; // @[:@144650.4]
  assign regs_16_reset = io_reset; // @[:@144651.4 RegFile.scala 76:16:@144658.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 75:16:@144657.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@144661.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@144655.4]
  assign regs_17_clock = clock; // @[:@144664.4]
  assign regs_17_reset = io_reset; // @[:@144665.4 RegFile.scala 76:16:@144672.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 75:16:@144671.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@144675.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@144669.4]
  assign regs_18_clock = clock; // @[:@144678.4]
  assign regs_18_reset = io_reset; // @[:@144679.4 RegFile.scala 76:16:@144686.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 75:16:@144685.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@144689.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@144683.4]
  assign regs_19_clock = clock; // @[:@144692.4]
  assign regs_19_reset = io_reset; // @[:@144693.4 RegFile.scala 76:16:@144700.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 75:16:@144699.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@144703.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@144697.4]
  assign regs_20_clock = clock; // @[:@144706.4]
  assign regs_20_reset = io_reset; // @[:@144707.4 RegFile.scala 76:16:@144714.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 75:16:@144713.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@144717.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@144711.4]
  assign regs_21_clock = clock; // @[:@144720.4]
  assign regs_21_reset = io_reset; // @[:@144721.4 RegFile.scala 76:16:@144728.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 75:16:@144727.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@144731.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@144725.4]
  assign regs_22_clock = clock; // @[:@144734.4]
  assign regs_22_reset = io_reset; // @[:@144735.4 RegFile.scala 76:16:@144742.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 75:16:@144741.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@144745.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@144739.4]
  assign regs_23_clock = clock; // @[:@144748.4]
  assign regs_23_reset = io_reset; // @[:@144749.4 RegFile.scala 76:16:@144756.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@144755.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@144759.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@144753.4]
  assign regs_24_clock = clock; // @[:@144762.4]
  assign regs_24_reset = io_reset; // @[:@144763.4 RegFile.scala 76:16:@144770.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@144769.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@144773.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@144767.4]
  assign regs_25_clock = clock; // @[:@144776.4]
  assign regs_25_reset = io_reset; // @[:@144777.4 RegFile.scala 76:16:@144784.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@144783.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@144787.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@144781.4]
  assign regs_26_clock = clock; // @[:@144790.4]
  assign regs_26_reset = io_reset; // @[:@144791.4 RegFile.scala 76:16:@144798.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@144797.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@144801.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@144795.4]
  assign regs_27_clock = clock; // @[:@144804.4]
  assign regs_27_reset = io_reset; // @[:@144805.4 RegFile.scala 76:16:@144812.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@144811.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@144815.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@144809.4]
  assign regs_28_clock = clock; // @[:@144818.4]
  assign regs_28_reset = io_reset; // @[:@144819.4 RegFile.scala 76:16:@144826.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@144825.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@144829.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@144823.4]
  assign regs_29_clock = clock; // @[:@144832.4]
  assign regs_29_reset = io_reset; // @[:@144833.4 RegFile.scala 76:16:@144840.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@144839.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@144843.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@144837.4]
  assign regs_30_clock = clock; // @[:@144846.4]
  assign regs_30_reset = io_reset; // @[:@144847.4 RegFile.scala 76:16:@144854.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@144853.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@144857.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@144851.4]
  assign regs_31_clock = clock; // @[:@144860.4]
  assign regs_31_reset = io_reset; // @[:@144861.4 RegFile.scala 76:16:@144868.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@144867.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@144871.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@144865.4]
  assign regs_32_clock = clock; // @[:@144874.4]
  assign regs_32_reset = io_reset; // @[:@144875.4 RegFile.scala 76:16:@144882.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@144881.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@144885.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@144879.4]
  assign regs_33_clock = clock; // @[:@144888.4]
  assign regs_33_reset = io_reset; // @[:@144889.4 RegFile.scala 76:16:@144896.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@144895.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@144899.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@144893.4]
  assign regs_34_clock = clock; // @[:@144902.4]
  assign regs_34_reset = io_reset; // @[:@144903.4 RegFile.scala 76:16:@144910.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@144909.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@144913.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@144907.4]
  assign regs_35_clock = clock; // @[:@144916.4]
  assign regs_35_reset = io_reset; // @[:@144917.4 RegFile.scala 76:16:@144924.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@144923.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@144927.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@144921.4]
  assign regs_36_clock = clock; // @[:@144930.4]
  assign regs_36_reset = io_reset; // @[:@144931.4 RegFile.scala 76:16:@144938.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@144937.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@144941.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@144935.4]
  assign regs_37_clock = clock; // @[:@144944.4]
  assign regs_37_reset = io_reset; // @[:@144945.4 RegFile.scala 76:16:@144952.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@144951.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@144955.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@144949.4]
  assign regs_38_clock = clock; // @[:@144958.4]
  assign regs_38_reset = io_reset; // @[:@144959.4 RegFile.scala 76:16:@144966.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@144965.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@144969.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@144963.4]
  assign regs_39_clock = clock; // @[:@144972.4]
  assign regs_39_reset = io_reset; // @[:@144973.4 RegFile.scala 76:16:@144980.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@144979.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@144983.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@144977.4]
  assign regs_40_clock = clock; // @[:@144986.4]
  assign regs_40_reset = io_reset; // @[:@144987.4 RegFile.scala 76:16:@144994.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@144993.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@144997.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@144991.4]
  assign regs_41_clock = clock; // @[:@145000.4]
  assign regs_41_reset = io_reset; // @[:@145001.4 RegFile.scala 76:16:@145008.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@145007.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@145011.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@145005.4]
  assign regs_42_clock = clock; // @[:@145014.4]
  assign regs_42_reset = io_reset; // @[:@145015.4 RegFile.scala 76:16:@145022.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@145021.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@145025.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@145019.4]
  assign regs_43_clock = clock; // @[:@145028.4]
  assign regs_43_reset = io_reset; // @[:@145029.4 RegFile.scala 76:16:@145036.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@145035.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@145039.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@145033.4]
  assign regs_44_clock = clock; // @[:@145042.4]
  assign regs_44_reset = io_reset; // @[:@145043.4 RegFile.scala 76:16:@145050.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@145049.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@145053.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@145047.4]
  assign regs_45_clock = clock; // @[:@145056.4]
  assign regs_45_reset = io_reset; // @[:@145057.4 RegFile.scala 76:16:@145064.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@145063.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@145067.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@145061.4]
  assign regs_46_clock = clock; // @[:@145070.4]
  assign regs_46_reset = io_reset; // @[:@145071.4 RegFile.scala 76:16:@145078.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@145077.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@145081.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@145075.4]
  assign regs_47_clock = clock; // @[:@145084.4]
  assign regs_47_reset = io_reset; // @[:@145085.4 RegFile.scala 76:16:@145092.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@145091.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@145095.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@145089.4]
  assign regs_48_clock = clock; // @[:@145098.4]
  assign regs_48_reset = io_reset; // @[:@145099.4 RegFile.scala 76:16:@145106.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@145105.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@145109.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@145103.4]
  assign regs_49_clock = clock; // @[:@145112.4]
  assign regs_49_reset = io_reset; // @[:@145113.4 RegFile.scala 76:16:@145120.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@145119.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@145123.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@145117.4]
  assign regs_50_clock = clock; // @[:@145126.4]
  assign regs_50_reset = io_reset; // @[:@145127.4 RegFile.scala 76:16:@145134.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@145133.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@145137.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@145131.4]
  assign regs_51_clock = clock; // @[:@145140.4]
  assign regs_51_reset = io_reset; // @[:@145141.4 RegFile.scala 76:16:@145148.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@145147.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@145151.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@145145.4]
  assign regs_52_clock = clock; // @[:@145154.4]
  assign regs_52_reset = io_reset; // @[:@145155.4 RegFile.scala 76:16:@145162.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@145161.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@145165.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@145159.4]
  assign regs_53_clock = clock; // @[:@145168.4]
  assign regs_53_reset = io_reset; // @[:@145169.4 RegFile.scala 76:16:@145176.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@145175.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@145179.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@145173.4]
  assign regs_54_clock = clock; // @[:@145182.4]
  assign regs_54_reset = io_reset; // @[:@145183.4 RegFile.scala 76:16:@145190.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@145189.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@145193.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@145187.4]
  assign regs_55_clock = clock; // @[:@145196.4]
  assign regs_55_reset = io_reset; // @[:@145197.4 RegFile.scala 76:16:@145204.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@145203.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@145207.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@145201.4]
  assign regs_56_clock = clock; // @[:@145210.4]
  assign regs_56_reset = io_reset; // @[:@145211.4 RegFile.scala 76:16:@145218.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@145217.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@145221.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@145215.4]
  assign regs_57_clock = clock; // @[:@145224.4]
  assign regs_57_reset = io_reset; // @[:@145225.4 RegFile.scala 76:16:@145232.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@145231.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@145235.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@145229.4]
  assign regs_58_clock = clock; // @[:@145238.4]
  assign regs_58_reset = io_reset; // @[:@145239.4 RegFile.scala 76:16:@145246.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@145245.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@145249.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@145243.4]
  assign regs_59_clock = clock; // @[:@145252.4]
  assign regs_59_reset = io_reset; // @[:@145253.4 RegFile.scala 76:16:@145260.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@145259.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@145263.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@145257.4]
  assign regs_60_clock = clock; // @[:@145266.4]
  assign regs_60_reset = io_reset; // @[:@145267.4 RegFile.scala 76:16:@145274.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@145273.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@145277.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@145271.4]
  assign regs_61_clock = clock; // @[:@145280.4]
  assign regs_61_reset = io_reset; // @[:@145281.4 RegFile.scala 76:16:@145288.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@145287.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@145291.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@145285.4]
  assign regs_62_clock = clock; // @[:@145294.4]
  assign regs_62_reset = io_reset; // @[:@145295.4 RegFile.scala 76:16:@145302.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@145301.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@145305.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@145299.4]
  assign regs_63_clock = clock; // @[:@145308.4]
  assign regs_63_reset = io_reset; // @[:@145309.4 RegFile.scala 76:16:@145316.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@145315.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@145319.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@145313.4]
  assign regs_64_clock = clock; // @[:@145322.4]
  assign regs_64_reset = io_reset; // @[:@145323.4 RegFile.scala 76:16:@145330.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@145329.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@145333.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@145327.4]
  assign regs_65_clock = clock; // @[:@145336.4]
  assign regs_65_reset = io_reset; // @[:@145337.4 RegFile.scala 76:16:@145344.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@145343.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@145347.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@145341.4]
  assign regs_66_clock = clock; // @[:@145350.4]
  assign regs_66_reset = io_reset; // @[:@145351.4 RegFile.scala 76:16:@145358.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@145357.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@145361.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@145355.4]
  assign regs_67_clock = clock; // @[:@145364.4]
  assign regs_67_reset = io_reset; // @[:@145365.4 RegFile.scala 76:16:@145372.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@145371.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@145375.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@145369.4]
  assign regs_68_clock = clock; // @[:@145378.4]
  assign regs_68_reset = io_reset; // @[:@145379.4 RegFile.scala 76:16:@145386.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@145385.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@145389.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@145383.4]
  assign regs_69_clock = clock; // @[:@145392.4]
  assign regs_69_reset = io_reset; // @[:@145393.4 RegFile.scala 76:16:@145400.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@145399.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@145403.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@145397.4]
  assign regs_70_clock = clock; // @[:@145406.4]
  assign regs_70_reset = io_reset; // @[:@145407.4 RegFile.scala 76:16:@145414.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@145413.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@145417.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@145411.4]
  assign regs_71_clock = clock; // @[:@145420.4]
  assign regs_71_reset = io_reset; // @[:@145421.4 RegFile.scala 76:16:@145428.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@145427.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@145431.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@145425.4]
  assign regs_72_clock = clock; // @[:@145434.4]
  assign regs_72_reset = io_reset; // @[:@145435.4 RegFile.scala 76:16:@145442.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@145441.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@145445.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@145439.4]
  assign regs_73_clock = clock; // @[:@145448.4]
  assign regs_73_reset = io_reset; // @[:@145449.4 RegFile.scala 76:16:@145456.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@145455.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@145459.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@145453.4]
  assign regs_74_clock = clock; // @[:@145462.4]
  assign regs_74_reset = io_reset; // @[:@145463.4 RegFile.scala 76:16:@145470.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@145469.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@145473.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@145467.4]
  assign regs_75_clock = clock; // @[:@145476.4]
  assign regs_75_reset = io_reset; // @[:@145477.4 RegFile.scala 76:16:@145484.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@145483.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@145487.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@145481.4]
  assign regs_76_clock = clock; // @[:@145490.4]
  assign regs_76_reset = io_reset; // @[:@145491.4 RegFile.scala 76:16:@145498.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@145497.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@145501.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@145495.4]
  assign regs_77_clock = clock; // @[:@145504.4]
  assign regs_77_reset = io_reset; // @[:@145505.4 RegFile.scala 76:16:@145512.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@145511.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@145515.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@145509.4]
  assign regs_78_clock = clock; // @[:@145518.4]
  assign regs_78_reset = io_reset; // @[:@145519.4 RegFile.scala 76:16:@145526.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@145525.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@145529.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@145523.4]
  assign regs_79_clock = clock; // @[:@145532.4]
  assign regs_79_reset = io_reset; // @[:@145533.4 RegFile.scala 76:16:@145540.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@145539.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@145543.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@145537.4]
  assign regs_80_clock = clock; // @[:@145546.4]
  assign regs_80_reset = io_reset; // @[:@145547.4 RegFile.scala 76:16:@145554.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@145553.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@145557.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@145551.4]
  assign regs_81_clock = clock; // @[:@145560.4]
  assign regs_81_reset = io_reset; // @[:@145561.4 RegFile.scala 76:16:@145568.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@145567.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@145571.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@145565.4]
  assign regs_82_clock = clock; // @[:@145574.4]
  assign regs_82_reset = io_reset; // @[:@145575.4 RegFile.scala 76:16:@145582.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@145581.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@145585.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@145579.4]
  assign regs_83_clock = clock; // @[:@145588.4]
  assign regs_83_reset = io_reset; // @[:@145589.4 RegFile.scala 76:16:@145596.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@145595.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@145599.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@145593.4]
  assign regs_84_clock = clock; // @[:@145602.4]
  assign regs_84_reset = io_reset; // @[:@145603.4 RegFile.scala 76:16:@145610.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@145609.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@145613.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@145607.4]
  assign regs_85_clock = clock; // @[:@145616.4]
  assign regs_85_reset = io_reset; // @[:@145617.4 RegFile.scala 76:16:@145624.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@145623.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@145627.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@145621.4]
  assign regs_86_clock = clock; // @[:@145630.4]
  assign regs_86_reset = io_reset; // @[:@145631.4 RegFile.scala 76:16:@145638.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@145637.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@145641.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@145635.4]
  assign regs_87_clock = clock; // @[:@145644.4]
  assign regs_87_reset = io_reset; // @[:@145645.4 RegFile.scala 76:16:@145652.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@145651.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@145655.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@145649.4]
  assign regs_88_clock = clock; // @[:@145658.4]
  assign regs_88_reset = io_reset; // @[:@145659.4 RegFile.scala 76:16:@145666.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@145665.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@145669.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@145663.4]
  assign regs_89_clock = clock; // @[:@145672.4]
  assign regs_89_reset = io_reset; // @[:@145673.4 RegFile.scala 76:16:@145680.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@145679.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@145683.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@145677.4]
  assign regs_90_clock = clock; // @[:@145686.4]
  assign regs_90_reset = io_reset; // @[:@145687.4 RegFile.scala 76:16:@145694.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@145693.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@145697.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@145691.4]
  assign regs_91_clock = clock; // @[:@145700.4]
  assign regs_91_reset = io_reset; // @[:@145701.4 RegFile.scala 76:16:@145708.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@145707.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@145711.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@145705.4]
  assign regs_92_clock = clock; // @[:@145714.4]
  assign regs_92_reset = io_reset; // @[:@145715.4 RegFile.scala 76:16:@145722.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@145721.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@145725.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@145719.4]
  assign regs_93_clock = clock; // @[:@145728.4]
  assign regs_93_reset = io_reset; // @[:@145729.4 RegFile.scala 76:16:@145736.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@145735.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@145739.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@145733.4]
  assign regs_94_clock = clock; // @[:@145742.4]
  assign regs_94_reset = io_reset; // @[:@145743.4 RegFile.scala 76:16:@145750.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@145749.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@145753.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@145747.4]
  assign regs_95_clock = clock; // @[:@145756.4]
  assign regs_95_reset = io_reset; // @[:@145757.4 RegFile.scala 76:16:@145764.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@145763.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@145767.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@145761.4]
  assign regs_96_clock = clock; // @[:@145770.4]
  assign regs_96_reset = io_reset; // @[:@145771.4 RegFile.scala 76:16:@145778.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@145777.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@145781.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@145775.4]
  assign regs_97_clock = clock; // @[:@145784.4]
  assign regs_97_reset = io_reset; // @[:@145785.4 RegFile.scala 76:16:@145792.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@145791.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@145795.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@145789.4]
  assign regs_98_clock = clock; // @[:@145798.4]
  assign regs_98_reset = io_reset; // @[:@145799.4 RegFile.scala 76:16:@145806.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@145805.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@145809.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@145803.4]
  assign regs_99_clock = clock; // @[:@145812.4]
  assign regs_99_reset = io_reset; // @[:@145813.4 RegFile.scala 76:16:@145820.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@145819.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@145823.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@145817.4]
  assign regs_100_clock = clock; // @[:@145826.4]
  assign regs_100_reset = io_reset; // @[:@145827.4 RegFile.scala 76:16:@145834.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@145833.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@145837.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@145831.4]
  assign regs_101_clock = clock; // @[:@145840.4]
  assign regs_101_reset = io_reset; // @[:@145841.4 RegFile.scala 76:16:@145848.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@145847.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@145851.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@145845.4]
  assign regs_102_clock = clock; // @[:@145854.4]
  assign regs_102_reset = io_reset; // @[:@145855.4 RegFile.scala 76:16:@145862.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@145861.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@145865.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@145859.4]
  assign regs_103_clock = clock; // @[:@145868.4]
  assign regs_103_reset = io_reset; // @[:@145869.4 RegFile.scala 76:16:@145876.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@145875.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@145879.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@145873.4]
  assign regs_104_clock = clock; // @[:@145882.4]
  assign regs_104_reset = io_reset; // @[:@145883.4 RegFile.scala 76:16:@145890.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@145889.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@145893.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@145887.4]
  assign regs_105_clock = clock; // @[:@145896.4]
  assign regs_105_reset = io_reset; // @[:@145897.4 RegFile.scala 76:16:@145904.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@145903.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@145907.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@145901.4]
  assign regs_106_clock = clock; // @[:@145910.4]
  assign regs_106_reset = io_reset; // @[:@145911.4 RegFile.scala 76:16:@145918.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@145917.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@145921.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@145915.4]
  assign regs_107_clock = clock; // @[:@145924.4]
  assign regs_107_reset = io_reset; // @[:@145925.4 RegFile.scala 76:16:@145932.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@145931.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@145935.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@145929.4]
  assign regs_108_clock = clock; // @[:@145938.4]
  assign regs_108_reset = io_reset; // @[:@145939.4 RegFile.scala 76:16:@145946.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@145945.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@145949.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@145943.4]
  assign regs_109_clock = clock; // @[:@145952.4]
  assign regs_109_reset = io_reset; // @[:@145953.4 RegFile.scala 76:16:@145960.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@145959.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@145963.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@145957.4]
  assign regs_110_clock = clock; // @[:@145966.4]
  assign regs_110_reset = io_reset; // @[:@145967.4 RegFile.scala 76:16:@145974.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@145973.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@145977.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@145971.4]
  assign regs_111_clock = clock; // @[:@145980.4]
  assign regs_111_reset = io_reset; // @[:@145981.4 RegFile.scala 76:16:@145988.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@145987.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@145991.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@145985.4]
  assign regs_112_clock = clock; // @[:@145994.4]
  assign regs_112_reset = io_reset; // @[:@145995.4 RegFile.scala 76:16:@146002.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@146001.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@146005.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@145999.4]
  assign regs_113_clock = clock; // @[:@146008.4]
  assign regs_113_reset = io_reset; // @[:@146009.4 RegFile.scala 76:16:@146016.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@146015.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@146019.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@146013.4]
  assign regs_114_clock = clock; // @[:@146022.4]
  assign regs_114_reset = io_reset; // @[:@146023.4 RegFile.scala 76:16:@146030.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@146029.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@146033.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@146027.4]
  assign regs_115_clock = clock; // @[:@146036.4]
  assign regs_115_reset = io_reset; // @[:@146037.4 RegFile.scala 76:16:@146044.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@146043.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@146047.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@146041.4]
  assign regs_116_clock = clock; // @[:@146050.4]
  assign regs_116_reset = io_reset; // @[:@146051.4 RegFile.scala 76:16:@146058.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@146057.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@146061.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@146055.4]
  assign regs_117_clock = clock; // @[:@146064.4]
  assign regs_117_reset = io_reset; // @[:@146065.4 RegFile.scala 76:16:@146072.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@146071.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@146075.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@146069.4]
  assign regs_118_clock = clock; // @[:@146078.4]
  assign regs_118_reset = io_reset; // @[:@146079.4 RegFile.scala 76:16:@146086.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@146085.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@146089.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@146083.4]
  assign regs_119_clock = clock; // @[:@146092.4]
  assign regs_119_reset = io_reset; // @[:@146093.4 RegFile.scala 76:16:@146100.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@146099.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@146103.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@146097.4]
  assign regs_120_clock = clock; // @[:@146106.4]
  assign regs_120_reset = io_reset; // @[:@146107.4 RegFile.scala 76:16:@146114.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@146113.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@146117.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@146111.4]
  assign regs_121_clock = clock; // @[:@146120.4]
  assign regs_121_reset = io_reset; // @[:@146121.4 RegFile.scala 76:16:@146128.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@146127.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@146131.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@146125.4]
  assign regs_122_clock = clock; // @[:@146134.4]
  assign regs_122_reset = io_reset; // @[:@146135.4 RegFile.scala 76:16:@146142.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@146141.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@146145.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@146139.4]
  assign regs_123_clock = clock; // @[:@146148.4]
  assign regs_123_reset = io_reset; // @[:@146149.4 RegFile.scala 76:16:@146156.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@146155.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@146159.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@146153.4]
  assign regs_124_clock = clock; // @[:@146162.4]
  assign regs_124_reset = io_reset; // @[:@146163.4 RegFile.scala 76:16:@146170.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@146169.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@146173.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@146167.4]
  assign regs_125_clock = clock; // @[:@146176.4]
  assign regs_125_reset = io_reset; // @[:@146177.4 RegFile.scala 76:16:@146184.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@146183.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@146187.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@146181.4]
  assign regs_126_clock = clock; // @[:@146190.4]
  assign regs_126_reset = io_reset; // @[:@146191.4 RegFile.scala 76:16:@146198.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@146197.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@146201.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@146195.4]
  assign regs_127_clock = clock; // @[:@146204.4]
  assign regs_127_reset = io_reset; // @[:@146205.4 RegFile.scala 76:16:@146212.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@146211.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@146215.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@146209.4]
  assign regs_128_clock = clock; // @[:@146218.4]
  assign regs_128_reset = io_reset; // @[:@146219.4 RegFile.scala 76:16:@146226.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@146225.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@146229.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@146223.4]
  assign regs_129_clock = clock; // @[:@146232.4]
  assign regs_129_reset = io_reset; // @[:@146233.4 RegFile.scala 76:16:@146240.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@146239.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@146243.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@146237.4]
  assign regs_130_clock = clock; // @[:@146246.4]
  assign regs_130_reset = io_reset; // @[:@146247.4 RegFile.scala 76:16:@146254.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@146253.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@146257.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@146251.4]
  assign regs_131_clock = clock; // @[:@146260.4]
  assign regs_131_reset = io_reset; // @[:@146261.4 RegFile.scala 76:16:@146268.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@146267.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@146271.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@146265.4]
  assign regs_132_clock = clock; // @[:@146274.4]
  assign regs_132_reset = io_reset; // @[:@146275.4 RegFile.scala 76:16:@146282.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@146281.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@146285.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@146279.4]
  assign regs_133_clock = clock; // @[:@146288.4]
  assign regs_133_reset = io_reset; // @[:@146289.4 RegFile.scala 76:16:@146296.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@146295.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@146299.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@146293.4]
  assign regs_134_clock = clock; // @[:@146302.4]
  assign regs_134_reset = io_reset; // @[:@146303.4 RegFile.scala 76:16:@146310.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@146309.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@146313.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@146307.4]
  assign regs_135_clock = clock; // @[:@146316.4]
  assign regs_135_reset = io_reset; // @[:@146317.4 RegFile.scala 76:16:@146324.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@146323.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@146327.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@146321.4]
  assign regs_136_clock = clock; // @[:@146330.4]
  assign regs_136_reset = io_reset; // @[:@146331.4 RegFile.scala 76:16:@146338.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@146337.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@146341.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@146335.4]
  assign regs_137_clock = clock; // @[:@146344.4]
  assign regs_137_reset = io_reset; // @[:@146345.4 RegFile.scala 76:16:@146352.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@146351.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@146355.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@146349.4]
  assign regs_138_clock = clock; // @[:@146358.4]
  assign regs_138_reset = io_reset; // @[:@146359.4 RegFile.scala 76:16:@146366.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@146365.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@146369.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@146363.4]
  assign regs_139_clock = clock; // @[:@146372.4]
  assign regs_139_reset = io_reset; // @[:@146373.4 RegFile.scala 76:16:@146380.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@146379.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@146383.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@146377.4]
  assign regs_140_clock = clock; // @[:@146386.4]
  assign regs_140_reset = io_reset; // @[:@146387.4 RegFile.scala 76:16:@146394.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@146393.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@146397.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@146391.4]
  assign regs_141_clock = clock; // @[:@146400.4]
  assign regs_141_reset = io_reset; // @[:@146401.4 RegFile.scala 76:16:@146408.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@146407.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@146411.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@146405.4]
  assign regs_142_clock = clock; // @[:@146414.4]
  assign regs_142_reset = io_reset; // @[:@146415.4 RegFile.scala 76:16:@146422.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@146421.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@146425.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@146419.4]
  assign regs_143_clock = clock; // @[:@146428.4]
  assign regs_143_reset = io_reset; // @[:@146429.4 RegFile.scala 76:16:@146436.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@146435.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@146439.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@146433.4]
  assign regs_144_clock = clock; // @[:@146442.4]
  assign regs_144_reset = io_reset; // @[:@146443.4 RegFile.scala 76:16:@146450.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@146449.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@146453.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@146447.4]
  assign regs_145_clock = clock; // @[:@146456.4]
  assign regs_145_reset = io_reset; // @[:@146457.4 RegFile.scala 76:16:@146464.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@146463.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@146467.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@146461.4]
  assign regs_146_clock = clock; // @[:@146470.4]
  assign regs_146_reset = io_reset; // @[:@146471.4 RegFile.scala 76:16:@146478.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@146477.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@146481.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@146475.4]
  assign regs_147_clock = clock; // @[:@146484.4]
  assign regs_147_reset = io_reset; // @[:@146485.4 RegFile.scala 76:16:@146492.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@146491.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@146495.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@146489.4]
  assign regs_148_clock = clock; // @[:@146498.4]
  assign regs_148_reset = io_reset; // @[:@146499.4 RegFile.scala 76:16:@146506.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@146505.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@146509.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@146503.4]
  assign regs_149_clock = clock; // @[:@146512.4]
  assign regs_149_reset = io_reset; // @[:@146513.4 RegFile.scala 76:16:@146520.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@146519.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@146523.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@146517.4]
  assign regs_150_clock = clock; // @[:@146526.4]
  assign regs_150_reset = io_reset; // @[:@146527.4 RegFile.scala 76:16:@146534.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@146533.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@146537.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@146531.4]
  assign regs_151_clock = clock; // @[:@146540.4]
  assign regs_151_reset = io_reset; // @[:@146541.4 RegFile.scala 76:16:@146548.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@146547.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@146551.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@146545.4]
  assign regs_152_clock = clock; // @[:@146554.4]
  assign regs_152_reset = io_reset; // @[:@146555.4 RegFile.scala 76:16:@146562.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@146561.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@146565.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@146559.4]
  assign regs_153_clock = clock; // @[:@146568.4]
  assign regs_153_reset = io_reset; // @[:@146569.4 RegFile.scala 76:16:@146576.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@146575.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@146579.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@146573.4]
  assign regs_154_clock = clock; // @[:@146582.4]
  assign regs_154_reset = io_reset; // @[:@146583.4 RegFile.scala 76:16:@146590.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@146589.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@146593.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@146587.4]
  assign regs_155_clock = clock; // @[:@146596.4]
  assign regs_155_reset = io_reset; // @[:@146597.4 RegFile.scala 76:16:@146604.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@146603.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@146607.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@146601.4]
  assign regs_156_clock = clock; // @[:@146610.4]
  assign regs_156_reset = io_reset; // @[:@146611.4 RegFile.scala 76:16:@146618.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@146617.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@146621.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@146615.4]
  assign regs_157_clock = clock; // @[:@146624.4]
  assign regs_157_reset = io_reset; // @[:@146625.4 RegFile.scala 76:16:@146632.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@146631.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@146635.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@146629.4]
  assign regs_158_clock = clock; // @[:@146638.4]
  assign regs_158_reset = io_reset; // @[:@146639.4 RegFile.scala 76:16:@146646.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@146645.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@146649.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@146643.4]
  assign regs_159_clock = clock; // @[:@146652.4]
  assign regs_159_reset = io_reset; // @[:@146653.4 RegFile.scala 76:16:@146660.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@146659.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@146663.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@146657.4]
  assign regs_160_clock = clock; // @[:@146666.4]
  assign regs_160_reset = io_reset; // @[:@146667.4 RegFile.scala 76:16:@146674.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@146673.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@146677.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@146671.4]
  assign regs_161_clock = clock; // @[:@146680.4]
  assign regs_161_reset = io_reset; // @[:@146681.4 RegFile.scala 76:16:@146688.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@146687.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@146691.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@146685.4]
  assign regs_162_clock = clock; // @[:@146694.4]
  assign regs_162_reset = io_reset; // @[:@146695.4 RegFile.scala 76:16:@146702.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@146701.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@146705.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@146699.4]
  assign regs_163_clock = clock; // @[:@146708.4]
  assign regs_163_reset = io_reset; // @[:@146709.4 RegFile.scala 76:16:@146716.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@146715.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@146719.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@146713.4]
  assign regs_164_clock = clock; // @[:@146722.4]
  assign regs_164_reset = io_reset; // @[:@146723.4 RegFile.scala 76:16:@146730.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@146729.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@146733.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@146727.4]
  assign regs_165_clock = clock; // @[:@146736.4]
  assign regs_165_reset = io_reset; // @[:@146737.4 RegFile.scala 76:16:@146744.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@146743.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@146747.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@146741.4]
  assign regs_166_clock = clock; // @[:@146750.4]
  assign regs_166_reset = io_reset; // @[:@146751.4 RegFile.scala 76:16:@146758.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@146757.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@146761.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@146755.4]
  assign regs_167_clock = clock; // @[:@146764.4]
  assign regs_167_reset = io_reset; // @[:@146765.4 RegFile.scala 76:16:@146772.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@146771.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@146775.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@146769.4]
  assign regs_168_clock = clock; // @[:@146778.4]
  assign regs_168_reset = io_reset; // @[:@146779.4 RegFile.scala 76:16:@146786.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@146785.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@146789.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@146783.4]
  assign regs_169_clock = clock; // @[:@146792.4]
  assign regs_169_reset = io_reset; // @[:@146793.4 RegFile.scala 76:16:@146800.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@146799.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@146803.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@146797.4]
  assign regs_170_clock = clock; // @[:@146806.4]
  assign regs_170_reset = io_reset; // @[:@146807.4 RegFile.scala 76:16:@146814.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@146813.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@146817.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@146811.4]
  assign regs_171_clock = clock; // @[:@146820.4]
  assign regs_171_reset = io_reset; // @[:@146821.4 RegFile.scala 76:16:@146828.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@146827.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@146831.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@146825.4]
  assign regs_172_clock = clock; // @[:@146834.4]
  assign regs_172_reset = io_reset; // @[:@146835.4 RegFile.scala 76:16:@146842.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@146841.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@146845.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@146839.4]
  assign regs_173_clock = clock; // @[:@146848.4]
  assign regs_173_reset = io_reset; // @[:@146849.4 RegFile.scala 76:16:@146856.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@146855.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@146859.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@146853.4]
  assign regs_174_clock = clock; // @[:@146862.4]
  assign regs_174_reset = io_reset; // @[:@146863.4 RegFile.scala 76:16:@146870.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@146869.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@146873.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@146867.4]
  assign regs_175_clock = clock; // @[:@146876.4]
  assign regs_175_reset = io_reset; // @[:@146877.4 RegFile.scala 76:16:@146884.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@146883.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@146887.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@146881.4]
  assign regs_176_clock = clock; // @[:@146890.4]
  assign regs_176_reset = io_reset; // @[:@146891.4 RegFile.scala 76:16:@146898.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@146897.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@146901.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@146895.4]
  assign regs_177_clock = clock; // @[:@146904.4]
  assign regs_177_reset = io_reset; // @[:@146905.4 RegFile.scala 76:16:@146912.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@146911.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@146915.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@146909.4]
  assign regs_178_clock = clock; // @[:@146918.4]
  assign regs_178_reset = io_reset; // @[:@146919.4 RegFile.scala 76:16:@146926.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@146925.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@146929.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@146923.4]
  assign regs_179_clock = clock; // @[:@146932.4]
  assign regs_179_reset = io_reset; // @[:@146933.4 RegFile.scala 76:16:@146940.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@146939.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@146943.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@146937.4]
  assign regs_180_clock = clock; // @[:@146946.4]
  assign regs_180_reset = io_reset; // @[:@146947.4 RegFile.scala 76:16:@146954.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@146953.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@146957.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@146951.4]
  assign regs_181_clock = clock; // @[:@146960.4]
  assign regs_181_reset = io_reset; // @[:@146961.4 RegFile.scala 76:16:@146968.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@146967.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@146971.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@146965.4]
  assign regs_182_clock = clock; // @[:@146974.4]
  assign regs_182_reset = io_reset; // @[:@146975.4 RegFile.scala 76:16:@146982.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@146981.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@146985.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@146979.4]
  assign regs_183_clock = clock; // @[:@146988.4]
  assign regs_183_reset = io_reset; // @[:@146989.4 RegFile.scala 76:16:@146996.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@146995.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@146999.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@146993.4]
  assign regs_184_clock = clock; // @[:@147002.4]
  assign regs_184_reset = io_reset; // @[:@147003.4 RegFile.scala 76:16:@147010.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@147009.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@147013.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@147007.4]
  assign regs_185_clock = clock; // @[:@147016.4]
  assign regs_185_reset = io_reset; // @[:@147017.4 RegFile.scala 76:16:@147024.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@147023.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@147027.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@147021.4]
  assign regs_186_clock = clock; // @[:@147030.4]
  assign regs_186_reset = io_reset; // @[:@147031.4 RegFile.scala 76:16:@147038.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@147037.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@147041.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@147035.4]
  assign regs_187_clock = clock; // @[:@147044.4]
  assign regs_187_reset = io_reset; // @[:@147045.4 RegFile.scala 76:16:@147052.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@147051.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@147055.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@147049.4]
  assign regs_188_clock = clock; // @[:@147058.4]
  assign regs_188_reset = io_reset; // @[:@147059.4 RegFile.scala 76:16:@147066.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@147065.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@147069.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@147063.4]
  assign regs_189_clock = clock; // @[:@147072.4]
  assign regs_189_reset = io_reset; // @[:@147073.4 RegFile.scala 76:16:@147080.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@147079.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@147083.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@147077.4]
  assign regs_190_clock = clock; // @[:@147086.4]
  assign regs_190_reset = io_reset; // @[:@147087.4 RegFile.scala 76:16:@147094.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@147093.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@147097.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@147091.4]
  assign regs_191_clock = clock; // @[:@147100.4]
  assign regs_191_reset = io_reset; // @[:@147101.4 RegFile.scala 76:16:@147108.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@147107.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@147111.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@147105.4]
  assign regs_192_clock = clock; // @[:@147114.4]
  assign regs_192_reset = io_reset; // @[:@147115.4 RegFile.scala 76:16:@147122.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@147121.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@147125.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@147119.4]
  assign regs_193_clock = clock; // @[:@147128.4]
  assign regs_193_reset = io_reset; // @[:@147129.4 RegFile.scala 76:16:@147136.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@147135.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@147139.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@147133.4]
  assign regs_194_clock = clock; // @[:@147142.4]
  assign regs_194_reset = io_reset; // @[:@147143.4 RegFile.scala 76:16:@147150.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@147149.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@147153.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@147147.4]
  assign regs_195_clock = clock; // @[:@147156.4]
  assign regs_195_reset = io_reset; // @[:@147157.4 RegFile.scala 76:16:@147164.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@147163.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@147167.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@147161.4]
  assign regs_196_clock = clock; // @[:@147170.4]
  assign regs_196_reset = io_reset; // @[:@147171.4 RegFile.scala 76:16:@147178.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@147177.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@147181.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@147175.4]
  assign regs_197_clock = clock; // @[:@147184.4]
  assign regs_197_reset = io_reset; // @[:@147185.4 RegFile.scala 76:16:@147192.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@147191.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@147195.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@147189.4]
  assign regs_198_clock = clock; // @[:@147198.4]
  assign regs_198_reset = io_reset; // @[:@147199.4 RegFile.scala 76:16:@147206.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@147205.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@147209.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@147203.4]
  assign regs_199_clock = clock; // @[:@147212.4]
  assign regs_199_reset = io_reset; // @[:@147213.4 RegFile.scala 76:16:@147220.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@147219.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@147223.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@147217.4]
  assign regs_200_clock = clock; // @[:@147226.4]
  assign regs_200_reset = io_reset; // @[:@147227.4 RegFile.scala 76:16:@147234.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@147233.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@147237.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@147231.4]
  assign regs_201_clock = clock; // @[:@147240.4]
  assign regs_201_reset = io_reset; // @[:@147241.4 RegFile.scala 76:16:@147248.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@147247.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@147251.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@147245.4]
  assign regs_202_clock = clock; // @[:@147254.4]
  assign regs_202_reset = io_reset; // @[:@147255.4 RegFile.scala 76:16:@147262.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@147261.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@147265.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@147259.4]
  assign regs_203_clock = clock; // @[:@147268.4]
  assign regs_203_reset = io_reset; // @[:@147269.4 RegFile.scala 76:16:@147276.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@147275.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@147279.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@147273.4]
  assign regs_204_clock = clock; // @[:@147282.4]
  assign regs_204_reset = io_reset; // @[:@147283.4 RegFile.scala 76:16:@147290.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@147289.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@147293.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@147287.4]
  assign regs_205_clock = clock; // @[:@147296.4]
  assign regs_205_reset = io_reset; // @[:@147297.4 RegFile.scala 76:16:@147304.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@147303.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@147307.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@147301.4]
  assign regs_206_clock = clock; // @[:@147310.4]
  assign regs_206_reset = io_reset; // @[:@147311.4 RegFile.scala 76:16:@147318.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@147317.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@147321.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@147315.4]
  assign regs_207_clock = clock; // @[:@147324.4]
  assign regs_207_reset = io_reset; // @[:@147325.4 RegFile.scala 76:16:@147332.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@147331.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@147335.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@147329.4]
  assign regs_208_clock = clock; // @[:@147338.4]
  assign regs_208_reset = io_reset; // @[:@147339.4 RegFile.scala 76:16:@147346.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@147345.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@147349.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@147343.4]
  assign regs_209_clock = clock; // @[:@147352.4]
  assign regs_209_reset = io_reset; // @[:@147353.4 RegFile.scala 76:16:@147360.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@147359.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@147363.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@147357.4]
  assign regs_210_clock = clock; // @[:@147366.4]
  assign regs_210_reset = io_reset; // @[:@147367.4 RegFile.scala 76:16:@147374.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@147373.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@147377.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@147371.4]
  assign regs_211_clock = clock; // @[:@147380.4]
  assign regs_211_reset = io_reset; // @[:@147381.4 RegFile.scala 76:16:@147388.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@147387.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@147391.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@147385.4]
  assign regs_212_clock = clock; // @[:@147394.4]
  assign regs_212_reset = io_reset; // @[:@147395.4 RegFile.scala 76:16:@147402.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@147401.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@147405.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@147399.4]
  assign regs_213_clock = clock; // @[:@147408.4]
  assign regs_213_reset = io_reset; // @[:@147409.4 RegFile.scala 76:16:@147416.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@147415.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@147419.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@147413.4]
  assign regs_214_clock = clock; // @[:@147422.4]
  assign regs_214_reset = io_reset; // @[:@147423.4 RegFile.scala 76:16:@147430.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@147429.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@147433.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@147427.4]
  assign regs_215_clock = clock; // @[:@147436.4]
  assign regs_215_reset = io_reset; // @[:@147437.4 RegFile.scala 76:16:@147444.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@147443.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@147447.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@147441.4]
  assign regs_216_clock = clock; // @[:@147450.4]
  assign regs_216_reset = io_reset; // @[:@147451.4 RegFile.scala 76:16:@147458.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@147457.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@147461.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@147455.4]
  assign regs_217_clock = clock; // @[:@147464.4]
  assign regs_217_reset = io_reset; // @[:@147465.4 RegFile.scala 76:16:@147472.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@147471.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@147475.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@147469.4]
  assign regs_218_clock = clock; // @[:@147478.4]
  assign regs_218_reset = io_reset; // @[:@147479.4 RegFile.scala 76:16:@147486.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@147485.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@147489.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@147483.4]
  assign regs_219_clock = clock; // @[:@147492.4]
  assign regs_219_reset = io_reset; // @[:@147493.4 RegFile.scala 76:16:@147500.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@147499.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@147503.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@147497.4]
  assign regs_220_clock = clock; // @[:@147506.4]
  assign regs_220_reset = io_reset; // @[:@147507.4 RegFile.scala 76:16:@147514.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@147513.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@147517.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@147511.4]
  assign regs_221_clock = clock; // @[:@147520.4]
  assign regs_221_reset = io_reset; // @[:@147521.4 RegFile.scala 76:16:@147528.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@147527.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@147531.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@147525.4]
  assign regs_222_clock = clock; // @[:@147534.4]
  assign regs_222_reset = io_reset; // @[:@147535.4 RegFile.scala 76:16:@147542.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@147541.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@147545.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@147539.4]
  assign regs_223_clock = clock; // @[:@147548.4]
  assign regs_223_reset = io_reset; // @[:@147549.4 RegFile.scala 76:16:@147556.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@147555.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@147559.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@147553.4]
  assign regs_224_clock = clock; // @[:@147562.4]
  assign regs_224_reset = io_reset; // @[:@147563.4 RegFile.scala 76:16:@147570.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@147569.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@147573.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@147567.4]
  assign regs_225_clock = clock; // @[:@147576.4]
  assign regs_225_reset = io_reset; // @[:@147577.4 RegFile.scala 76:16:@147584.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@147583.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@147587.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@147581.4]
  assign regs_226_clock = clock; // @[:@147590.4]
  assign regs_226_reset = io_reset; // @[:@147591.4 RegFile.scala 76:16:@147598.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@147597.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@147601.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@147595.4]
  assign regs_227_clock = clock; // @[:@147604.4]
  assign regs_227_reset = io_reset; // @[:@147605.4 RegFile.scala 76:16:@147612.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@147611.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@147615.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@147609.4]
  assign regs_228_clock = clock; // @[:@147618.4]
  assign regs_228_reset = io_reset; // @[:@147619.4 RegFile.scala 76:16:@147626.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@147625.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@147629.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@147623.4]
  assign regs_229_clock = clock; // @[:@147632.4]
  assign regs_229_reset = io_reset; // @[:@147633.4 RegFile.scala 76:16:@147640.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@147639.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@147643.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@147637.4]
  assign regs_230_clock = clock; // @[:@147646.4]
  assign regs_230_reset = io_reset; // @[:@147647.4 RegFile.scala 76:16:@147654.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@147653.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@147657.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@147651.4]
  assign regs_231_clock = clock; // @[:@147660.4]
  assign regs_231_reset = io_reset; // @[:@147661.4 RegFile.scala 76:16:@147668.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@147667.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@147671.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@147665.4]
  assign regs_232_clock = clock; // @[:@147674.4]
  assign regs_232_reset = io_reset; // @[:@147675.4 RegFile.scala 76:16:@147682.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@147681.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@147685.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@147679.4]
  assign regs_233_clock = clock; // @[:@147688.4]
  assign regs_233_reset = io_reset; // @[:@147689.4 RegFile.scala 76:16:@147696.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@147695.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@147699.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@147693.4]
  assign regs_234_clock = clock; // @[:@147702.4]
  assign regs_234_reset = io_reset; // @[:@147703.4 RegFile.scala 76:16:@147710.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@147709.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@147713.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@147707.4]
  assign regs_235_clock = clock; // @[:@147716.4]
  assign regs_235_reset = io_reset; // @[:@147717.4 RegFile.scala 76:16:@147724.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@147723.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@147727.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@147721.4]
  assign regs_236_clock = clock; // @[:@147730.4]
  assign regs_236_reset = io_reset; // @[:@147731.4 RegFile.scala 76:16:@147738.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@147737.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@147741.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@147735.4]
  assign regs_237_clock = clock; // @[:@147744.4]
  assign regs_237_reset = io_reset; // @[:@147745.4 RegFile.scala 76:16:@147752.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@147751.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@147755.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@147749.4]
  assign regs_238_clock = clock; // @[:@147758.4]
  assign regs_238_reset = io_reset; // @[:@147759.4 RegFile.scala 76:16:@147766.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@147765.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@147769.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@147763.4]
  assign regs_239_clock = clock; // @[:@147772.4]
  assign regs_239_reset = io_reset; // @[:@147773.4 RegFile.scala 76:16:@147780.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@147779.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@147783.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@147777.4]
  assign regs_240_clock = clock; // @[:@147786.4]
  assign regs_240_reset = io_reset; // @[:@147787.4 RegFile.scala 76:16:@147794.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@147793.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@147797.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@147791.4]
  assign regs_241_clock = clock; // @[:@147800.4]
  assign regs_241_reset = io_reset; // @[:@147801.4 RegFile.scala 76:16:@147808.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@147807.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@147811.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@147805.4]
  assign regs_242_clock = clock; // @[:@147814.4]
  assign regs_242_reset = io_reset; // @[:@147815.4 RegFile.scala 76:16:@147822.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@147821.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@147825.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@147819.4]
  assign regs_243_clock = clock; // @[:@147828.4]
  assign regs_243_reset = io_reset; // @[:@147829.4 RegFile.scala 76:16:@147836.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@147835.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@147839.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@147833.4]
  assign regs_244_clock = clock; // @[:@147842.4]
  assign regs_244_reset = io_reset; // @[:@147843.4 RegFile.scala 76:16:@147850.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@147849.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@147853.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@147847.4]
  assign regs_245_clock = clock; // @[:@147856.4]
  assign regs_245_reset = io_reset; // @[:@147857.4 RegFile.scala 76:16:@147864.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@147863.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@147867.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@147861.4]
  assign regs_246_clock = clock; // @[:@147870.4]
  assign regs_246_reset = io_reset; // @[:@147871.4 RegFile.scala 76:16:@147878.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@147877.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@147881.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@147875.4]
  assign regs_247_clock = clock; // @[:@147884.4]
  assign regs_247_reset = io_reset; // @[:@147885.4 RegFile.scala 76:16:@147892.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@147891.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@147895.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@147889.4]
  assign regs_248_clock = clock; // @[:@147898.4]
  assign regs_248_reset = io_reset; // @[:@147899.4 RegFile.scala 76:16:@147906.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@147905.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@147909.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@147903.4]
  assign regs_249_clock = clock; // @[:@147912.4]
  assign regs_249_reset = io_reset; // @[:@147913.4 RegFile.scala 76:16:@147920.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@147919.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@147923.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@147917.4]
  assign regs_250_clock = clock; // @[:@147926.4]
  assign regs_250_reset = io_reset; // @[:@147927.4 RegFile.scala 76:16:@147934.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@147933.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@147937.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@147931.4]
  assign regs_251_clock = clock; // @[:@147940.4]
  assign regs_251_reset = io_reset; // @[:@147941.4 RegFile.scala 76:16:@147948.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@147947.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@147951.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@147945.4]
  assign regs_252_clock = clock; // @[:@147954.4]
  assign regs_252_reset = io_reset; // @[:@147955.4 RegFile.scala 76:16:@147962.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@147961.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@147965.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@147959.4]
  assign regs_253_clock = clock; // @[:@147968.4]
  assign regs_253_reset = io_reset; // @[:@147969.4 RegFile.scala 76:16:@147976.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@147975.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@147979.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@147973.4]
  assign regs_254_clock = clock; // @[:@147982.4]
  assign regs_254_reset = io_reset; // @[:@147983.4 RegFile.scala 76:16:@147990.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@147989.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@147993.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@147987.4]
  assign regs_255_clock = clock; // @[:@147996.4]
  assign regs_255_reset = io_reset; // @[:@147997.4 RegFile.scala 76:16:@148004.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@148003.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@148007.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@148001.4]
  assign regs_256_clock = clock; // @[:@148010.4]
  assign regs_256_reset = io_reset; // @[:@148011.4 RegFile.scala 76:16:@148018.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@148017.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@148021.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@148015.4]
  assign regs_257_clock = clock; // @[:@148024.4]
  assign regs_257_reset = io_reset; // @[:@148025.4 RegFile.scala 76:16:@148032.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@148031.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@148035.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@148029.4]
  assign regs_258_clock = clock; // @[:@148038.4]
  assign regs_258_reset = io_reset; // @[:@148039.4 RegFile.scala 76:16:@148046.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@148045.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@148049.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@148043.4]
  assign regs_259_clock = clock; // @[:@148052.4]
  assign regs_259_reset = io_reset; // @[:@148053.4 RegFile.scala 76:16:@148060.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@148059.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@148063.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@148057.4]
  assign regs_260_clock = clock; // @[:@148066.4]
  assign regs_260_reset = io_reset; // @[:@148067.4 RegFile.scala 76:16:@148074.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@148073.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@148077.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@148071.4]
  assign regs_261_clock = clock; // @[:@148080.4]
  assign regs_261_reset = io_reset; // @[:@148081.4 RegFile.scala 76:16:@148088.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@148087.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@148091.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@148085.4]
  assign regs_262_clock = clock; // @[:@148094.4]
  assign regs_262_reset = io_reset; // @[:@148095.4 RegFile.scala 76:16:@148102.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@148101.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@148105.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@148099.4]
  assign regs_263_clock = clock; // @[:@148108.4]
  assign regs_263_reset = io_reset; // @[:@148109.4 RegFile.scala 76:16:@148116.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@148115.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@148119.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@148113.4]
  assign regs_264_clock = clock; // @[:@148122.4]
  assign regs_264_reset = io_reset; // @[:@148123.4 RegFile.scala 76:16:@148130.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@148129.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@148133.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@148127.4]
  assign regs_265_clock = clock; // @[:@148136.4]
  assign regs_265_reset = io_reset; // @[:@148137.4 RegFile.scala 76:16:@148144.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@148143.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@148147.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@148141.4]
  assign regs_266_clock = clock; // @[:@148150.4]
  assign regs_266_reset = io_reset; // @[:@148151.4 RegFile.scala 76:16:@148158.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@148157.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@148161.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@148155.4]
  assign regs_267_clock = clock; // @[:@148164.4]
  assign regs_267_reset = io_reset; // @[:@148165.4 RegFile.scala 76:16:@148172.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@148171.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@148175.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@148169.4]
  assign regs_268_clock = clock; // @[:@148178.4]
  assign regs_268_reset = io_reset; // @[:@148179.4 RegFile.scala 76:16:@148186.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@148185.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@148189.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@148183.4]
  assign regs_269_clock = clock; // @[:@148192.4]
  assign regs_269_reset = io_reset; // @[:@148193.4 RegFile.scala 76:16:@148200.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@148199.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@148203.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@148197.4]
  assign regs_270_clock = clock; // @[:@148206.4]
  assign regs_270_reset = io_reset; // @[:@148207.4 RegFile.scala 76:16:@148214.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@148213.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@148217.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@148211.4]
  assign regs_271_clock = clock; // @[:@148220.4]
  assign regs_271_reset = io_reset; // @[:@148221.4 RegFile.scala 76:16:@148228.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@148227.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@148231.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@148225.4]
  assign regs_272_clock = clock; // @[:@148234.4]
  assign regs_272_reset = io_reset; // @[:@148235.4 RegFile.scala 76:16:@148242.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@148241.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@148245.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@148239.4]
  assign regs_273_clock = clock; // @[:@148248.4]
  assign regs_273_reset = io_reset; // @[:@148249.4 RegFile.scala 76:16:@148256.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@148255.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@148259.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@148253.4]
  assign regs_274_clock = clock; // @[:@148262.4]
  assign regs_274_reset = io_reset; // @[:@148263.4 RegFile.scala 76:16:@148270.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@148269.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@148273.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@148267.4]
  assign regs_275_clock = clock; // @[:@148276.4]
  assign regs_275_reset = io_reset; // @[:@148277.4 RegFile.scala 76:16:@148284.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@148283.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@148287.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@148281.4]
  assign regs_276_clock = clock; // @[:@148290.4]
  assign regs_276_reset = io_reset; // @[:@148291.4 RegFile.scala 76:16:@148298.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@148297.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@148301.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@148295.4]
  assign regs_277_clock = clock; // @[:@148304.4]
  assign regs_277_reset = io_reset; // @[:@148305.4 RegFile.scala 76:16:@148312.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@148311.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@148315.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@148309.4]
  assign regs_278_clock = clock; // @[:@148318.4]
  assign regs_278_reset = io_reset; // @[:@148319.4 RegFile.scala 76:16:@148326.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@148325.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@148329.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@148323.4]
  assign regs_279_clock = clock; // @[:@148332.4]
  assign regs_279_reset = io_reset; // @[:@148333.4 RegFile.scala 76:16:@148340.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@148339.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@148343.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@148337.4]
  assign regs_280_clock = clock; // @[:@148346.4]
  assign regs_280_reset = io_reset; // @[:@148347.4 RegFile.scala 76:16:@148354.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@148353.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@148357.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@148351.4]
  assign regs_281_clock = clock; // @[:@148360.4]
  assign regs_281_reset = io_reset; // @[:@148361.4 RegFile.scala 76:16:@148368.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@148367.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@148371.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@148365.4]
  assign regs_282_clock = clock; // @[:@148374.4]
  assign regs_282_reset = io_reset; // @[:@148375.4 RegFile.scala 76:16:@148382.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@148381.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@148385.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@148379.4]
  assign regs_283_clock = clock; // @[:@148388.4]
  assign regs_283_reset = io_reset; // @[:@148389.4 RegFile.scala 76:16:@148396.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@148395.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@148399.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@148393.4]
  assign regs_284_clock = clock; // @[:@148402.4]
  assign regs_284_reset = io_reset; // @[:@148403.4 RegFile.scala 76:16:@148410.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@148409.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@148413.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@148407.4]
  assign regs_285_clock = clock; // @[:@148416.4]
  assign regs_285_reset = io_reset; // @[:@148417.4 RegFile.scala 76:16:@148424.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@148423.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@148427.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@148421.4]
  assign regs_286_clock = clock; // @[:@148430.4]
  assign regs_286_reset = io_reset; // @[:@148431.4 RegFile.scala 76:16:@148438.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@148437.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@148441.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@148435.4]
  assign regs_287_clock = clock; // @[:@148444.4]
  assign regs_287_reset = io_reset; // @[:@148445.4 RegFile.scala 76:16:@148452.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@148451.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@148455.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@148449.4]
  assign regs_288_clock = clock; // @[:@148458.4]
  assign regs_288_reset = io_reset; // @[:@148459.4 RegFile.scala 76:16:@148466.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@148465.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@148469.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@148463.4]
  assign regs_289_clock = clock; // @[:@148472.4]
  assign regs_289_reset = io_reset; // @[:@148473.4 RegFile.scala 76:16:@148480.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@148479.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@148483.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@148477.4]
  assign regs_290_clock = clock; // @[:@148486.4]
  assign regs_290_reset = io_reset; // @[:@148487.4 RegFile.scala 76:16:@148494.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@148493.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@148497.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@148491.4]
  assign regs_291_clock = clock; // @[:@148500.4]
  assign regs_291_reset = io_reset; // @[:@148501.4 RegFile.scala 76:16:@148508.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@148507.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@148511.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@148505.4]
  assign regs_292_clock = clock; // @[:@148514.4]
  assign regs_292_reset = io_reset; // @[:@148515.4 RegFile.scala 76:16:@148522.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@148521.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@148525.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@148519.4]
  assign regs_293_clock = clock; // @[:@148528.4]
  assign regs_293_reset = io_reset; // @[:@148529.4 RegFile.scala 76:16:@148536.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@148535.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@148539.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@148533.4]
  assign regs_294_clock = clock; // @[:@148542.4]
  assign regs_294_reset = io_reset; // @[:@148543.4 RegFile.scala 76:16:@148550.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@148549.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@148553.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@148547.4]
  assign regs_295_clock = clock; // @[:@148556.4]
  assign regs_295_reset = io_reset; // @[:@148557.4 RegFile.scala 76:16:@148564.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@148563.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@148567.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@148561.4]
  assign regs_296_clock = clock; // @[:@148570.4]
  assign regs_296_reset = io_reset; // @[:@148571.4 RegFile.scala 76:16:@148578.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@148577.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@148581.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@148575.4]
  assign regs_297_clock = clock; // @[:@148584.4]
  assign regs_297_reset = io_reset; // @[:@148585.4 RegFile.scala 76:16:@148592.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@148591.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@148595.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@148589.4]
  assign regs_298_clock = clock; // @[:@148598.4]
  assign regs_298_reset = io_reset; // @[:@148599.4 RegFile.scala 76:16:@148606.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@148605.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@148609.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@148603.4]
  assign regs_299_clock = clock; // @[:@148612.4]
  assign regs_299_reset = io_reset; // @[:@148613.4 RegFile.scala 76:16:@148620.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@148619.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@148623.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@148617.4]
  assign regs_300_clock = clock; // @[:@148626.4]
  assign regs_300_reset = io_reset; // @[:@148627.4 RegFile.scala 76:16:@148634.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@148633.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@148637.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@148631.4]
  assign regs_301_clock = clock; // @[:@148640.4]
  assign regs_301_reset = io_reset; // @[:@148641.4 RegFile.scala 76:16:@148648.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@148647.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@148651.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@148645.4]
  assign regs_302_clock = clock; // @[:@148654.4]
  assign regs_302_reset = io_reset; // @[:@148655.4 RegFile.scala 76:16:@148662.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@148661.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@148665.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@148659.4]
  assign regs_303_clock = clock; // @[:@148668.4]
  assign regs_303_reset = io_reset; // @[:@148669.4 RegFile.scala 76:16:@148676.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@148675.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@148679.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@148673.4]
  assign regs_304_clock = clock; // @[:@148682.4]
  assign regs_304_reset = io_reset; // @[:@148683.4 RegFile.scala 76:16:@148690.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@148689.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@148693.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@148687.4]
  assign regs_305_clock = clock; // @[:@148696.4]
  assign regs_305_reset = io_reset; // @[:@148697.4 RegFile.scala 76:16:@148704.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@148703.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@148707.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@148701.4]
  assign regs_306_clock = clock; // @[:@148710.4]
  assign regs_306_reset = io_reset; // @[:@148711.4 RegFile.scala 76:16:@148718.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@148717.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@148721.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@148715.4]
  assign regs_307_clock = clock; // @[:@148724.4]
  assign regs_307_reset = io_reset; // @[:@148725.4 RegFile.scala 76:16:@148732.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@148731.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@148735.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@148729.4]
  assign regs_308_clock = clock; // @[:@148738.4]
  assign regs_308_reset = io_reset; // @[:@148739.4 RegFile.scala 76:16:@148746.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@148745.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@148749.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@148743.4]
  assign regs_309_clock = clock; // @[:@148752.4]
  assign regs_309_reset = io_reset; // @[:@148753.4 RegFile.scala 76:16:@148760.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@148759.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@148763.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@148757.4]
  assign regs_310_clock = clock; // @[:@148766.4]
  assign regs_310_reset = io_reset; // @[:@148767.4 RegFile.scala 76:16:@148774.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@148773.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@148777.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@148771.4]
  assign regs_311_clock = clock; // @[:@148780.4]
  assign regs_311_reset = io_reset; // @[:@148781.4 RegFile.scala 76:16:@148788.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@148787.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@148791.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@148785.4]
  assign regs_312_clock = clock; // @[:@148794.4]
  assign regs_312_reset = io_reset; // @[:@148795.4 RegFile.scala 76:16:@148802.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@148801.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@148805.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@148799.4]
  assign regs_313_clock = clock; // @[:@148808.4]
  assign regs_313_reset = io_reset; // @[:@148809.4 RegFile.scala 76:16:@148816.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@148815.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@148819.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@148813.4]
  assign regs_314_clock = clock; // @[:@148822.4]
  assign regs_314_reset = io_reset; // @[:@148823.4 RegFile.scala 76:16:@148830.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@148829.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@148833.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@148827.4]
  assign regs_315_clock = clock; // @[:@148836.4]
  assign regs_315_reset = io_reset; // @[:@148837.4 RegFile.scala 76:16:@148844.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@148843.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@148847.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@148841.4]
  assign regs_316_clock = clock; // @[:@148850.4]
  assign regs_316_reset = io_reset; // @[:@148851.4 RegFile.scala 76:16:@148858.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@148857.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@148861.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@148855.4]
  assign regs_317_clock = clock; // @[:@148864.4]
  assign regs_317_reset = io_reset; // @[:@148865.4 RegFile.scala 76:16:@148872.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@148871.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@148875.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@148869.4]
  assign regs_318_clock = clock; // @[:@148878.4]
  assign regs_318_reset = io_reset; // @[:@148879.4 RegFile.scala 76:16:@148886.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@148885.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@148889.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@148883.4]
  assign regs_319_clock = clock; // @[:@148892.4]
  assign regs_319_reset = io_reset; // @[:@148893.4 RegFile.scala 76:16:@148900.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@148899.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@148903.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@148897.4]
  assign regs_320_clock = clock; // @[:@148906.4]
  assign regs_320_reset = io_reset; // @[:@148907.4 RegFile.scala 76:16:@148914.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@148913.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@148917.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@148911.4]
  assign regs_321_clock = clock; // @[:@148920.4]
  assign regs_321_reset = io_reset; // @[:@148921.4 RegFile.scala 76:16:@148928.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@148927.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@148931.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@148925.4]
  assign regs_322_clock = clock; // @[:@148934.4]
  assign regs_322_reset = io_reset; // @[:@148935.4 RegFile.scala 76:16:@148942.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@148941.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@148945.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@148939.4]
  assign regs_323_clock = clock; // @[:@148948.4]
  assign regs_323_reset = io_reset; // @[:@148949.4 RegFile.scala 76:16:@148956.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@148955.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@148959.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@148953.4]
  assign regs_324_clock = clock; // @[:@148962.4]
  assign regs_324_reset = io_reset; // @[:@148963.4 RegFile.scala 76:16:@148970.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@148969.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@148973.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@148967.4]
  assign regs_325_clock = clock; // @[:@148976.4]
  assign regs_325_reset = io_reset; // @[:@148977.4 RegFile.scala 76:16:@148984.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@148983.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@148987.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@148981.4]
  assign regs_326_clock = clock; // @[:@148990.4]
  assign regs_326_reset = io_reset; // @[:@148991.4 RegFile.scala 76:16:@148998.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@148997.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@149001.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@148995.4]
  assign regs_327_clock = clock; // @[:@149004.4]
  assign regs_327_reset = io_reset; // @[:@149005.4 RegFile.scala 76:16:@149012.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@149011.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@149015.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@149009.4]
  assign regs_328_clock = clock; // @[:@149018.4]
  assign regs_328_reset = io_reset; // @[:@149019.4 RegFile.scala 76:16:@149026.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@149025.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@149029.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@149023.4]
  assign regs_329_clock = clock; // @[:@149032.4]
  assign regs_329_reset = io_reset; // @[:@149033.4 RegFile.scala 76:16:@149040.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@149039.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@149043.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@149037.4]
  assign regs_330_clock = clock; // @[:@149046.4]
  assign regs_330_reset = io_reset; // @[:@149047.4 RegFile.scala 76:16:@149054.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@149053.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@149057.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@149051.4]
  assign regs_331_clock = clock; // @[:@149060.4]
  assign regs_331_reset = io_reset; // @[:@149061.4 RegFile.scala 76:16:@149068.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@149067.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@149071.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@149065.4]
  assign regs_332_clock = clock; // @[:@149074.4]
  assign regs_332_reset = io_reset; // @[:@149075.4 RegFile.scala 76:16:@149082.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@149081.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@149085.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@149079.4]
  assign regs_333_clock = clock; // @[:@149088.4]
  assign regs_333_reset = io_reset; // @[:@149089.4 RegFile.scala 76:16:@149096.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@149095.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@149099.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@149093.4]
  assign regs_334_clock = clock; // @[:@149102.4]
  assign regs_334_reset = io_reset; // @[:@149103.4 RegFile.scala 76:16:@149110.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@149109.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@149113.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@149107.4]
  assign regs_335_clock = clock; // @[:@149116.4]
  assign regs_335_reset = io_reset; // @[:@149117.4 RegFile.scala 76:16:@149124.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@149123.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@149127.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@149121.4]
  assign regs_336_clock = clock; // @[:@149130.4]
  assign regs_336_reset = io_reset; // @[:@149131.4 RegFile.scala 76:16:@149138.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@149137.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@149141.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@149135.4]
  assign regs_337_clock = clock; // @[:@149144.4]
  assign regs_337_reset = io_reset; // @[:@149145.4 RegFile.scala 76:16:@149152.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@149151.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@149155.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@149149.4]
  assign regs_338_clock = clock; // @[:@149158.4]
  assign regs_338_reset = io_reset; // @[:@149159.4 RegFile.scala 76:16:@149166.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@149165.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@149169.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@149163.4]
  assign regs_339_clock = clock; // @[:@149172.4]
  assign regs_339_reset = io_reset; // @[:@149173.4 RegFile.scala 76:16:@149180.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@149179.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@149183.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@149177.4]
  assign regs_340_clock = clock; // @[:@149186.4]
  assign regs_340_reset = io_reset; // @[:@149187.4 RegFile.scala 76:16:@149194.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@149193.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@149197.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@149191.4]
  assign regs_341_clock = clock; // @[:@149200.4]
  assign regs_341_reset = io_reset; // @[:@149201.4 RegFile.scala 76:16:@149208.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@149207.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@149211.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@149205.4]
  assign regs_342_clock = clock; // @[:@149214.4]
  assign regs_342_reset = io_reset; // @[:@149215.4 RegFile.scala 76:16:@149222.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@149221.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@149225.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@149219.4]
  assign regs_343_clock = clock; // @[:@149228.4]
  assign regs_343_reset = io_reset; // @[:@149229.4 RegFile.scala 76:16:@149236.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@149235.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@149239.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@149233.4]
  assign regs_344_clock = clock; // @[:@149242.4]
  assign regs_344_reset = io_reset; // @[:@149243.4 RegFile.scala 76:16:@149250.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@149249.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@149253.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@149247.4]
  assign regs_345_clock = clock; // @[:@149256.4]
  assign regs_345_reset = io_reset; // @[:@149257.4 RegFile.scala 76:16:@149264.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@149263.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@149267.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@149261.4]
  assign regs_346_clock = clock; // @[:@149270.4]
  assign regs_346_reset = io_reset; // @[:@149271.4 RegFile.scala 76:16:@149278.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@149277.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@149281.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@149275.4]
  assign regs_347_clock = clock; // @[:@149284.4]
  assign regs_347_reset = io_reset; // @[:@149285.4 RegFile.scala 76:16:@149292.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@149291.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@149295.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@149289.4]
  assign regs_348_clock = clock; // @[:@149298.4]
  assign regs_348_reset = io_reset; // @[:@149299.4 RegFile.scala 76:16:@149306.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@149305.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@149309.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@149303.4]
  assign regs_349_clock = clock; // @[:@149312.4]
  assign regs_349_reset = io_reset; // @[:@149313.4 RegFile.scala 76:16:@149320.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@149319.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@149323.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@149317.4]
  assign regs_350_clock = clock; // @[:@149326.4]
  assign regs_350_reset = io_reset; // @[:@149327.4 RegFile.scala 76:16:@149334.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@149333.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@149337.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@149331.4]
  assign regs_351_clock = clock; // @[:@149340.4]
  assign regs_351_reset = io_reset; // @[:@149341.4 RegFile.scala 76:16:@149348.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@149347.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@149351.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@149345.4]
  assign regs_352_clock = clock; // @[:@149354.4]
  assign regs_352_reset = io_reset; // @[:@149355.4 RegFile.scala 76:16:@149362.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@149361.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@149365.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@149359.4]
  assign regs_353_clock = clock; // @[:@149368.4]
  assign regs_353_reset = io_reset; // @[:@149369.4 RegFile.scala 76:16:@149376.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@149375.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@149379.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@149373.4]
  assign regs_354_clock = clock; // @[:@149382.4]
  assign regs_354_reset = io_reset; // @[:@149383.4 RegFile.scala 76:16:@149390.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@149389.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@149393.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@149387.4]
  assign regs_355_clock = clock; // @[:@149396.4]
  assign regs_355_reset = io_reset; // @[:@149397.4 RegFile.scala 76:16:@149404.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@149403.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@149407.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@149401.4]
  assign regs_356_clock = clock; // @[:@149410.4]
  assign regs_356_reset = io_reset; // @[:@149411.4 RegFile.scala 76:16:@149418.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@149417.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@149421.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@149415.4]
  assign regs_357_clock = clock; // @[:@149424.4]
  assign regs_357_reset = io_reset; // @[:@149425.4 RegFile.scala 76:16:@149432.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@149431.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@149435.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@149429.4]
  assign regs_358_clock = clock; // @[:@149438.4]
  assign regs_358_reset = io_reset; // @[:@149439.4 RegFile.scala 76:16:@149446.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@149445.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@149449.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@149443.4]
  assign regs_359_clock = clock; // @[:@149452.4]
  assign regs_359_reset = io_reset; // @[:@149453.4 RegFile.scala 76:16:@149460.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@149459.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@149463.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@149457.4]
  assign regs_360_clock = clock; // @[:@149466.4]
  assign regs_360_reset = io_reset; // @[:@149467.4 RegFile.scala 76:16:@149474.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@149473.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@149477.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@149471.4]
  assign regs_361_clock = clock; // @[:@149480.4]
  assign regs_361_reset = io_reset; // @[:@149481.4 RegFile.scala 76:16:@149488.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@149487.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@149491.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@149485.4]
  assign regs_362_clock = clock; // @[:@149494.4]
  assign regs_362_reset = io_reset; // @[:@149495.4 RegFile.scala 76:16:@149502.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@149501.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@149505.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@149499.4]
  assign regs_363_clock = clock; // @[:@149508.4]
  assign regs_363_reset = io_reset; // @[:@149509.4 RegFile.scala 76:16:@149516.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@149515.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@149519.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@149513.4]
  assign regs_364_clock = clock; // @[:@149522.4]
  assign regs_364_reset = io_reset; // @[:@149523.4 RegFile.scala 76:16:@149530.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@149529.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@149533.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@149527.4]
  assign regs_365_clock = clock; // @[:@149536.4]
  assign regs_365_reset = io_reset; // @[:@149537.4 RegFile.scala 76:16:@149544.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@149543.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@149547.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@149541.4]
  assign regs_366_clock = clock; // @[:@149550.4]
  assign regs_366_reset = io_reset; // @[:@149551.4 RegFile.scala 76:16:@149558.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@149557.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@149561.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@149555.4]
  assign regs_367_clock = clock; // @[:@149564.4]
  assign regs_367_reset = io_reset; // @[:@149565.4 RegFile.scala 76:16:@149572.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@149571.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@149575.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@149569.4]
  assign regs_368_clock = clock; // @[:@149578.4]
  assign regs_368_reset = io_reset; // @[:@149579.4 RegFile.scala 76:16:@149586.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@149585.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@149589.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@149583.4]
  assign regs_369_clock = clock; // @[:@149592.4]
  assign regs_369_reset = io_reset; // @[:@149593.4 RegFile.scala 76:16:@149600.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@149599.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@149603.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@149597.4]
  assign regs_370_clock = clock; // @[:@149606.4]
  assign regs_370_reset = io_reset; // @[:@149607.4 RegFile.scala 76:16:@149614.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@149613.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@149617.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@149611.4]
  assign regs_371_clock = clock; // @[:@149620.4]
  assign regs_371_reset = io_reset; // @[:@149621.4 RegFile.scala 76:16:@149628.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@149627.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@149631.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@149625.4]
  assign regs_372_clock = clock; // @[:@149634.4]
  assign regs_372_reset = io_reset; // @[:@149635.4 RegFile.scala 76:16:@149642.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@149641.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@149645.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@149639.4]
  assign regs_373_clock = clock; // @[:@149648.4]
  assign regs_373_reset = io_reset; // @[:@149649.4 RegFile.scala 76:16:@149656.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@149655.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@149659.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@149653.4]
  assign regs_374_clock = clock; // @[:@149662.4]
  assign regs_374_reset = io_reset; // @[:@149663.4 RegFile.scala 76:16:@149670.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@149669.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@149673.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@149667.4]
  assign regs_375_clock = clock; // @[:@149676.4]
  assign regs_375_reset = io_reset; // @[:@149677.4 RegFile.scala 76:16:@149684.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@149683.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@149687.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@149681.4]
  assign regs_376_clock = clock; // @[:@149690.4]
  assign regs_376_reset = io_reset; // @[:@149691.4 RegFile.scala 76:16:@149698.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@149697.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@149701.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@149695.4]
  assign regs_377_clock = clock; // @[:@149704.4]
  assign regs_377_reset = io_reset; // @[:@149705.4 RegFile.scala 76:16:@149712.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@149711.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@149715.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@149709.4]
  assign regs_378_clock = clock; // @[:@149718.4]
  assign regs_378_reset = io_reset; // @[:@149719.4 RegFile.scala 76:16:@149726.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@149725.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@149729.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@149723.4]
  assign regs_379_clock = clock; // @[:@149732.4]
  assign regs_379_reset = io_reset; // @[:@149733.4 RegFile.scala 76:16:@149740.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@149739.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@149743.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@149737.4]
  assign regs_380_clock = clock; // @[:@149746.4]
  assign regs_380_reset = io_reset; // @[:@149747.4 RegFile.scala 76:16:@149754.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@149753.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@149757.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@149751.4]
  assign regs_381_clock = clock; // @[:@149760.4]
  assign regs_381_reset = io_reset; // @[:@149761.4 RegFile.scala 76:16:@149768.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@149767.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@149771.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@149765.4]
  assign regs_382_clock = clock; // @[:@149774.4]
  assign regs_382_reset = io_reset; // @[:@149775.4 RegFile.scala 76:16:@149782.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@149781.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@149785.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@149779.4]
  assign regs_383_clock = clock; // @[:@149788.4]
  assign regs_383_reset = io_reset; // @[:@149789.4 RegFile.scala 76:16:@149796.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@149795.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@149799.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@149793.4]
  assign regs_384_clock = clock; // @[:@149802.4]
  assign regs_384_reset = io_reset; // @[:@149803.4 RegFile.scala 76:16:@149810.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@149809.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@149813.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@149807.4]
  assign regs_385_clock = clock; // @[:@149816.4]
  assign regs_385_reset = io_reset; // @[:@149817.4 RegFile.scala 76:16:@149824.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@149823.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@149827.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@149821.4]
  assign regs_386_clock = clock; // @[:@149830.4]
  assign regs_386_reset = io_reset; // @[:@149831.4 RegFile.scala 76:16:@149838.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@149837.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@149841.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@149835.4]
  assign regs_387_clock = clock; // @[:@149844.4]
  assign regs_387_reset = io_reset; // @[:@149845.4 RegFile.scala 76:16:@149852.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@149851.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@149855.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@149849.4]
  assign regs_388_clock = clock; // @[:@149858.4]
  assign regs_388_reset = io_reset; // @[:@149859.4 RegFile.scala 76:16:@149866.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@149865.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@149869.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@149863.4]
  assign regs_389_clock = clock; // @[:@149872.4]
  assign regs_389_reset = io_reset; // @[:@149873.4 RegFile.scala 76:16:@149880.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@149879.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@149883.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@149877.4]
  assign regs_390_clock = clock; // @[:@149886.4]
  assign regs_390_reset = io_reset; // @[:@149887.4 RegFile.scala 76:16:@149894.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@149893.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@149897.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@149891.4]
  assign regs_391_clock = clock; // @[:@149900.4]
  assign regs_391_reset = io_reset; // @[:@149901.4 RegFile.scala 76:16:@149908.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@149907.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@149911.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@149905.4]
  assign regs_392_clock = clock; // @[:@149914.4]
  assign regs_392_reset = io_reset; // @[:@149915.4 RegFile.scala 76:16:@149922.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@149921.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@149925.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@149919.4]
  assign regs_393_clock = clock; // @[:@149928.4]
  assign regs_393_reset = io_reset; // @[:@149929.4 RegFile.scala 76:16:@149936.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@149935.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@149939.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@149933.4]
  assign regs_394_clock = clock; // @[:@149942.4]
  assign regs_394_reset = io_reset; // @[:@149943.4 RegFile.scala 76:16:@149950.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@149949.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@149953.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@149947.4]
  assign regs_395_clock = clock; // @[:@149956.4]
  assign regs_395_reset = io_reset; // @[:@149957.4 RegFile.scala 76:16:@149964.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@149963.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@149967.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@149961.4]
  assign regs_396_clock = clock; // @[:@149970.4]
  assign regs_396_reset = io_reset; // @[:@149971.4 RegFile.scala 76:16:@149978.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@149977.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@149981.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@149975.4]
  assign regs_397_clock = clock; // @[:@149984.4]
  assign regs_397_reset = io_reset; // @[:@149985.4 RegFile.scala 76:16:@149992.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@149991.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@149995.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@149989.4]
  assign regs_398_clock = clock; // @[:@149998.4]
  assign regs_398_reset = io_reset; // @[:@149999.4 RegFile.scala 76:16:@150006.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@150005.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@150009.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@150003.4]
  assign regs_399_clock = clock; // @[:@150012.4]
  assign regs_399_reset = io_reset; // @[:@150013.4 RegFile.scala 76:16:@150020.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@150019.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@150023.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@150017.4]
  assign regs_400_clock = clock; // @[:@150026.4]
  assign regs_400_reset = io_reset; // @[:@150027.4 RegFile.scala 76:16:@150034.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@150033.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@150037.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@150031.4]
  assign regs_401_clock = clock; // @[:@150040.4]
  assign regs_401_reset = io_reset; // @[:@150041.4 RegFile.scala 76:16:@150048.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@150047.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@150051.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@150045.4]
  assign regs_402_clock = clock; // @[:@150054.4]
  assign regs_402_reset = io_reset; // @[:@150055.4 RegFile.scala 76:16:@150062.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@150061.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@150065.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@150059.4]
  assign regs_403_clock = clock; // @[:@150068.4]
  assign regs_403_reset = io_reset; // @[:@150069.4 RegFile.scala 76:16:@150076.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@150075.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@150079.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@150073.4]
  assign regs_404_clock = clock; // @[:@150082.4]
  assign regs_404_reset = io_reset; // @[:@150083.4 RegFile.scala 76:16:@150090.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@150089.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@150093.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@150087.4]
  assign regs_405_clock = clock; // @[:@150096.4]
  assign regs_405_reset = io_reset; // @[:@150097.4 RegFile.scala 76:16:@150104.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@150103.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@150107.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@150101.4]
  assign regs_406_clock = clock; // @[:@150110.4]
  assign regs_406_reset = io_reset; // @[:@150111.4 RegFile.scala 76:16:@150118.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@150117.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@150121.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@150115.4]
  assign regs_407_clock = clock; // @[:@150124.4]
  assign regs_407_reset = io_reset; // @[:@150125.4 RegFile.scala 76:16:@150132.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@150131.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@150135.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@150129.4]
  assign regs_408_clock = clock; // @[:@150138.4]
  assign regs_408_reset = io_reset; // @[:@150139.4 RegFile.scala 76:16:@150146.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@150145.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@150149.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@150143.4]
  assign regs_409_clock = clock; // @[:@150152.4]
  assign regs_409_reset = io_reset; // @[:@150153.4 RegFile.scala 76:16:@150160.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@150159.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@150163.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@150157.4]
  assign regs_410_clock = clock; // @[:@150166.4]
  assign regs_410_reset = io_reset; // @[:@150167.4 RegFile.scala 76:16:@150174.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@150173.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@150177.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@150171.4]
  assign regs_411_clock = clock; // @[:@150180.4]
  assign regs_411_reset = io_reset; // @[:@150181.4 RegFile.scala 76:16:@150188.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@150187.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@150191.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@150185.4]
  assign regs_412_clock = clock; // @[:@150194.4]
  assign regs_412_reset = io_reset; // @[:@150195.4 RegFile.scala 76:16:@150202.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@150201.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@150205.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@150199.4]
  assign regs_413_clock = clock; // @[:@150208.4]
  assign regs_413_reset = io_reset; // @[:@150209.4 RegFile.scala 76:16:@150216.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@150215.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@150219.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@150213.4]
  assign regs_414_clock = clock; // @[:@150222.4]
  assign regs_414_reset = io_reset; // @[:@150223.4 RegFile.scala 76:16:@150230.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@150229.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@150233.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@150227.4]
  assign regs_415_clock = clock; // @[:@150236.4]
  assign regs_415_reset = io_reset; // @[:@150237.4 RegFile.scala 76:16:@150244.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@150243.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@150247.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@150241.4]
  assign regs_416_clock = clock; // @[:@150250.4]
  assign regs_416_reset = io_reset; // @[:@150251.4 RegFile.scala 76:16:@150258.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@150257.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@150261.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@150255.4]
  assign regs_417_clock = clock; // @[:@150264.4]
  assign regs_417_reset = io_reset; // @[:@150265.4 RegFile.scala 76:16:@150272.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@150271.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@150275.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@150269.4]
  assign regs_418_clock = clock; // @[:@150278.4]
  assign regs_418_reset = io_reset; // @[:@150279.4 RegFile.scala 76:16:@150286.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@150285.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@150289.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@150283.4]
  assign regs_419_clock = clock; // @[:@150292.4]
  assign regs_419_reset = io_reset; // @[:@150293.4 RegFile.scala 76:16:@150300.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@150299.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@150303.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@150297.4]
  assign regs_420_clock = clock; // @[:@150306.4]
  assign regs_420_reset = io_reset; // @[:@150307.4 RegFile.scala 76:16:@150314.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@150313.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@150317.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@150311.4]
  assign regs_421_clock = clock; // @[:@150320.4]
  assign regs_421_reset = io_reset; // @[:@150321.4 RegFile.scala 76:16:@150328.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@150327.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@150331.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@150325.4]
  assign regs_422_clock = clock; // @[:@150334.4]
  assign regs_422_reset = io_reset; // @[:@150335.4 RegFile.scala 76:16:@150342.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@150341.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@150345.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@150339.4]
  assign regs_423_clock = clock; // @[:@150348.4]
  assign regs_423_reset = io_reset; // @[:@150349.4 RegFile.scala 76:16:@150356.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@150355.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@150359.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@150353.4]
  assign regs_424_clock = clock; // @[:@150362.4]
  assign regs_424_reset = io_reset; // @[:@150363.4 RegFile.scala 76:16:@150370.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@150369.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@150373.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@150367.4]
  assign regs_425_clock = clock; // @[:@150376.4]
  assign regs_425_reset = io_reset; // @[:@150377.4 RegFile.scala 76:16:@150384.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@150383.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@150387.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@150381.4]
  assign regs_426_clock = clock; // @[:@150390.4]
  assign regs_426_reset = io_reset; // @[:@150391.4 RegFile.scala 76:16:@150398.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@150397.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@150401.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@150395.4]
  assign regs_427_clock = clock; // @[:@150404.4]
  assign regs_427_reset = io_reset; // @[:@150405.4 RegFile.scala 76:16:@150412.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@150411.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@150415.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@150409.4]
  assign regs_428_clock = clock; // @[:@150418.4]
  assign regs_428_reset = io_reset; // @[:@150419.4 RegFile.scala 76:16:@150426.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@150425.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@150429.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@150423.4]
  assign regs_429_clock = clock; // @[:@150432.4]
  assign regs_429_reset = io_reset; // @[:@150433.4 RegFile.scala 76:16:@150440.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@150439.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@150443.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@150437.4]
  assign regs_430_clock = clock; // @[:@150446.4]
  assign regs_430_reset = io_reset; // @[:@150447.4 RegFile.scala 76:16:@150454.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@150453.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@150457.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@150451.4]
  assign regs_431_clock = clock; // @[:@150460.4]
  assign regs_431_reset = io_reset; // @[:@150461.4 RegFile.scala 76:16:@150468.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@150467.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@150471.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@150465.4]
  assign regs_432_clock = clock; // @[:@150474.4]
  assign regs_432_reset = io_reset; // @[:@150475.4 RegFile.scala 76:16:@150482.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@150481.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@150485.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@150479.4]
  assign regs_433_clock = clock; // @[:@150488.4]
  assign regs_433_reset = io_reset; // @[:@150489.4 RegFile.scala 76:16:@150496.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@150495.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@150499.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@150493.4]
  assign regs_434_clock = clock; // @[:@150502.4]
  assign regs_434_reset = io_reset; // @[:@150503.4 RegFile.scala 76:16:@150510.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@150509.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@150513.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@150507.4]
  assign regs_435_clock = clock; // @[:@150516.4]
  assign regs_435_reset = io_reset; // @[:@150517.4 RegFile.scala 76:16:@150524.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@150523.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@150527.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@150521.4]
  assign regs_436_clock = clock; // @[:@150530.4]
  assign regs_436_reset = io_reset; // @[:@150531.4 RegFile.scala 76:16:@150538.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@150537.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@150541.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@150535.4]
  assign regs_437_clock = clock; // @[:@150544.4]
  assign regs_437_reset = io_reset; // @[:@150545.4 RegFile.scala 76:16:@150552.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@150551.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@150555.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@150549.4]
  assign regs_438_clock = clock; // @[:@150558.4]
  assign regs_438_reset = io_reset; // @[:@150559.4 RegFile.scala 76:16:@150566.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@150565.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@150569.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@150563.4]
  assign regs_439_clock = clock; // @[:@150572.4]
  assign regs_439_reset = io_reset; // @[:@150573.4 RegFile.scala 76:16:@150580.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@150579.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@150583.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@150577.4]
  assign regs_440_clock = clock; // @[:@150586.4]
  assign regs_440_reset = io_reset; // @[:@150587.4 RegFile.scala 76:16:@150594.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@150593.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@150597.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@150591.4]
  assign regs_441_clock = clock; // @[:@150600.4]
  assign regs_441_reset = io_reset; // @[:@150601.4 RegFile.scala 76:16:@150608.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@150607.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@150611.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@150605.4]
  assign regs_442_clock = clock; // @[:@150614.4]
  assign regs_442_reset = io_reset; // @[:@150615.4 RegFile.scala 76:16:@150622.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@150621.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@150625.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@150619.4]
  assign regs_443_clock = clock; // @[:@150628.4]
  assign regs_443_reset = io_reset; // @[:@150629.4 RegFile.scala 76:16:@150636.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@150635.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@150639.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@150633.4]
  assign regs_444_clock = clock; // @[:@150642.4]
  assign regs_444_reset = io_reset; // @[:@150643.4 RegFile.scala 76:16:@150650.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@150649.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@150653.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@150647.4]
  assign regs_445_clock = clock; // @[:@150656.4]
  assign regs_445_reset = io_reset; // @[:@150657.4 RegFile.scala 76:16:@150664.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@150663.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@150667.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@150661.4]
  assign regs_446_clock = clock; // @[:@150670.4]
  assign regs_446_reset = io_reset; // @[:@150671.4 RegFile.scala 76:16:@150678.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@150677.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@150681.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@150675.4]
  assign regs_447_clock = clock; // @[:@150684.4]
  assign regs_447_reset = io_reset; // @[:@150685.4 RegFile.scala 76:16:@150692.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@150691.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@150695.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@150689.4]
  assign regs_448_clock = clock; // @[:@150698.4]
  assign regs_448_reset = io_reset; // @[:@150699.4 RegFile.scala 76:16:@150706.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@150705.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@150709.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@150703.4]
  assign regs_449_clock = clock; // @[:@150712.4]
  assign regs_449_reset = io_reset; // @[:@150713.4 RegFile.scala 76:16:@150720.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@150719.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@150723.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@150717.4]
  assign regs_450_clock = clock; // @[:@150726.4]
  assign regs_450_reset = io_reset; // @[:@150727.4 RegFile.scala 76:16:@150734.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@150733.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@150737.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@150731.4]
  assign regs_451_clock = clock; // @[:@150740.4]
  assign regs_451_reset = io_reset; // @[:@150741.4 RegFile.scala 76:16:@150748.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@150747.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@150751.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@150745.4]
  assign regs_452_clock = clock; // @[:@150754.4]
  assign regs_452_reset = io_reset; // @[:@150755.4 RegFile.scala 76:16:@150762.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@150761.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@150765.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@150759.4]
  assign regs_453_clock = clock; // @[:@150768.4]
  assign regs_453_reset = io_reset; // @[:@150769.4 RegFile.scala 76:16:@150776.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@150775.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@150779.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@150773.4]
  assign regs_454_clock = clock; // @[:@150782.4]
  assign regs_454_reset = io_reset; // @[:@150783.4 RegFile.scala 76:16:@150790.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@150789.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@150793.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@150787.4]
  assign regs_455_clock = clock; // @[:@150796.4]
  assign regs_455_reset = io_reset; // @[:@150797.4 RegFile.scala 76:16:@150804.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@150803.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@150807.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@150801.4]
  assign regs_456_clock = clock; // @[:@150810.4]
  assign regs_456_reset = io_reset; // @[:@150811.4 RegFile.scala 76:16:@150818.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@150817.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@150821.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@150815.4]
  assign regs_457_clock = clock; // @[:@150824.4]
  assign regs_457_reset = io_reset; // @[:@150825.4 RegFile.scala 76:16:@150832.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@150831.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@150835.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@150829.4]
  assign regs_458_clock = clock; // @[:@150838.4]
  assign regs_458_reset = io_reset; // @[:@150839.4 RegFile.scala 76:16:@150846.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@150845.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@150849.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@150843.4]
  assign regs_459_clock = clock; // @[:@150852.4]
  assign regs_459_reset = io_reset; // @[:@150853.4 RegFile.scala 76:16:@150860.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@150859.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@150863.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@150857.4]
  assign regs_460_clock = clock; // @[:@150866.4]
  assign regs_460_reset = io_reset; // @[:@150867.4 RegFile.scala 76:16:@150874.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@150873.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@150877.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@150871.4]
  assign regs_461_clock = clock; // @[:@150880.4]
  assign regs_461_reset = io_reset; // @[:@150881.4 RegFile.scala 76:16:@150888.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@150887.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@150891.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@150885.4]
  assign regs_462_clock = clock; // @[:@150894.4]
  assign regs_462_reset = io_reset; // @[:@150895.4 RegFile.scala 76:16:@150902.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@150901.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@150905.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@150899.4]
  assign regs_463_clock = clock; // @[:@150908.4]
  assign regs_463_reset = io_reset; // @[:@150909.4 RegFile.scala 76:16:@150916.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@150915.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@150919.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@150913.4]
  assign regs_464_clock = clock; // @[:@150922.4]
  assign regs_464_reset = io_reset; // @[:@150923.4 RegFile.scala 76:16:@150930.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@150929.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@150933.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@150927.4]
  assign regs_465_clock = clock; // @[:@150936.4]
  assign regs_465_reset = io_reset; // @[:@150937.4 RegFile.scala 76:16:@150944.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@150943.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@150947.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@150941.4]
  assign regs_466_clock = clock; // @[:@150950.4]
  assign regs_466_reset = io_reset; // @[:@150951.4 RegFile.scala 76:16:@150958.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@150957.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@150961.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@150955.4]
  assign regs_467_clock = clock; // @[:@150964.4]
  assign regs_467_reset = io_reset; // @[:@150965.4 RegFile.scala 76:16:@150972.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@150971.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@150975.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@150969.4]
  assign regs_468_clock = clock; // @[:@150978.4]
  assign regs_468_reset = io_reset; // @[:@150979.4 RegFile.scala 76:16:@150986.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@150985.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@150989.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@150983.4]
  assign regs_469_clock = clock; // @[:@150992.4]
  assign regs_469_reset = io_reset; // @[:@150993.4 RegFile.scala 76:16:@151000.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@150999.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@151003.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@150997.4]
  assign regs_470_clock = clock; // @[:@151006.4]
  assign regs_470_reset = io_reset; // @[:@151007.4 RegFile.scala 76:16:@151014.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@151013.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@151017.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@151011.4]
  assign regs_471_clock = clock; // @[:@151020.4]
  assign regs_471_reset = io_reset; // @[:@151021.4 RegFile.scala 76:16:@151028.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@151027.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@151031.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@151025.4]
  assign regs_472_clock = clock; // @[:@151034.4]
  assign regs_472_reset = io_reset; // @[:@151035.4 RegFile.scala 76:16:@151042.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@151041.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@151045.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@151039.4]
  assign regs_473_clock = clock; // @[:@151048.4]
  assign regs_473_reset = io_reset; // @[:@151049.4 RegFile.scala 76:16:@151056.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@151055.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@151059.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@151053.4]
  assign regs_474_clock = clock; // @[:@151062.4]
  assign regs_474_reset = io_reset; // @[:@151063.4 RegFile.scala 76:16:@151070.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@151069.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@151073.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@151067.4]
  assign regs_475_clock = clock; // @[:@151076.4]
  assign regs_475_reset = io_reset; // @[:@151077.4 RegFile.scala 76:16:@151084.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@151083.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@151087.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@151081.4]
  assign regs_476_clock = clock; // @[:@151090.4]
  assign regs_476_reset = io_reset; // @[:@151091.4 RegFile.scala 76:16:@151098.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@151097.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@151101.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@151095.4]
  assign regs_477_clock = clock; // @[:@151104.4]
  assign regs_477_reset = io_reset; // @[:@151105.4 RegFile.scala 76:16:@151112.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@151111.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@151115.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@151109.4]
  assign regs_478_clock = clock; // @[:@151118.4]
  assign regs_478_reset = io_reset; // @[:@151119.4 RegFile.scala 76:16:@151126.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@151125.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@151129.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@151123.4]
  assign regs_479_clock = clock; // @[:@151132.4]
  assign regs_479_reset = io_reset; // @[:@151133.4 RegFile.scala 76:16:@151140.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@151139.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@151143.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@151137.4]
  assign regs_480_clock = clock; // @[:@151146.4]
  assign regs_480_reset = io_reset; // @[:@151147.4 RegFile.scala 76:16:@151154.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@151153.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@151157.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@151151.4]
  assign regs_481_clock = clock; // @[:@151160.4]
  assign regs_481_reset = io_reset; // @[:@151161.4 RegFile.scala 76:16:@151168.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@151167.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@151171.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@151165.4]
  assign regs_482_clock = clock; // @[:@151174.4]
  assign regs_482_reset = io_reset; // @[:@151175.4 RegFile.scala 76:16:@151182.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@151181.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@151185.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@151179.4]
  assign regs_483_clock = clock; // @[:@151188.4]
  assign regs_483_reset = io_reset; // @[:@151189.4 RegFile.scala 76:16:@151196.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@151195.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@151199.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@151193.4]
  assign regs_484_clock = clock; // @[:@151202.4]
  assign regs_484_reset = io_reset; // @[:@151203.4 RegFile.scala 76:16:@151210.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@151209.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@151213.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@151207.4]
  assign regs_485_clock = clock; // @[:@151216.4]
  assign regs_485_reset = io_reset; // @[:@151217.4 RegFile.scala 76:16:@151224.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@151223.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@151227.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@151221.4]
  assign regs_486_clock = clock; // @[:@151230.4]
  assign regs_486_reset = io_reset; // @[:@151231.4 RegFile.scala 76:16:@151238.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@151237.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@151241.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@151235.4]
  assign regs_487_clock = clock; // @[:@151244.4]
  assign regs_487_reset = io_reset; // @[:@151245.4 RegFile.scala 76:16:@151252.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@151251.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@151255.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@151249.4]
  assign regs_488_clock = clock; // @[:@151258.4]
  assign regs_488_reset = io_reset; // @[:@151259.4 RegFile.scala 76:16:@151266.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@151265.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@151269.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@151263.4]
  assign regs_489_clock = clock; // @[:@151272.4]
  assign regs_489_reset = io_reset; // @[:@151273.4 RegFile.scala 76:16:@151280.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@151279.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@151283.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@151277.4]
  assign regs_490_clock = clock; // @[:@151286.4]
  assign regs_490_reset = io_reset; // @[:@151287.4 RegFile.scala 76:16:@151294.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@151293.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@151297.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@151291.4]
  assign regs_491_clock = clock; // @[:@151300.4]
  assign regs_491_reset = io_reset; // @[:@151301.4 RegFile.scala 76:16:@151308.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@151307.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@151311.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@151305.4]
  assign regs_492_clock = clock; // @[:@151314.4]
  assign regs_492_reset = io_reset; // @[:@151315.4 RegFile.scala 76:16:@151322.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@151321.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@151325.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@151319.4]
  assign regs_493_clock = clock; // @[:@151328.4]
  assign regs_493_reset = io_reset; // @[:@151329.4 RegFile.scala 76:16:@151336.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@151335.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@151339.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@151333.4]
  assign regs_494_clock = clock; // @[:@151342.4]
  assign regs_494_reset = io_reset; // @[:@151343.4 RegFile.scala 76:16:@151350.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@151349.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@151353.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@151347.4]
  assign regs_495_clock = clock; // @[:@151356.4]
  assign regs_495_reset = io_reset; // @[:@151357.4 RegFile.scala 76:16:@151364.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@151363.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@151367.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@151361.4]
  assign regs_496_clock = clock; // @[:@151370.4]
  assign regs_496_reset = io_reset; // @[:@151371.4 RegFile.scala 76:16:@151378.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@151377.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@151381.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@151375.4]
  assign regs_497_clock = clock; // @[:@151384.4]
  assign regs_497_reset = io_reset; // @[:@151385.4 RegFile.scala 76:16:@151392.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@151391.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@151395.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@151389.4]
  assign regs_498_clock = clock; // @[:@151398.4]
  assign regs_498_reset = io_reset; // @[:@151399.4 RegFile.scala 76:16:@151406.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@151405.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@151409.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@151403.4]
  assign regs_499_clock = clock; // @[:@151412.4]
  assign regs_499_reset = io_reset; // @[:@151413.4 RegFile.scala 76:16:@151420.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@151419.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@151423.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@151417.4]
  assign regs_500_clock = clock; // @[:@151426.4]
  assign regs_500_reset = io_reset; // @[:@151427.4 RegFile.scala 76:16:@151434.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@151433.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@151437.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@151431.4]
  assign regs_501_clock = clock; // @[:@151440.4]
  assign regs_501_reset = io_reset; // @[:@151441.4 RegFile.scala 76:16:@151448.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@151447.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@151451.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@151445.4]
  assign regs_502_clock = clock; // @[:@151454.4]
  assign regs_502_reset = io_reset; // @[:@151455.4 RegFile.scala 76:16:@151462.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@151461.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@151465.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@151459.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@151974.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@151975.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@151976.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@151977.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@151978.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@151979.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@151980.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@151981.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@151982.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@151983.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@151984.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@151985.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@151986.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@151987.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@151988.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@151989.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@151990.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@151991.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@151992.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@151993.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@151994.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@151995.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@151996.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@151997.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@151998.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@151999.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@152000.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@152001.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@152002.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@152003.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@152004.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@152005.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@152006.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@152007.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@152008.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@152009.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@152010.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@152011.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@152012.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@152013.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@152014.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@152015.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@152016.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@152017.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@152018.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@152019.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@152020.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@152021.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@152022.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@152023.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@152024.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@152025.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@152026.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@152027.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@152028.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@152029.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@152030.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@152031.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@152032.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@152033.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@152034.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@152035.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@152036.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@152037.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@152038.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@152039.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@152040.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@152041.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@152042.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@152043.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@152044.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@152045.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@152046.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@152047.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@152048.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@152049.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@152050.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@152051.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@152052.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@152053.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@152054.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@152055.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@152056.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@152057.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@152058.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@152059.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@152060.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@152061.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@152062.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@152063.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@152064.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@152065.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@152066.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@152067.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@152068.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@152069.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@152070.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@152071.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@152072.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@152073.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@152074.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@152075.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@152076.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@152077.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@152078.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@152079.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@152080.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@152081.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@152082.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@152083.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@152084.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@152085.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@152086.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@152087.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@152088.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@152089.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@152090.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@152091.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@152092.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@152093.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@152094.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@152095.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@152096.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@152097.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@152098.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@152099.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@152100.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@152101.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@152102.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@152103.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@152104.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@152105.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@152106.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@152107.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@152108.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@152109.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@152110.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@152111.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@152112.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@152113.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@152114.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@152115.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@152116.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@152117.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@152118.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@152119.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@152120.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@152121.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@152122.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@152123.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@152124.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@152125.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@152126.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@152127.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@152128.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@152129.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@152130.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@152131.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@152132.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@152133.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@152134.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@152135.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@152136.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@152137.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@152138.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@152139.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@152140.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@152141.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@152142.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@152143.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@152144.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@152145.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@152146.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@152147.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@152148.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@152149.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@152150.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@152151.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@152152.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@152153.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@152154.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@152155.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@152156.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@152157.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@152158.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@152159.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@152160.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@152161.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@152162.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@152163.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@152164.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@152165.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@152166.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@152167.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@152168.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@152169.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@152170.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@152171.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@152172.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@152173.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@152174.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@152175.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@152176.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@152177.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@152178.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@152179.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@152180.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@152181.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@152182.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@152183.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@152184.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@152185.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@152186.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@152187.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@152188.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@152189.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@152190.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@152191.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@152192.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@152193.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@152194.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@152195.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@152196.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@152197.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@152198.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@152199.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@152200.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@152201.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@152202.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@152203.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@152204.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@152205.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@152206.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@152207.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@152208.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@152209.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@152210.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@152211.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@152212.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@152213.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@152214.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@152215.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@152216.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@152217.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@152218.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@152219.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@152220.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@152221.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@152222.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@152223.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@152224.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@152225.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@152226.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@152227.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@152228.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@152229.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@152230.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@152231.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@152232.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@152233.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@152234.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@152235.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@152236.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@152237.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@152238.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@152239.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@152240.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@152241.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@152242.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@152243.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@152244.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@152245.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@152246.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@152247.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@152248.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@152249.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@152250.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@152251.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@152252.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@152253.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@152254.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@152255.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@152256.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@152257.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@152258.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@152259.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@152260.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@152261.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@152262.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@152263.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@152264.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@152265.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@152266.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@152267.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@152268.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@152269.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@152270.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@152271.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@152272.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@152273.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@152274.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@152275.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@152276.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@152277.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@152278.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@152279.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@152280.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@152281.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@152282.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@152283.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@152284.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@152285.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@152286.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@152287.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@152288.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@152289.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@152290.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@152291.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@152292.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@152293.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@152294.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@152295.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@152296.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@152297.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@152298.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@152299.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@152300.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@152301.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@152302.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@152303.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@152304.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@152305.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@152306.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@152307.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@152308.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@152309.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@152310.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@152311.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@152312.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@152313.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@152314.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@152315.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@152316.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@152317.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@152318.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@152319.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@152320.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@152321.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@152322.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@152323.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@152324.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@152325.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@152326.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@152327.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@152328.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@152329.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@152330.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@152331.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@152332.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@152333.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@152334.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@152335.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@152336.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@152337.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@152338.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@152339.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@152340.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@152341.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@152342.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@152343.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@152344.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@152345.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@152346.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@152347.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@152348.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@152349.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@152350.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@152351.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@152352.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@152353.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@152354.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@152355.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@152356.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@152357.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@152358.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@152359.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@152360.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@152361.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@152362.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@152363.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@152364.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@152365.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@152366.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@152367.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@152368.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@152369.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@152370.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@152371.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@152372.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@152373.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@152374.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@152375.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@152376.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@152377.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@152378.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@152379.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@152380.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@152381.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@152382.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@152383.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@152384.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@152385.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@152386.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@152387.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@152388.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@152389.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@152390.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@152391.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@152392.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@152393.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@152394.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@152395.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@152396.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@152397.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@152398.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@152399.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@152400.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@152401.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@152402.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@152403.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@152404.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@152405.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@152406.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@152407.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@152408.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@152409.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@152410.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@152411.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@152412.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@152413.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@152414.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@152415.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@152416.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@152417.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@152418.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@152419.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@152420.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@152421.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@152422.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@152423.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@152424.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@152425.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@152426.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@152427.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@152428.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@152429.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@152430.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@152431.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@152432.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@152433.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@152434.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@152435.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@152436.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@152437.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@152438.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@152439.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@152440.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@152441.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@152442.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@152443.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@152444.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@152445.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@152446.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@152447.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@152448.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@152449.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@152450.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@152451.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@152452.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@152453.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@152454.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@152455.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@152456.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@152457.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@152458.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@152459.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@152460.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@152461.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@152462.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@152463.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@152464.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@152465.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@152466.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@152467.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@152468.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@152469.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@152470.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@152471.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@152472.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@152473.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@152474.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@152475.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@152476.4]
  assign rport_io_sel = io_raddr[8:0]; // @[RegFile.scala 106:18:@152477.4]
endmodule
module RetimeWrapper_1012( // @[:@152501.2]
  input         clock, // @[:@152502.4]
  input         reset, // @[:@152503.4]
  input  [39:0] io_in, // @[:@152504.4]
  output [39:0] io_out // @[:@152504.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@152506.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@152506.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@152506.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@152506.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@152506.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@152506.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@152506.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@152519.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@152518.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@152517.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@152516.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@152515.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@152513.4]
endmodule
module FringeFF_503( // @[:@152521.2]
  input         clock, // @[:@152522.4]
  input         reset, // @[:@152523.4]
  input  [39:0] io_in, // @[:@152524.4]
  output [39:0] io_out, // @[:@152524.4]
  input         io_enable // @[:@152524.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@152527.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@152527.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@152527.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@152527.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@152532.4 package.scala 96:25:@152533.4]
  RetimeWrapper_1012 RetimeWrapper ( // @[package.scala 93:22:@152527.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@152532.4 package.scala 96:25:@152533.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@152544.4]
  assign RetimeWrapper_clock = clock; // @[:@152528.4]
  assign RetimeWrapper_reset = reset; // @[:@152529.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@152530.4]
endmodule
module FringeCounter( // @[:@152546.2]
  input   clock, // @[:@152547.4]
  input   reset, // @[:@152548.4]
  input   io_enable, // @[:@152549.4]
  output  io_done // @[:@152549.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@152551.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@152551.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@152551.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@152551.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@152551.4]
  wire [40:0] count; // @[Cat.scala 30:58:@152558.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@152559.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@152560.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@152561.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@152563.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@152551.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@152558.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@152559.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@152560.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@152561.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@152563.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@152574.4]
  assign reg$_clock = clock; // @[:@152552.4]
  assign reg$_reset = reset; // @[:@152553.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@152565.6 FringeCounter.scala 37:15:@152568.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@152556.4]
endmodule
module FringeFF_504( // @[:@152608.2]
  input   clock, // @[:@152609.4]
  input   reset, // @[:@152610.4]
  input   io_in, // @[:@152611.4]
  input   io_reset, // @[:@152611.4]
  output  io_out, // @[:@152611.4]
  input   io_enable // @[:@152611.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@152614.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@152614.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@152614.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@152614.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@152614.4]
  wire  _T_18; // @[package.scala 96:25:@152619.4 package.scala 96:25:@152620.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@152625.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@152614.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@152619.4 package.scala 96:25:@152620.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@152625.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@152631.4]
  assign RetimeWrapper_clock = clock; // @[:@152615.4]
  assign RetimeWrapper_reset = reset; // @[:@152616.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@152618.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@152617.4]
endmodule
module Depulser( // @[:@152633.2]
  input   clock, // @[:@152634.4]
  input   reset, // @[:@152635.4]
  input   io_in, // @[:@152636.4]
  input   io_rst, // @[:@152636.4]
  output  io_out // @[:@152636.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@152638.4]
  wire  r_reset; // @[Depulser.scala 14:17:@152638.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@152638.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@152638.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@152638.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@152638.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@152638.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@152647.4]
  assign r_clock = clock; // @[:@152639.4]
  assign r_reset = reset; // @[:@152640.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@152642.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@152646.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@152645.4]
endmodule
module Fringe( // @[:@152649.2]
  input         clock, // @[:@152650.4]
  input         reset, // @[:@152651.4]
  input  [31:0] io_raddr, // @[:@152652.4]
  input         io_wen, // @[:@152652.4]
  input  [31:0] io_waddr, // @[:@152652.4]
  input  [63:0] io_wdata, // @[:@152652.4]
  output [63:0] io_rdata, // @[:@152652.4]
  output        io_enable, // @[:@152652.4]
  input         io_done, // @[:@152652.4]
  output        io_reset, // @[:@152652.4]
  output [63:0] io_argIns_0, // @[:@152652.4]
  output [63:0] io_argIns_1, // @[:@152652.4]
  input         io_argOuts_0_valid, // @[:@152652.4]
  input  [63:0] io_argOuts_0_bits, // @[:@152652.4]
  output        io_memStreams_stores_0_cmd_ready, // @[:@152652.4]
  input         io_memStreams_stores_0_cmd_valid, // @[:@152652.4]
  input  [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@152652.4]
  input  [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@152652.4]
  output        io_memStreams_stores_0_data_ready, // @[:@152652.4]
  input         io_memStreams_stores_0_data_valid, // @[:@152652.4]
  input  [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@152652.4]
  input         io_memStreams_stores_0_data_bits_wstrb, // @[:@152652.4]
  input         io_memStreams_stores_0_wresp_ready, // @[:@152652.4]
  output        io_memStreams_stores_0_wresp_valid, // @[:@152652.4]
  output        io_memStreams_stores_0_wresp_bits, // @[:@152652.4]
  input         io_dram_0_cmd_ready, // @[:@152652.4]
  output        io_dram_0_cmd_valid, // @[:@152652.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@152652.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@152652.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@152652.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@152652.4]
  input         io_dram_0_wdata_ready, // @[:@152652.4]
  output        io_dram_0_wdata_valid, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_0, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_1, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_2, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_3, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_4, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_5, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_6, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_7, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_8, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_9, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_10, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_11, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_12, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_13, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_14, // @[:@152652.4]
  output [31:0] io_dram_0_wdata_bits_wdata_15, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@152652.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@152652.4]
  output        io_dram_0_rresp_ready, // @[:@152652.4]
  output        io_dram_0_wresp_ready, // @[:@152652.4]
  input         io_dram_0_wresp_valid, // @[:@152652.4]
  input  [31:0] io_dram_0_wresp_bits_tag, // @[:@152652.4]
  input         io_dram_1_cmd_ready, // @[:@152652.4]
  output        io_dram_1_cmd_valid, // @[:@152652.4]
  output [63:0] io_dram_1_cmd_bits_addr, // @[:@152652.4]
  output [31:0] io_dram_1_cmd_bits_size, // @[:@152652.4]
  output        io_dram_1_cmd_bits_isWr, // @[:@152652.4]
  output [31:0] io_dram_1_cmd_bits_tag, // @[:@152652.4]
  input         io_dram_1_wdata_ready, // @[:@152652.4]
  output        io_dram_1_wdata_valid, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_0, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_1, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_2, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_3, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_4, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_5, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_6, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_7, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_8, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_9, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_10, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_11, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_12, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_13, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_14, // @[:@152652.4]
  output [31:0] io_dram_1_wdata_bits_wdata_15, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_0, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_1, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_2, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_3, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_4, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_5, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_6, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_7, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_8, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_9, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_10, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_11, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_12, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_13, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_14, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_15, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_16, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_17, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_18, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_19, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_20, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_21, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_22, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_23, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_24, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_25, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_26, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_27, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_28, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_29, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_30, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_31, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_32, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_33, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_34, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_35, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_36, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_37, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_38, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_39, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_40, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_41, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_42, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_43, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_44, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_45, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_46, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_47, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_48, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_49, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_50, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_51, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_52, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_53, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_54, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_55, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_56, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_57, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_58, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_59, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_60, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_61, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_62, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wstrb_63, // @[:@152652.4]
  output        io_dram_1_wdata_bits_wlast, // @[:@152652.4]
  output        io_dram_1_rresp_ready, // @[:@152652.4]
  output        io_dram_1_wresp_ready, // @[:@152652.4]
  input         io_dram_1_wresp_valid, // @[:@152652.4]
  input  [31:0] io_dram_1_wresp_bits_tag, // @[:@152652.4]
  input         io_dram_2_cmd_ready, // @[:@152652.4]
  output        io_dram_2_cmd_valid, // @[:@152652.4]
  output [63:0] io_dram_2_cmd_bits_addr, // @[:@152652.4]
  output [31:0] io_dram_2_cmd_bits_size, // @[:@152652.4]
  output        io_dram_2_cmd_bits_isWr, // @[:@152652.4]
  output [31:0] io_dram_2_cmd_bits_tag, // @[:@152652.4]
  input         io_dram_2_wdata_ready, // @[:@152652.4]
  output        io_dram_2_wdata_valid, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_0, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_1, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_2, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_3, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_4, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_5, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_6, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_7, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_8, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_9, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_10, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_11, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_12, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_13, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_14, // @[:@152652.4]
  output [31:0] io_dram_2_wdata_bits_wdata_15, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_0, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_1, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_2, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_3, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_4, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_5, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_6, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_7, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_8, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_9, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_10, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_11, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_12, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_13, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_14, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_15, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_16, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_17, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_18, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_19, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_20, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_21, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_22, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_23, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_24, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_25, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_26, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_27, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_28, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_29, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_30, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_31, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_32, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_33, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_34, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_35, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_36, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_37, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_38, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_39, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_40, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_41, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_42, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_43, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_44, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_45, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_46, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_47, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_48, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_49, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_50, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_51, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_52, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_53, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_54, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_55, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_56, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_57, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_58, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_59, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_60, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_61, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_62, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wstrb_63, // @[:@152652.4]
  output        io_dram_2_wdata_bits_wlast, // @[:@152652.4]
  output        io_dram_2_rresp_ready, // @[:@152652.4]
  output        io_dram_2_wresp_ready, // @[:@152652.4]
  input         io_dram_2_wresp_valid, // @[:@152652.4]
  input  [31:0] io_dram_2_wresp_bits_tag, // @[:@152652.4]
  input         io_dram_3_cmd_ready, // @[:@152652.4]
  output        io_dram_3_cmd_valid, // @[:@152652.4]
  output [63:0] io_dram_3_cmd_bits_addr, // @[:@152652.4]
  output [31:0] io_dram_3_cmd_bits_size, // @[:@152652.4]
  output        io_dram_3_cmd_bits_isWr, // @[:@152652.4]
  output [31:0] io_dram_3_cmd_bits_tag, // @[:@152652.4]
  input         io_dram_3_wdata_ready, // @[:@152652.4]
  output        io_dram_3_wdata_valid, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_0, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_1, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_2, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_3, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_4, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_5, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_6, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_7, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_8, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_9, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_10, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_11, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_12, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_13, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_14, // @[:@152652.4]
  output [31:0] io_dram_3_wdata_bits_wdata_15, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_0, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_1, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_2, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_3, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_4, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_5, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_6, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_7, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_8, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_9, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_10, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_11, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_12, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_13, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_14, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_15, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_16, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_17, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_18, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_19, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_20, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_21, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_22, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_23, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_24, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_25, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_26, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_27, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_28, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_29, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_30, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_31, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_32, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_33, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_34, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_35, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_36, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_37, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_38, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_39, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_40, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_41, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_42, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_43, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_44, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_45, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_46, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_47, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_48, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_49, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_50, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_51, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_52, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_53, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_54, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_55, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_56, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_57, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_58, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_59, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_60, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_61, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_62, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wstrb_63, // @[:@152652.4]
  output        io_dram_3_wdata_bits_wlast, // @[:@152652.4]
  output        io_dram_3_rresp_ready, // @[:@152652.4]
  output        io_dram_3_wresp_ready, // @[:@152652.4]
  input         io_dram_3_wresp_valid, // @[:@152652.4]
  input  [31:0] io_dram_3_wresp_bits_tag, // @[:@152652.4]
  input         io_heap_0_req_valid, // @[:@152652.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@152652.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@152652.4]
  output        io_heap_0_resp_valid, // @[:@152652.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@152652.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@152652.4]
);
  wire  dramArbs_0_clock; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_reset; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_enable; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@152658.4]
  wire [63:0] dramArbs_0_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_app_stores_0_wresp_ready; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_cmd_ready; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 91:25:@152658.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_ready; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_0_io_dram_wresp_valid; // @[Fringe.scala 91:25:@152658.4]
  wire [31:0] dramArbs_0_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@152658.4]
  wire  dramArbs_1_clock; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_reset; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_enable; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_cmd_ready; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 91:25:@153651.4]
  wire [63:0] dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_ready; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_1_io_dram_wresp_valid; // @[Fringe.scala 91:25:@153651.4]
  wire [31:0] dramArbs_1_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@153651.4]
  wire  dramArbs_2_clock; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_reset; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_enable; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_cmd_ready; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 91:25:@154611.4]
  wire [63:0] dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_ready; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_2_io_dram_wresp_valid; // @[Fringe.scala 91:25:@154611.4]
  wire [31:0] dramArbs_2_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@154611.4]
  wire  dramArbs_3_clock; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_reset; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_enable; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_cmd_ready; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 91:25:@155571.4]
  wire [63:0] dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_ready; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 91:25:@155571.4]
  wire  dramArbs_3_io_dram_wresp_valid; // @[Fringe.scala 91:25:@155571.4]
  wire [31:0] dramArbs_3_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@155571.4]
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@156531.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@156531.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@156531.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@156531.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@156531.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@156531.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@156531.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@156531.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@156531.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@156531.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@156531.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@156531.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@156540.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@156540.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@156540.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@156540.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@156540.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@156540.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@156540.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@156540.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@156540.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@156540.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@156540.4]
  wire [63:0] regs_io_argIns_3; // @[Fringe.scala 116:20:@156540.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@156540.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@156540.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@156540.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@156540.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@158590.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@158590.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@158590.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@158590.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@158609.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@158609.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@158609.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@158609.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@158609.4]
  wire [63:0] _T_1020; // @[:@158567.4 :@158568.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@158569.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@158571.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@158573.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@158575.4]
  wire  _T_1025; // @[Fringe.scala 134:28:@158577.4]
  wire  _T_1029; // @[Fringe.scala 134:42:@158579.4]
  wire  _T_1030; // @[Fringe.scala 135:27:@158581.4]
  wire [63:0] _T_1040; // @[Fringe.scala 156:22:@158617.4]
  reg  _T_1047; // @[package.scala 152:20:@158620.4]
  reg [31:0] _RAND_0;
  wire  _T_1048; // @[package.scala 153:13:@158622.4]
  wire  _T_1049; // @[package.scala 153:8:@158623.4]
  wire  _T_1052; // @[Fringe.scala 160:55:@158627.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@158628.4]
  wire  _T_1055; // @[Fringe.scala 161:58:@158631.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@158632.4]
  wire [1:0] _T_1059; // @[Fringe.scala 162:57:@158634.4]
  wire [1:0] _T_1061; // @[Fringe.scala 162:34:@158635.4]
  wire [63:0] _T_1063; // @[Fringe.scala 163:30:@158637.4]
  wire [1:0] _T_1064; // @[Fringe.scala 171:37:@158640.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@158619.4 Fringe.scala 163:24:@158638.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@158619.4 Fringe.scala 162:28:@158636.4]
  wire [61:0] _T_1065; // @[Fringe.scala 171:37:@158641.4]
  wire  alloc; // @[Fringe.scala 202:38:@160271.4]
  wire  dealloc; // @[Fringe.scala 203:40:@160272.4]
  wire  _T_1569; // @[Fringe.scala 204:37:@160273.4]
  reg  _T_1572; // @[package.scala 152:20:@160274.4]
  reg [31:0] _RAND_1;
  wire  _T_1573; // @[package.scala 153:13:@160276.4]
  DRAMArbiter dramArbs_0 ( // @[Fringe.scala 91:25:@152658.4]
    .clock(dramArbs_0_clock),
    .reset(dramArbs_0_reset),
    .io_enable(dramArbs_0_io_enable),
    .io_app_stores_0_cmd_ready(dramArbs_0_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_0_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_0_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_0_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_0_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_0_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_0_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_0_io_app_stores_0_data_bits_wstrb),
    .io_app_stores_0_wresp_ready(dramArbs_0_io_app_stores_0_wresp_ready),
    .io_app_stores_0_wresp_valid(dramArbs_0_io_app_stores_0_wresp_valid),
    .io_app_stores_0_wresp_bits(dramArbs_0_io_app_stores_0_wresp_bits),
    .io_dram_cmd_ready(dramArbs_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_0_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_0_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_0_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_0_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_0_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_0_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_0_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_0_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_0_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_0_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_0_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_0_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_0_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_0_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_0_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_0_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_0_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_0_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_0_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_0_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_0_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_0_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_0_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_0_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_0_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_0_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_0_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_0_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_0_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_0_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_0_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_0_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_0_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_0_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_0_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_0_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_0_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_0_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_0_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_0_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_0_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_0_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_0_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_0_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_0_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_0_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_0_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_0_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_0_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_0_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_0_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_0_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_0_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_0_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_0_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_0_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_0_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_0_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_0_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_0_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_0_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_0_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_0_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_0_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_0_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_0_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_0_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_0_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_0_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_0_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_0_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_0_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_0_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_0_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_1 ( // @[Fringe.scala 91:25:@153651.4]
    .clock(dramArbs_1_clock),
    .reset(dramArbs_1_reset),
    .io_enable(dramArbs_1_io_enable),
    .io_dram_cmd_ready(dramArbs_1_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_1_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_1_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_1_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_1_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_1_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_1_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_1_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_1_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_1_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_1_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_1_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_1_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_1_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_1_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_1_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_1_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_1_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_1_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_1_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_1_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_1_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_1_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_1_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_1_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_1_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_1_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_1_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_1_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_1_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_1_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_1_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_1_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_1_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_1_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_1_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_1_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_1_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_1_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_1_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_1_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_1_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_1_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_1_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_1_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_1_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_1_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_1_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_1_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_1_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_1_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_1_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_1_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_1_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_1_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_1_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_1_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_1_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_1_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_1_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_1_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_1_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_1_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_1_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_1_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_1_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_1_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_1_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_1_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_1_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_1_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_1_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_1_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_1_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_1_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_1_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_1_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_1_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_1_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_1_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_1_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_1_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_1_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_1_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_1_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_1_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_1_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_1_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_1_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_1_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_1_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_1_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_1_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_2 ( // @[Fringe.scala 91:25:@154611.4]
    .clock(dramArbs_2_clock),
    .reset(dramArbs_2_reset),
    .io_enable(dramArbs_2_io_enable),
    .io_dram_cmd_ready(dramArbs_2_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_2_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_2_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_2_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_2_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_2_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_2_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_2_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_2_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_2_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_2_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_2_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_2_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_2_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_2_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_2_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_2_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_2_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_2_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_2_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_2_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_2_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_2_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_2_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_2_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_2_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_2_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_2_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_2_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_2_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_2_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_2_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_2_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_2_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_2_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_2_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_2_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_2_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_2_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_2_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_2_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_2_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_2_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_2_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_2_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_2_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_2_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_2_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_2_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_2_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_2_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_2_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_2_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_2_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_2_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_2_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_2_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_2_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_2_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_2_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_2_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_2_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_2_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_2_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_2_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_2_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_2_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_2_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_2_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_2_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_2_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_2_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_2_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_2_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_2_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_2_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_2_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_2_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_2_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_2_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_2_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_2_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_2_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_2_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_2_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_2_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_2_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_2_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_2_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_2_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_2_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_2_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_2_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_3 ( // @[Fringe.scala 91:25:@155571.4]
    .clock(dramArbs_3_clock),
    .reset(dramArbs_3_reset),
    .io_enable(dramArbs_3_io_enable),
    .io_dram_cmd_ready(dramArbs_3_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_3_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_3_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_3_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_3_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_3_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_3_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_3_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_3_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_3_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_3_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_3_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_3_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_3_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_3_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_3_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_3_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_3_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_3_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_3_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_3_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_3_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_3_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_3_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_3_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_3_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_3_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_3_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_3_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_3_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_3_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_3_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_3_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_3_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_3_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_3_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_3_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_3_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_3_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_3_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_3_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_3_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_3_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_3_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_3_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_3_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_3_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_3_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_3_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_3_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_3_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_3_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_3_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_3_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_3_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_3_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_3_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_3_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_3_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_3_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_3_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_3_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_3_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_3_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_3_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_3_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_3_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_3_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_3_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_3_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_3_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_3_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_3_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_3_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_3_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_3_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_3_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_3_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_3_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_3_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_3_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_3_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_3_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_3_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_3_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_3_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_3_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_3_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_3_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_3_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_3_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_3_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_3_io_dram_wresp_bits_tag)
  );
  DRAMHeap heap ( // @[Fringe.scala 107:20:@156531.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@156540.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@158590.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@158609.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_1020 = regs_io_argIns_1; // @[:@158567.4 :@158568.4]
  assign curStatus_done = _T_1020[0]; // @[Fringe.scala 133:45:@158569.4]
  assign curStatus_timeout = _T_1020[1]; // @[Fringe.scala 133:45:@158571.4]
  assign curStatus_allocDealloc = _T_1020[4:2]; // @[Fringe.scala 133:45:@158573.4]
  assign curStatus_sizeAddr = _T_1020[63:5]; // @[Fringe.scala 133:45:@158575.4]
  assign _T_1025 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@158577.4]
  assign _T_1029 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@158579.4]
  assign _T_1030 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@158581.4]
  assign _T_1040 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@158617.4]
  assign _T_1048 = _T_1047 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@158622.4]
  assign _T_1049 = heap_io_host_0_req_valid & _T_1048; // @[package.scala 153:8:@158623.4]
  assign _T_1052 = _T_1025 & depulser_io_out; // @[Fringe.scala 160:55:@158627.4]
  assign status_bits_done = depulser_io_out ? _T_1052 : curStatus_done; // @[Fringe.scala 160:26:@158628.4]
  assign _T_1055 = _T_1025 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@158631.4]
  assign status_bits_timeout = depulser_io_out ? _T_1055 : curStatus_timeout; // @[Fringe.scala 161:29:@158632.4]
  assign _T_1059 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@158634.4]
  assign _T_1061 = heap_io_host_0_req_valid ? _T_1059 : 2'h0; // @[Fringe.scala 162:34:@158635.4]
  assign _T_1063 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@158637.4]
  assign _T_1064 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@158640.4]
  assign status_bits_sizeAddr = _T_1063[58:0]; // @[Fringe.scala 158:20:@158619.4 Fringe.scala 163:24:@158638.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_1061}; // @[Fringe.scala 158:20:@158619.4 Fringe.scala 162:28:@158636.4]
  assign _T_1065 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@158641.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@160271.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@160272.4]
  assign _T_1569 = alloc | dealloc; // @[Fringe.scala 204:37:@160273.4]
  assign _T_1573 = _T_1572 ^ _T_1569; // @[package.scala 153:13:@160276.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@158565.4]
  assign io_enable = _T_1025 & _T_1029; // @[Fringe.scala 136:13:@158585.4]
  assign io_reset = _T_1030 | reset; // @[Fringe.scala 137:12:@158586.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@158607.4]
  assign io_argIns_1 = regs_io_argIns_3; // @[Fringe.scala 151:51:@158608.4]
  assign io_memStreams_stores_0_cmd_ready = dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 101:72:@153577.4]
  assign io_memStreams_stores_0_data_ready = dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 101:72:@153573.4]
  assign io_memStreams_stores_0_wresp_valid = dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 101:72:@153568.4]
  assign io_memStreams_stores_0_wresp_bits = dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 101:72:@153567.4]
  assign io_dram_0_cmd_valid = dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 195:72:@159769.4]
  assign io_dram_0_cmd_bits_addr = dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@159768.4]
  assign io_dram_0_cmd_bits_size = dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@159767.4]
  assign io_dram_0_cmd_bits_isWr = dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@159765.4]
  assign io_dram_0_cmd_bits_tag = dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@159764.4]
  assign io_dram_0_wdata_valid = dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 195:72:@159762.4]
  assign io_dram_0_wdata_bits_wdata_0 = dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@159746.4]
  assign io_dram_0_wdata_bits_wdata_1 = dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@159747.4]
  assign io_dram_0_wdata_bits_wdata_2 = dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@159748.4]
  assign io_dram_0_wdata_bits_wdata_3 = dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@159749.4]
  assign io_dram_0_wdata_bits_wdata_4 = dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@159750.4]
  assign io_dram_0_wdata_bits_wdata_5 = dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@159751.4]
  assign io_dram_0_wdata_bits_wdata_6 = dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@159752.4]
  assign io_dram_0_wdata_bits_wdata_7 = dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@159753.4]
  assign io_dram_0_wdata_bits_wdata_8 = dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@159754.4]
  assign io_dram_0_wdata_bits_wdata_9 = dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@159755.4]
  assign io_dram_0_wdata_bits_wdata_10 = dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@159756.4]
  assign io_dram_0_wdata_bits_wdata_11 = dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@159757.4]
  assign io_dram_0_wdata_bits_wdata_12 = dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@159758.4]
  assign io_dram_0_wdata_bits_wdata_13 = dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@159759.4]
  assign io_dram_0_wdata_bits_wdata_14 = dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@159760.4]
  assign io_dram_0_wdata_bits_wdata_15 = dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@159761.4]
  assign io_dram_0_wdata_bits_wstrb_0 = dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@159682.4]
  assign io_dram_0_wdata_bits_wstrb_1 = dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@159683.4]
  assign io_dram_0_wdata_bits_wstrb_2 = dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@159684.4]
  assign io_dram_0_wdata_bits_wstrb_3 = dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@159685.4]
  assign io_dram_0_wdata_bits_wstrb_4 = dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@159686.4]
  assign io_dram_0_wdata_bits_wstrb_5 = dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@159687.4]
  assign io_dram_0_wdata_bits_wstrb_6 = dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@159688.4]
  assign io_dram_0_wdata_bits_wstrb_7 = dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@159689.4]
  assign io_dram_0_wdata_bits_wstrb_8 = dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@159690.4]
  assign io_dram_0_wdata_bits_wstrb_9 = dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@159691.4]
  assign io_dram_0_wdata_bits_wstrb_10 = dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@159692.4]
  assign io_dram_0_wdata_bits_wstrb_11 = dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@159693.4]
  assign io_dram_0_wdata_bits_wstrb_12 = dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@159694.4]
  assign io_dram_0_wdata_bits_wstrb_13 = dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@159695.4]
  assign io_dram_0_wdata_bits_wstrb_14 = dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@159696.4]
  assign io_dram_0_wdata_bits_wstrb_15 = dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@159697.4]
  assign io_dram_0_wdata_bits_wstrb_16 = dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@159698.4]
  assign io_dram_0_wdata_bits_wstrb_17 = dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@159699.4]
  assign io_dram_0_wdata_bits_wstrb_18 = dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@159700.4]
  assign io_dram_0_wdata_bits_wstrb_19 = dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@159701.4]
  assign io_dram_0_wdata_bits_wstrb_20 = dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@159702.4]
  assign io_dram_0_wdata_bits_wstrb_21 = dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@159703.4]
  assign io_dram_0_wdata_bits_wstrb_22 = dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@159704.4]
  assign io_dram_0_wdata_bits_wstrb_23 = dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@159705.4]
  assign io_dram_0_wdata_bits_wstrb_24 = dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@159706.4]
  assign io_dram_0_wdata_bits_wstrb_25 = dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@159707.4]
  assign io_dram_0_wdata_bits_wstrb_26 = dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@159708.4]
  assign io_dram_0_wdata_bits_wstrb_27 = dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@159709.4]
  assign io_dram_0_wdata_bits_wstrb_28 = dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@159710.4]
  assign io_dram_0_wdata_bits_wstrb_29 = dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@159711.4]
  assign io_dram_0_wdata_bits_wstrb_30 = dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@159712.4]
  assign io_dram_0_wdata_bits_wstrb_31 = dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@159713.4]
  assign io_dram_0_wdata_bits_wstrb_32 = dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@159714.4]
  assign io_dram_0_wdata_bits_wstrb_33 = dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@159715.4]
  assign io_dram_0_wdata_bits_wstrb_34 = dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@159716.4]
  assign io_dram_0_wdata_bits_wstrb_35 = dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@159717.4]
  assign io_dram_0_wdata_bits_wstrb_36 = dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@159718.4]
  assign io_dram_0_wdata_bits_wstrb_37 = dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@159719.4]
  assign io_dram_0_wdata_bits_wstrb_38 = dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@159720.4]
  assign io_dram_0_wdata_bits_wstrb_39 = dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@159721.4]
  assign io_dram_0_wdata_bits_wstrb_40 = dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@159722.4]
  assign io_dram_0_wdata_bits_wstrb_41 = dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@159723.4]
  assign io_dram_0_wdata_bits_wstrb_42 = dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@159724.4]
  assign io_dram_0_wdata_bits_wstrb_43 = dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@159725.4]
  assign io_dram_0_wdata_bits_wstrb_44 = dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@159726.4]
  assign io_dram_0_wdata_bits_wstrb_45 = dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@159727.4]
  assign io_dram_0_wdata_bits_wstrb_46 = dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@159728.4]
  assign io_dram_0_wdata_bits_wstrb_47 = dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@159729.4]
  assign io_dram_0_wdata_bits_wstrb_48 = dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@159730.4]
  assign io_dram_0_wdata_bits_wstrb_49 = dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@159731.4]
  assign io_dram_0_wdata_bits_wstrb_50 = dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@159732.4]
  assign io_dram_0_wdata_bits_wstrb_51 = dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@159733.4]
  assign io_dram_0_wdata_bits_wstrb_52 = dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@159734.4]
  assign io_dram_0_wdata_bits_wstrb_53 = dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@159735.4]
  assign io_dram_0_wdata_bits_wstrb_54 = dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@159736.4]
  assign io_dram_0_wdata_bits_wstrb_55 = dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@159737.4]
  assign io_dram_0_wdata_bits_wstrb_56 = dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@159738.4]
  assign io_dram_0_wdata_bits_wstrb_57 = dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@159739.4]
  assign io_dram_0_wdata_bits_wstrb_58 = dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@159740.4]
  assign io_dram_0_wdata_bits_wstrb_59 = dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@159741.4]
  assign io_dram_0_wdata_bits_wstrb_60 = dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@159742.4]
  assign io_dram_0_wdata_bits_wstrb_61 = dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@159743.4]
  assign io_dram_0_wdata_bits_wstrb_62 = dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@159744.4]
  assign io_dram_0_wdata_bits_wstrb_63 = dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@159745.4]
  assign io_dram_0_wdata_bits_wlast = dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@159681.4]
  assign io_dram_0_rresp_ready = dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 195:72:@159680.4]
  assign io_dram_0_wresp_ready = dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 195:72:@159661.4]
  assign io_dram_1_cmd_valid = dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 195:72:@159881.4]
  assign io_dram_1_cmd_bits_addr = dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@159880.4]
  assign io_dram_1_cmd_bits_size = dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@159879.4]
  assign io_dram_1_cmd_bits_isWr = dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@159877.4]
  assign io_dram_1_cmd_bits_tag = dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@159876.4]
  assign io_dram_1_wdata_valid = dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 195:72:@159874.4]
  assign io_dram_1_wdata_bits_wdata_0 = dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@159858.4]
  assign io_dram_1_wdata_bits_wdata_1 = dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@159859.4]
  assign io_dram_1_wdata_bits_wdata_2 = dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@159860.4]
  assign io_dram_1_wdata_bits_wdata_3 = dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@159861.4]
  assign io_dram_1_wdata_bits_wdata_4 = dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@159862.4]
  assign io_dram_1_wdata_bits_wdata_5 = dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@159863.4]
  assign io_dram_1_wdata_bits_wdata_6 = dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@159864.4]
  assign io_dram_1_wdata_bits_wdata_7 = dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@159865.4]
  assign io_dram_1_wdata_bits_wdata_8 = dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@159866.4]
  assign io_dram_1_wdata_bits_wdata_9 = dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@159867.4]
  assign io_dram_1_wdata_bits_wdata_10 = dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@159868.4]
  assign io_dram_1_wdata_bits_wdata_11 = dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@159869.4]
  assign io_dram_1_wdata_bits_wdata_12 = dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@159870.4]
  assign io_dram_1_wdata_bits_wdata_13 = dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@159871.4]
  assign io_dram_1_wdata_bits_wdata_14 = dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@159872.4]
  assign io_dram_1_wdata_bits_wdata_15 = dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@159873.4]
  assign io_dram_1_wdata_bits_wstrb_0 = dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@159794.4]
  assign io_dram_1_wdata_bits_wstrb_1 = dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@159795.4]
  assign io_dram_1_wdata_bits_wstrb_2 = dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@159796.4]
  assign io_dram_1_wdata_bits_wstrb_3 = dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@159797.4]
  assign io_dram_1_wdata_bits_wstrb_4 = dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@159798.4]
  assign io_dram_1_wdata_bits_wstrb_5 = dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@159799.4]
  assign io_dram_1_wdata_bits_wstrb_6 = dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@159800.4]
  assign io_dram_1_wdata_bits_wstrb_7 = dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@159801.4]
  assign io_dram_1_wdata_bits_wstrb_8 = dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@159802.4]
  assign io_dram_1_wdata_bits_wstrb_9 = dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@159803.4]
  assign io_dram_1_wdata_bits_wstrb_10 = dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@159804.4]
  assign io_dram_1_wdata_bits_wstrb_11 = dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@159805.4]
  assign io_dram_1_wdata_bits_wstrb_12 = dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@159806.4]
  assign io_dram_1_wdata_bits_wstrb_13 = dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@159807.4]
  assign io_dram_1_wdata_bits_wstrb_14 = dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@159808.4]
  assign io_dram_1_wdata_bits_wstrb_15 = dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@159809.4]
  assign io_dram_1_wdata_bits_wstrb_16 = dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@159810.4]
  assign io_dram_1_wdata_bits_wstrb_17 = dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@159811.4]
  assign io_dram_1_wdata_bits_wstrb_18 = dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@159812.4]
  assign io_dram_1_wdata_bits_wstrb_19 = dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@159813.4]
  assign io_dram_1_wdata_bits_wstrb_20 = dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@159814.4]
  assign io_dram_1_wdata_bits_wstrb_21 = dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@159815.4]
  assign io_dram_1_wdata_bits_wstrb_22 = dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@159816.4]
  assign io_dram_1_wdata_bits_wstrb_23 = dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@159817.4]
  assign io_dram_1_wdata_bits_wstrb_24 = dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@159818.4]
  assign io_dram_1_wdata_bits_wstrb_25 = dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@159819.4]
  assign io_dram_1_wdata_bits_wstrb_26 = dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@159820.4]
  assign io_dram_1_wdata_bits_wstrb_27 = dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@159821.4]
  assign io_dram_1_wdata_bits_wstrb_28 = dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@159822.4]
  assign io_dram_1_wdata_bits_wstrb_29 = dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@159823.4]
  assign io_dram_1_wdata_bits_wstrb_30 = dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@159824.4]
  assign io_dram_1_wdata_bits_wstrb_31 = dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@159825.4]
  assign io_dram_1_wdata_bits_wstrb_32 = dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@159826.4]
  assign io_dram_1_wdata_bits_wstrb_33 = dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@159827.4]
  assign io_dram_1_wdata_bits_wstrb_34 = dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@159828.4]
  assign io_dram_1_wdata_bits_wstrb_35 = dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@159829.4]
  assign io_dram_1_wdata_bits_wstrb_36 = dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@159830.4]
  assign io_dram_1_wdata_bits_wstrb_37 = dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@159831.4]
  assign io_dram_1_wdata_bits_wstrb_38 = dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@159832.4]
  assign io_dram_1_wdata_bits_wstrb_39 = dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@159833.4]
  assign io_dram_1_wdata_bits_wstrb_40 = dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@159834.4]
  assign io_dram_1_wdata_bits_wstrb_41 = dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@159835.4]
  assign io_dram_1_wdata_bits_wstrb_42 = dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@159836.4]
  assign io_dram_1_wdata_bits_wstrb_43 = dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@159837.4]
  assign io_dram_1_wdata_bits_wstrb_44 = dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@159838.4]
  assign io_dram_1_wdata_bits_wstrb_45 = dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@159839.4]
  assign io_dram_1_wdata_bits_wstrb_46 = dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@159840.4]
  assign io_dram_1_wdata_bits_wstrb_47 = dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@159841.4]
  assign io_dram_1_wdata_bits_wstrb_48 = dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@159842.4]
  assign io_dram_1_wdata_bits_wstrb_49 = dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@159843.4]
  assign io_dram_1_wdata_bits_wstrb_50 = dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@159844.4]
  assign io_dram_1_wdata_bits_wstrb_51 = dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@159845.4]
  assign io_dram_1_wdata_bits_wstrb_52 = dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@159846.4]
  assign io_dram_1_wdata_bits_wstrb_53 = dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@159847.4]
  assign io_dram_1_wdata_bits_wstrb_54 = dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@159848.4]
  assign io_dram_1_wdata_bits_wstrb_55 = dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@159849.4]
  assign io_dram_1_wdata_bits_wstrb_56 = dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@159850.4]
  assign io_dram_1_wdata_bits_wstrb_57 = dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@159851.4]
  assign io_dram_1_wdata_bits_wstrb_58 = dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@159852.4]
  assign io_dram_1_wdata_bits_wstrb_59 = dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@159853.4]
  assign io_dram_1_wdata_bits_wstrb_60 = dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@159854.4]
  assign io_dram_1_wdata_bits_wstrb_61 = dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@159855.4]
  assign io_dram_1_wdata_bits_wstrb_62 = dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@159856.4]
  assign io_dram_1_wdata_bits_wstrb_63 = dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@159857.4]
  assign io_dram_1_wdata_bits_wlast = dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@159793.4]
  assign io_dram_1_rresp_ready = dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 195:72:@159792.4]
  assign io_dram_1_wresp_ready = dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 195:72:@159773.4]
  assign io_dram_2_cmd_valid = dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 195:72:@159993.4]
  assign io_dram_2_cmd_bits_addr = dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@159992.4]
  assign io_dram_2_cmd_bits_size = dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@159991.4]
  assign io_dram_2_cmd_bits_isWr = dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@159989.4]
  assign io_dram_2_cmd_bits_tag = dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@159988.4]
  assign io_dram_2_wdata_valid = dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 195:72:@159986.4]
  assign io_dram_2_wdata_bits_wdata_0 = dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@159970.4]
  assign io_dram_2_wdata_bits_wdata_1 = dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@159971.4]
  assign io_dram_2_wdata_bits_wdata_2 = dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@159972.4]
  assign io_dram_2_wdata_bits_wdata_3 = dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@159973.4]
  assign io_dram_2_wdata_bits_wdata_4 = dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@159974.4]
  assign io_dram_2_wdata_bits_wdata_5 = dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@159975.4]
  assign io_dram_2_wdata_bits_wdata_6 = dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@159976.4]
  assign io_dram_2_wdata_bits_wdata_7 = dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@159977.4]
  assign io_dram_2_wdata_bits_wdata_8 = dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@159978.4]
  assign io_dram_2_wdata_bits_wdata_9 = dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@159979.4]
  assign io_dram_2_wdata_bits_wdata_10 = dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@159980.4]
  assign io_dram_2_wdata_bits_wdata_11 = dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@159981.4]
  assign io_dram_2_wdata_bits_wdata_12 = dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@159982.4]
  assign io_dram_2_wdata_bits_wdata_13 = dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@159983.4]
  assign io_dram_2_wdata_bits_wdata_14 = dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@159984.4]
  assign io_dram_2_wdata_bits_wdata_15 = dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@159985.4]
  assign io_dram_2_wdata_bits_wstrb_0 = dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@159906.4]
  assign io_dram_2_wdata_bits_wstrb_1 = dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@159907.4]
  assign io_dram_2_wdata_bits_wstrb_2 = dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@159908.4]
  assign io_dram_2_wdata_bits_wstrb_3 = dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@159909.4]
  assign io_dram_2_wdata_bits_wstrb_4 = dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@159910.4]
  assign io_dram_2_wdata_bits_wstrb_5 = dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@159911.4]
  assign io_dram_2_wdata_bits_wstrb_6 = dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@159912.4]
  assign io_dram_2_wdata_bits_wstrb_7 = dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@159913.4]
  assign io_dram_2_wdata_bits_wstrb_8 = dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@159914.4]
  assign io_dram_2_wdata_bits_wstrb_9 = dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@159915.4]
  assign io_dram_2_wdata_bits_wstrb_10 = dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@159916.4]
  assign io_dram_2_wdata_bits_wstrb_11 = dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@159917.4]
  assign io_dram_2_wdata_bits_wstrb_12 = dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@159918.4]
  assign io_dram_2_wdata_bits_wstrb_13 = dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@159919.4]
  assign io_dram_2_wdata_bits_wstrb_14 = dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@159920.4]
  assign io_dram_2_wdata_bits_wstrb_15 = dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@159921.4]
  assign io_dram_2_wdata_bits_wstrb_16 = dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@159922.4]
  assign io_dram_2_wdata_bits_wstrb_17 = dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@159923.4]
  assign io_dram_2_wdata_bits_wstrb_18 = dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@159924.4]
  assign io_dram_2_wdata_bits_wstrb_19 = dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@159925.4]
  assign io_dram_2_wdata_bits_wstrb_20 = dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@159926.4]
  assign io_dram_2_wdata_bits_wstrb_21 = dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@159927.4]
  assign io_dram_2_wdata_bits_wstrb_22 = dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@159928.4]
  assign io_dram_2_wdata_bits_wstrb_23 = dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@159929.4]
  assign io_dram_2_wdata_bits_wstrb_24 = dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@159930.4]
  assign io_dram_2_wdata_bits_wstrb_25 = dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@159931.4]
  assign io_dram_2_wdata_bits_wstrb_26 = dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@159932.4]
  assign io_dram_2_wdata_bits_wstrb_27 = dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@159933.4]
  assign io_dram_2_wdata_bits_wstrb_28 = dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@159934.4]
  assign io_dram_2_wdata_bits_wstrb_29 = dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@159935.4]
  assign io_dram_2_wdata_bits_wstrb_30 = dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@159936.4]
  assign io_dram_2_wdata_bits_wstrb_31 = dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@159937.4]
  assign io_dram_2_wdata_bits_wstrb_32 = dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@159938.4]
  assign io_dram_2_wdata_bits_wstrb_33 = dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@159939.4]
  assign io_dram_2_wdata_bits_wstrb_34 = dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@159940.4]
  assign io_dram_2_wdata_bits_wstrb_35 = dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@159941.4]
  assign io_dram_2_wdata_bits_wstrb_36 = dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@159942.4]
  assign io_dram_2_wdata_bits_wstrb_37 = dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@159943.4]
  assign io_dram_2_wdata_bits_wstrb_38 = dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@159944.4]
  assign io_dram_2_wdata_bits_wstrb_39 = dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@159945.4]
  assign io_dram_2_wdata_bits_wstrb_40 = dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@159946.4]
  assign io_dram_2_wdata_bits_wstrb_41 = dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@159947.4]
  assign io_dram_2_wdata_bits_wstrb_42 = dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@159948.4]
  assign io_dram_2_wdata_bits_wstrb_43 = dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@159949.4]
  assign io_dram_2_wdata_bits_wstrb_44 = dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@159950.4]
  assign io_dram_2_wdata_bits_wstrb_45 = dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@159951.4]
  assign io_dram_2_wdata_bits_wstrb_46 = dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@159952.4]
  assign io_dram_2_wdata_bits_wstrb_47 = dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@159953.4]
  assign io_dram_2_wdata_bits_wstrb_48 = dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@159954.4]
  assign io_dram_2_wdata_bits_wstrb_49 = dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@159955.4]
  assign io_dram_2_wdata_bits_wstrb_50 = dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@159956.4]
  assign io_dram_2_wdata_bits_wstrb_51 = dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@159957.4]
  assign io_dram_2_wdata_bits_wstrb_52 = dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@159958.4]
  assign io_dram_2_wdata_bits_wstrb_53 = dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@159959.4]
  assign io_dram_2_wdata_bits_wstrb_54 = dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@159960.4]
  assign io_dram_2_wdata_bits_wstrb_55 = dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@159961.4]
  assign io_dram_2_wdata_bits_wstrb_56 = dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@159962.4]
  assign io_dram_2_wdata_bits_wstrb_57 = dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@159963.4]
  assign io_dram_2_wdata_bits_wstrb_58 = dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@159964.4]
  assign io_dram_2_wdata_bits_wstrb_59 = dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@159965.4]
  assign io_dram_2_wdata_bits_wstrb_60 = dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@159966.4]
  assign io_dram_2_wdata_bits_wstrb_61 = dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@159967.4]
  assign io_dram_2_wdata_bits_wstrb_62 = dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@159968.4]
  assign io_dram_2_wdata_bits_wstrb_63 = dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@159969.4]
  assign io_dram_2_wdata_bits_wlast = dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@159905.4]
  assign io_dram_2_rresp_ready = dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 195:72:@159904.4]
  assign io_dram_2_wresp_ready = dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 195:72:@159885.4]
  assign io_dram_3_cmd_valid = dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 195:72:@160105.4]
  assign io_dram_3_cmd_bits_addr = dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@160104.4]
  assign io_dram_3_cmd_bits_size = dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@160103.4]
  assign io_dram_3_cmd_bits_isWr = dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@160101.4]
  assign io_dram_3_cmd_bits_tag = dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@160100.4]
  assign io_dram_3_wdata_valid = dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 195:72:@160098.4]
  assign io_dram_3_wdata_bits_wdata_0 = dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@160082.4]
  assign io_dram_3_wdata_bits_wdata_1 = dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@160083.4]
  assign io_dram_3_wdata_bits_wdata_2 = dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@160084.4]
  assign io_dram_3_wdata_bits_wdata_3 = dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@160085.4]
  assign io_dram_3_wdata_bits_wdata_4 = dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@160086.4]
  assign io_dram_3_wdata_bits_wdata_5 = dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@160087.4]
  assign io_dram_3_wdata_bits_wdata_6 = dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@160088.4]
  assign io_dram_3_wdata_bits_wdata_7 = dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@160089.4]
  assign io_dram_3_wdata_bits_wdata_8 = dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@160090.4]
  assign io_dram_3_wdata_bits_wdata_9 = dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@160091.4]
  assign io_dram_3_wdata_bits_wdata_10 = dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@160092.4]
  assign io_dram_3_wdata_bits_wdata_11 = dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@160093.4]
  assign io_dram_3_wdata_bits_wdata_12 = dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@160094.4]
  assign io_dram_3_wdata_bits_wdata_13 = dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@160095.4]
  assign io_dram_3_wdata_bits_wdata_14 = dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@160096.4]
  assign io_dram_3_wdata_bits_wdata_15 = dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@160097.4]
  assign io_dram_3_wdata_bits_wstrb_0 = dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@160018.4]
  assign io_dram_3_wdata_bits_wstrb_1 = dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@160019.4]
  assign io_dram_3_wdata_bits_wstrb_2 = dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@160020.4]
  assign io_dram_3_wdata_bits_wstrb_3 = dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@160021.4]
  assign io_dram_3_wdata_bits_wstrb_4 = dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@160022.4]
  assign io_dram_3_wdata_bits_wstrb_5 = dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@160023.4]
  assign io_dram_3_wdata_bits_wstrb_6 = dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@160024.4]
  assign io_dram_3_wdata_bits_wstrb_7 = dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@160025.4]
  assign io_dram_3_wdata_bits_wstrb_8 = dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@160026.4]
  assign io_dram_3_wdata_bits_wstrb_9 = dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@160027.4]
  assign io_dram_3_wdata_bits_wstrb_10 = dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@160028.4]
  assign io_dram_3_wdata_bits_wstrb_11 = dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@160029.4]
  assign io_dram_3_wdata_bits_wstrb_12 = dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@160030.4]
  assign io_dram_3_wdata_bits_wstrb_13 = dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@160031.4]
  assign io_dram_3_wdata_bits_wstrb_14 = dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@160032.4]
  assign io_dram_3_wdata_bits_wstrb_15 = dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@160033.4]
  assign io_dram_3_wdata_bits_wstrb_16 = dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@160034.4]
  assign io_dram_3_wdata_bits_wstrb_17 = dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@160035.4]
  assign io_dram_3_wdata_bits_wstrb_18 = dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@160036.4]
  assign io_dram_3_wdata_bits_wstrb_19 = dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@160037.4]
  assign io_dram_3_wdata_bits_wstrb_20 = dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@160038.4]
  assign io_dram_3_wdata_bits_wstrb_21 = dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@160039.4]
  assign io_dram_3_wdata_bits_wstrb_22 = dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@160040.4]
  assign io_dram_3_wdata_bits_wstrb_23 = dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@160041.4]
  assign io_dram_3_wdata_bits_wstrb_24 = dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@160042.4]
  assign io_dram_3_wdata_bits_wstrb_25 = dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@160043.4]
  assign io_dram_3_wdata_bits_wstrb_26 = dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@160044.4]
  assign io_dram_3_wdata_bits_wstrb_27 = dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@160045.4]
  assign io_dram_3_wdata_bits_wstrb_28 = dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@160046.4]
  assign io_dram_3_wdata_bits_wstrb_29 = dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@160047.4]
  assign io_dram_3_wdata_bits_wstrb_30 = dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@160048.4]
  assign io_dram_3_wdata_bits_wstrb_31 = dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@160049.4]
  assign io_dram_3_wdata_bits_wstrb_32 = dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@160050.4]
  assign io_dram_3_wdata_bits_wstrb_33 = dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@160051.4]
  assign io_dram_3_wdata_bits_wstrb_34 = dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@160052.4]
  assign io_dram_3_wdata_bits_wstrb_35 = dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@160053.4]
  assign io_dram_3_wdata_bits_wstrb_36 = dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@160054.4]
  assign io_dram_3_wdata_bits_wstrb_37 = dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@160055.4]
  assign io_dram_3_wdata_bits_wstrb_38 = dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@160056.4]
  assign io_dram_3_wdata_bits_wstrb_39 = dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@160057.4]
  assign io_dram_3_wdata_bits_wstrb_40 = dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@160058.4]
  assign io_dram_3_wdata_bits_wstrb_41 = dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@160059.4]
  assign io_dram_3_wdata_bits_wstrb_42 = dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@160060.4]
  assign io_dram_3_wdata_bits_wstrb_43 = dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@160061.4]
  assign io_dram_3_wdata_bits_wstrb_44 = dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@160062.4]
  assign io_dram_3_wdata_bits_wstrb_45 = dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@160063.4]
  assign io_dram_3_wdata_bits_wstrb_46 = dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@160064.4]
  assign io_dram_3_wdata_bits_wstrb_47 = dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@160065.4]
  assign io_dram_3_wdata_bits_wstrb_48 = dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@160066.4]
  assign io_dram_3_wdata_bits_wstrb_49 = dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@160067.4]
  assign io_dram_3_wdata_bits_wstrb_50 = dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@160068.4]
  assign io_dram_3_wdata_bits_wstrb_51 = dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@160069.4]
  assign io_dram_3_wdata_bits_wstrb_52 = dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@160070.4]
  assign io_dram_3_wdata_bits_wstrb_53 = dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@160071.4]
  assign io_dram_3_wdata_bits_wstrb_54 = dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@160072.4]
  assign io_dram_3_wdata_bits_wstrb_55 = dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@160073.4]
  assign io_dram_3_wdata_bits_wstrb_56 = dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@160074.4]
  assign io_dram_3_wdata_bits_wstrb_57 = dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@160075.4]
  assign io_dram_3_wdata_bits_wstrb_58 = dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@160076.4]
  assign io_dram_3_wdata_bits_wstrb_59 = dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@160077.4]
  assign io_dram_3_wdata_bits_wstrb_60 = dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@160078.4]
  assign io_dram_3_wdata_bits_wstrb_61 = dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@160079.4]
  assign io_dram_3_wdata_bits_wstrb_62 = dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@160080.4]
  assign io_dram_3_wdata_bits_wstrb_63 = dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@160081.4]
  assign io_dram_3_wdata_bits_wlast = dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@160017.4]
  assign io_dram_3_rresp_ready = dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 195:72:@160016.4]
  assign io_dram_3_wresp_ready = dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 195:72:@159997.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@156536.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@156535.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@156534.4]
  assign dramArbs_0_clock = clock; // @[:@152659.4]
  assign dramArbs_0_reset = _T_1030 | reset; // @[:@152660.4 Fringe.scala 187:30:@159651.4]
  assign dramArbs_0_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@159655.4]
  assign dramArbs_0_io_app_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[Fringe.scala 101:72:@153576.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[Fringe.scala 101:72:@153575.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[Fringe.scala 101:72:@153574.4]
  assign dramArbs_0_io_app_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[Fringe.scala 101:72:@153572.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[Fringe.scala 101:72:@153571.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[Fringe.scala 101:72:@153570.4]
  assign dramArbs_0_io_app_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[Fringe.scala 101:72:@153569.4]
  assign dramArbs_0_io_dram_cmd_ready = io_dram_0_cmd_ready; // @[Fringe.scala 195:72:@159770.4]
  assign dramArbs_0_io_dram_wdata_ready = io_dram_0_wdata_ready; // @[Fringe.scala 195:72:@159763.4]
  assign dramArbs_0_io_dram_wresp_valid = io_dram_0_wresp_valid; // @[Fringe.scala 195:72:@159660.4]
  assign dramArbs_0_io_dram_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[Fringe.scala 195:72:@159659.4]
  assign dramArbs_1_clock = clock; // @[:@153652.4]
  assign dramArbs_1_reset = _T_1030 | reset; // @[:@153653.4 Fringe.scala 187:30:@159652.4]
  assign dramArbs_1_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@159656.4]
  assign dramArbs_1_io_dram_cmd_ready = io_dram_1_cmd_ready; // @[Fringe.scala 195:72:@159882.4]
  assign dramArbs_1_io_dram_wdata_ready = io_dram_1_wdata_ready; // @[Fringe.scala 195:72:@159875.4]
  assign dramArbs_1_io_dram_wresp_valid = io_dram_1_wresp_valid; // @[Fringe.scala 195:72:@159772.4]
  assign dramArbs_1_io_dram_wresp_bits_tag = io_dram_1_wresp_bits_tag; // @[Fringe.scala 195:72:@159771.4]
  assign dramArbs_2_clock = clock; // @[:@154612.4]
  assign dramArbs_2_reset = _T_1030 | reset; // @[:@154613.4 Fringe.scala 187:30:@159653.4]
  assign dramArbs_2_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@159657.4]
  assign dramArbs_2_io_dram_cmd_ready = io_dram_2_cmd_ready; // @[Fringe.scala 195:72:@159994.4]
  assign dramArbs_2_io_dram_wdata_ready = io_dram_2_wdata_ready; // @[Fringe.scala 195:72:@159987.4]
  assign dramArbs_2_io_dram_wresp_valid = io_dram_2_wresp_valid; // @[Fringe.scala 195:72:@159884.4]
  assign dramArbs_2_io_dram_wresp_bits_tag = io_dram_2_wresp_bits_tag; // @[Fringe.scala 195:72:@159883.4]
  assign dramArbs_3_clock = clock; // @[:@155572.4]
  assign dramArbs_3_reset = _T_1030 | reset; // @[:@155573.4 Fringe.scala 187:30:@159654.4]
  assign dramArbs_3_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@159658.4]
  assign dramArbs_3_io_dram_cmd_ready = io_dram_3_cmd_ready; // @[Fringe.scala 195:72:@160106.4]
  assign dramArbs_3_io_dram_wdata_ready = io_dram_3_wdata_ready; // @[Fringe.scala 195:72:@160099.4]
  assign dramArbs_3_io_dram_wresp_valid = io_dram_3_wresp_valid; // @[Fringe.scala 195:72:@159996.4]
  assign dramArbs_3_io_dram_wresp_bits_tag = io_dram_3_wresp_bits_tag; // @[Fringe.scala 195:72:@159995.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@156539.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@156538.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@156537.4]
  assign heap_io_host_0_resp_valid = _T_1569 & _T_1573; // @[Fringe.scala 204:22:@160278.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@160279.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@160280.4]
  assign regs_clock = clock; // @[:@156541.4]
  assign regs_reset = reset; // @[:@156542.4 Fringe.scala 139:14:@158589.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@158561.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@158563.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@158562.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@158564.4]
  assign regs_io_reset = _T_1030 | reset; // @[Fringe.scala 138:17:@158587.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_1049; // @[Fringe.scala 170:23:@158639.4]
  assign regs_io_argOuts_0_bits = {_T_1065,_T_1064}; // @[Fringe.scala 171:22:@158643.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@158646.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@158645.4]
  assign timeoutCtr_clock = clock; // @[:@158591.4]
  assign timeoutCtr_reset = reset; // @[:@158592.4]
  assign timeoutCtr_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 149:24:@158606.4]
  assign depulser_clock = clock; // @[:@158610.4]
  assign depulser_reset = reset; // @[:@158611.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@158616.4]
  assign depulser_io_rst = _T_1040[0]; // @[Fringe.scala 156:19:@158618.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1047 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1572 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1047 <= 1'h0;
    end else begin
      _T_1047 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1572 <= 1'h0;
    end else begin
      _T_1572 <= _T_1569;
    end
  end
endmodule
module AXI4LiteToRFBridge( // @[:@160295.2]
  input         clock, // @[:@160296.4]
  input         reset, // @[:@160297.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@160298.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@160298.4]
  input         io_S_AXI_AWVALID, // @[:@160298.4]
  output        io_S_AXI_AWREADY, // @[:@160298.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@160298.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@160298.4]
  input         io_S_AXI_ARVALID, // @[:@160298.4]
  output        io_S_AXI_ARREADY, // @[:@160298.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@160298.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@160298.4]
  input         io_S_AXI_WVALID, // @[:@160298.4]
  output        io_S_AXI_WREADY, // @[:@160298.4]
  output [31:0] io_S_AXI_RDATA, // @[:@160298.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@160298.4]
  output        io_S_AXI_RVALID, // @[:@160298.4]
  input         io_S_AXI_RREADY, // @[:@160298.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@160298.4]
  output        io_S_AXI_BVALID, // @[:@160298.4]
  input         io_S_AXI_BREADY, // @[:@160298.4]
  output [31:0] io_raddr, // @[:@160298.4]
  output        io_wen, // @[:@160298.4]
  output [31:0] io_waddr, // @[:@160298.4]
  output [31:0] io_wdata, // @[:@160298.4]
  input  [31:0] io_rdata // @[:@160298.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 36:17:@160300.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 38:14:@160324.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 38:14:@160320.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 38:14:@160316.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 38:14:@160315.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 38:14:@160314.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 38:14:@160313.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 38:14:@160311.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 38:14:@160310.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 42:12:@160332.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 45:12:@160335.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 43:12:@160333.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 44:12:@160334.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 46:17:@160336.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 40:22:@160331.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 39:19:@160328.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 38:14:@160327.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 38:14:@160326.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 38:14:@160325.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 38:14:@160323.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 38:14:@160322.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 38:14:@160321.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 38:14:@160319.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 38:14:@160318.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 38:14:@160317.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 38:14:@160312.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 38:14:@160309.4]
endmodule
module MAGToAXI4Bridge( // @[:@160338.2]
  output         io_in_cmd_ready, // @[:@160341.4]
  input          io_in_cmd_valid, // @[:@160341.4]
  input  [63:0]  io_in_cmd_bits_addr, // @[:@160341.4]
  input  [31:0]  io_in_cmd_bits_size, // @[:@160341.4]
  input          io_in_cmd_bits_isWr, // @[:@160341.4]
  input  [31:0]  io_in_cmd_bits_tag, // @[:@160341.4]
  output         io_in_wdata_ready, // @[:@160341.4]
  input          io_in_wdata_valid, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_0, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_1, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_2, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_3, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_4, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_5, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_6, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_7, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_8, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_9, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_10, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_11, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_12, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_13, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_14, // @[:@160341.4]
  input  [31:0]  io_in_wdata_bits_wdata_15, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_0, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_1, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_2, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_3, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_4, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_5, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_6, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_7, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_8, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_9, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_10, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_11, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_12, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_13, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_14, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_15, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_16, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_17, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_18, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_19, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_20, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_21, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_22, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_23, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_24, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_25, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_26, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_27, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_28, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_29, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_30, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_31, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_32, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_33, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_34, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_35, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_36, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_37, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_38, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_39, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_40, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_41, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_42, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_43, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_44, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_45, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_46, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_47, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_48, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_49, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_50, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_51, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_52, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_53, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_54, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_55, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_56, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_57, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_58, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_59, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_60, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_61, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_62, // @[:@160341.4]
  input          io_in_wdata_bits_wstrb_63, // @[:@160341.4]
  input          io_in_wdata_bits_wlast, // @[:@160341.4]
  input          io_in_rresp_ready, // @[:@160341.4]
  input          io_in_wresp_ready, // @[:@160341.4]
  output         io_in_wresp_valid, // @[:@160341.4]
  output [31:0]  io_in_wresp_bits_tag, // @[:@160341.4]
  output [31:0]  io_M_AXI_AWID, // @[:@160341.4]
  output [31:0]  io_M_AXI_AWADDR, // @[:@160341.4]
  output [7:0]   io_M_AXI_AWLEN, // @[:@160341.4]
  output         io_M_AXI_AWVALID, // @[:@160341.4]
  input          io_M_AXI_AWREADY, // @[:@160341.4]
  output [31:0]  io_M_AXI_ARID, // @[:@160341.4]
  output [31:0]  io_M_AXI_ARADDR, // @[:@160341.4]
  output [7:0]   io_M_AXI_ARLEN, // @[:@160341.4]
  output         io_M_AXI_ARVALID, // @[:@160341.4]
  input          io_M_AXI_ARREADY, // @[:@160341.4]
  output [511:0] io_M_AXI_WDATA, // @[:@160341.4]
  output [63:0]  io_M_AXI_WSTRB, // @[:@160341.4]
  output         io_M_AXI_WLAST, // @[:@160341.4]
  output         io_M_AXI_WVALID, // @[:@160341.4]
  input          io_M_AXI_WREADY, // @[:@160341.4]
  output         io_M_AXI_RREADY, // @[:@160341.4]
  input  [31:0]  io_M_AXI_BID, // @[:@160341.4]
  input          io_M_AXI_BVALID, // @[:@160341.4]
  output         io_M_AXI_BREADY // @[:@160341.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@160498.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@160499.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@160500.4]
  wire  _T_228; // @[MAGToAXI4Bridge.scala 35:42:@160508.4]
  wire [319:0] _T_250; // @[Cat.scala 30:58:@160535.4]
  wire [479:0] _T_255; // @[Cat.scala 30:58:@160540.4]
  wire [9:0] _T_265; // @[Cat.scala 30:58:@160551.4]
  wire [18:0] _T_274; // @[Cat.scala 30:58:@160560.4]
  wire [27:0] _T_283; // @[Cat.scala 30:58:@160569.4]
  wire [36:0] _T_292; // @[Cat.scala 30:58:@160578.4]
  wire [45:0] _T_301; // @[Cat.scala 30:58:@160587.4]
  wire [54:0] _T_310; // @[Cat.scala 30:58:@160596.4]
  wire [62:0] _T_318; // @[Cat.scala 30:58:@160604.4]
  assign _T_218 = io_in_cmd_bits_size - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@160498.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@160499.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@160500.4]
  assign _T_228 = io_in_cmd_bits_isWr == 1'h0; // @[MAGToAXI4Bridge.scala 35:42:@160508.4]
  assign _T_250 = {io_in_wdata_bits_wdata_15,io_in_wdata_bits_wdata_14,io_in_wdata_bits_wdata_13,io_in_wdata_bits_wdata_12,io_in_wdata_bits_wdata_11,io_in_wdata_bits_wdata_10,io_in_wdata_bits_wdata_9,io_in_wdata_bits_wdata_8,io_in_wdata_bits_wdata_7,io_in_wdata_bits_wdata_6}; // @[Cat.scala 30:58:@160535.4]
  assign _T_255 = {_T_250,io_in_wdata_bits_wdata_5,io_in_wdata_bits_wdata_4,io_in_wdata_bits_wdata_3,io_in_wdata_bits_wdata_2,io_in_wdata_bits_wdata_1}; // @[Cat.scala 30:58:@160540.4]
  assign _T_265 = {io_in_wdata_bits_wstrb_63,io_in_wdata_bits_wstrb_62,io_in_wdata_bits_wstrb_61,io_in_wdata_bits_wstrb_60,io_in_wdata_bits_wstrb_59,io_in_wdata_bits_wstrb_58,io_in_wdata_bits_wstrb_57,io_in_wdata_bits_wstrb_56,io_in_wdata_bits_wstrb_55,io_in_wdata_bits_wstrb_54}; // @[Cat.scala 30:58:@160551.4]
  assign _T_274 = {_T_265,io_in_wdata_bits_wstrb_53,io_in_wdata_bits_wstrb_52,io_in_wdata_bits_wstrb_51,io_in_wdata_bits_wstrb_50,io_in_wdata_bits_wstrb_49,io_in_wdata_bits_wstrb_48,io_in_wdata_bits_wstrb_47,io_in_wdata_bits_wstrb_46,io_in_wdata_bits_wstrb_45}; // @[Cat.scala 30:58:@160560.4]
  assign _T_283 = {_T_274,io_in_wdata_bits_wstrb_44,io_in_wdata_bits_wstrb_43,io_in_wdata_bits_wstrb_42,io_in_wdata_bits_wstrb_41,io_in_wdata_bits_wstrb_40,io_in_wdata_bits_wstrb_39,io_in_wdata_bits_wstrb_38,io_in_wdata_bits_wstrb_37,io_in_wdata_bits_wstrb_36}; // @[Cat.scala 30:58:@160569.4]
  assign _T_292 = {_T_283,io_in_wdata_bits_wstrb_35,io_in_wdata_bits_wstrb_34,io_in_wdata_bits_wstrb_33,io_in_wdata_bits_wstrb_32,io_in_wdata_bits_wstrb_31,io_in_wdata_bits_wstrb_30,io_in_wdata_bits_wstrb_29,io_in_wdata_bits_wstrb_28,io_in_wdata_bits_wstrb_27}; // @[Cat.scala 30:58:@160578.4]
  assign _T_301 = {_T_292,io_in_wdata_bits_wstrb_26,io_in_wdata_bits_wstrb_25,io_in_wdata_bits_wstrb_24,io_in_wdata_bits_wstrb_23,io_in_wdata_bits_wstrb_22,io_in_wdata_bits_wstrb_21,io_in_wdata_bits_wstrb_20,io_in_wdata_bits_wstrb_19,io_in_wdata_bits_wstrb_18}; // @[Cat.scala 30:58:@160587.4]
  assign _T_310 = {_T_301,io_in_wdata_bits_wstrb_17,io_in_wdata_bits_wstrb_16,io_in_wdata_bits_wstrb_15,io_in_wdata_bits_wstrb_14,io_in_wdata_bits_wstrb_13,io_in_wdata_bits_wstrb_12,io_in_wdata_bits_wstrb_11,io_in_wdata_bits_wstrb_10,io_in_wdata_bits_wstrb_9}; // @[Cat.scala 30:58:@160596.4]
  assign _T_318 = {_T_310,io_in_wdata_bits_wstrb_8,io_in_wdata_bits_wstrb_7,io_in_wdata_bits_wstrb_6,io_in_wdata_bits_wstrb_5,io_in_wdata_bits_wstrb_4,io_in_wdata_bits_wstrb_3,io_in_wdata_bits_wstrb_2,io_in_wdata_bits_wstrb_1}; // @[Cat.scala 30:58:@160604.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? io_M_AXI_AWREADY : io_M_AXI_ARREADY; // @[MAGToAXI4Bridge.scala 36:21:@160512.4]
  assign io_in_wdata_ready = io_M_AXI_WREADY; // @[MAGToAXI4Bridge.scala 56:21:@160609.4]
  assign io_in_wresp_valid = io_M_AXI_BVALID; // @[MAGToAXI4Bridge.scala 71:21:@160662.4]
  assign io_in_wresp_bits_tag = io_M_AXI_BID; // @[MAGToAXI4Bridge.scala 74:24:@160664.4]
  assign io_M_AXI_AWID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 39:21:@160513.4]
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 40:21:@160514.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@160518.4]
  assign io_M_AXI_AWVALID = io_in_cmd_valid & io_in_cmd_bits_isWr; // @[MAGToAXI4Bridge.scala 49:21:@160526.4]
  assign io_M_AXI_ARID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 25:21:@160496.4]
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 26:21:@160497.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@160501.4]
  assign io_M_AXI_ARVALID = io_in_cmd_valid & _T_228; // @[MAGToAXI4Bridge.scala 35:21:@160510.4]
  assign io_M_AXI_WDATA = {_T_255,io_in_wdata_bits_wdata_0}; // @[MAGToAXI4Bridge.scala 52:21:@160542.4]
  assign io_M_AXI_WSTRB = {_T_318,io_in_wdata_bits_wstrb_0}; // @[MAGToAXI4Bridge.scala 53:21:@160606.4]
  assign io_M_AXI_WLAST = io_in_wdata_bits_wlast; // @[MAGToAXI4Bridge.scala 54:21:@160607.4]
  assign io_M_AXI_WVALID = io_in_wdata_valid; // @[MAGToAXI4Bridge.scala 55:21:@160608.4]
  assign io_M_AXI_RREADY = io_in_rresp_ready; // @[MAGToAXI4Bridge.scala 64:19:@160659.4]
  assign io_M_AXI_BREADY = io_in_wresp_ready; // @[MAGToAXI4Bridge.scala 67:19:@160660.4]
endmodule
module FringeZynq( // @[:@161650.2]
  input          clock, // @[:@161651.4]
  input          reset, // @[:@161652.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@161653.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@161653.4]
  input          io_S_AXI_AWVALID, // @[:@161653.4]
  output         io_S_AXI_AWREADY, // @[:@161653.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@161653.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@161653.4]
  input          io_S_AXI_ARVALID, // @[:@161653.4]
  output         io_S_AXI_ARREADY, // @[:@161653.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@161653.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@161653.4]
  input          io_S_AXI_WVALID, // @[:@161653.4]
  output         io_S_AXI_WREADY, // @[:@161653.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@161653.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@161653.4]
  output         io_S_AXI_RVALID, // @[:@161653.4]
  input          io_S_AXI_RREADY, // @[:@161653.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@161653.4]
  output         io_S_AXI_BVALID, // @[:@161653.4]
  input          io_S_AXI_BREADY, // @[:@161653.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@161653.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@161653.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@161653.4]
  output         io_M_AXI_0_AWVALID, // @[:@161653.4]
  input          io_M_AXI_0_AWREADY, // @[:@161653.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@161653.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@161653.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@161653.4]
  output         io_M_AXI_0_ARVALID, // @[:@161653.4]
  input          io_M_AXI_0_ARREADY, // @[:@161653.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@161653.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@161653.4]
  output         io_M_AXI_0_WLAST, // @[:@161653.4]
  output         io_M_AXI_0_WVALID, // @[:@161653.4]
  input          io_M_AXI_0_WREADY, // @[:@161653.4]
  output         io_M_AXI_0_RREADY, // @[:@161653.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@161653.4]
  input          io_M_AXI_0_BVALID, // @[:@161653.4]
  output         io_M_AXI_0_BREADY, // @[:@161653.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@161653.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@161653.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@161653.4]
  output         io_M_AXI_1_AWVALID, // @[:@161653.4]
  input          io_M_AXI_1_AWREADY, // @[:@161653.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@161653.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@161653.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@161653.4]
  output         io_M_AXI_1_ARVALID, // @[:@161653.4]
  input          io_M_AXI_1_ARREADY, // @[:@161653.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@161653.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@161653.4]
  output         io_M_AXI_1_WLAST, // @[:@161653.4]
  output         io_M_AXI_1_WVALID, // @[:@161653.4]
  input          io_M_AXI_1_WREADY, // @[:@161653.4]
  output         io_M_AXI_1_RREADY, // @[:@161653.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@161653.4]
  input          io_M_AXI_1_BVALID, // @[:@161653.4]
  output         io_M_AXI_1_BREADY, // @[:@161653.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@161653.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@161653.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@161653.4]
  output         io_M_AXI_2_AWVALID, // @[:@161653.4]
  input          io_M_AXI_2_AWREADY, // @[:@161653.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@161653.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@161653.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@161653.4]
  output         io_M_AXI_2_ARVALID, // @[:@161653.4]
  input          io_M_AXI_2_ARREADY, // @[:@161653.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@161653.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@161653.4]
  output         io_M_AXI_2_WLAST, // @[:@161653.4]
  output         io_M_AXI_2_WVALID, // @[:@161653.4]
  input          io_M_AXI_2_WREADY, // @[:@161653.4]
  output         io_M_AXI_2_RREADY, // @[:@161653.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@161653.4]
  input          io_M_AXI_2_BVALID, // @[:@161653.4]
  output         io_M_AXI_2_BREADY, // @[:@161653.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@161653.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@161653.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@161653.4]
  output         io_M_AXI_3_AWVALID, // @[:@161653.4]
  input          io_M_AXI_3_AWREADY, // @[:@161653.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@161653.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@161653.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@161653.4]
  output         io_M_AXI_3_ARVALID, // @[:@161653.4]
  input          io_M_AXI_3_ARREADY, // @[:@161653.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@161653.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@161653.4]
  output         io_M_AXI_3_WLAST, // @[:@161653.4]
  output         io_M_AXI_3_WVALID, // @[:@161653.4]
  input          io_M_AXI_3_WREADY, // @[:@161653.4]
  output         io_M_AXI_3_RREADY, // @[:@161653.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@161653.4]
  input          io_M_AXI_3_BVALID, // @[:@161653.4]
  output         io_M_AXI_3_BREADY, // @[:@161653.4]
  output         io_enable, // @[:@161653.4]
  input          io_done, // @[:@161653.4]
  output         io_reset, // @[:@161653.4]
  output [63:0]  io_argIns_0, // @[:@161653.4]
  output [63:0]  io_argIns_1, // @[:@161653.4]
  input          io_argOuts_0_valid, // @[:@161653.4]
  input  [63:0]  io_argOuts_0_bits, // @[:@161653.4]
  output         io_memStreams_stores_0_cmd_ready, // @[:@161653.4]
  input          io_memStreams_stores_0_cmd_valid, // @[:@161653.4]
  input  [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@161653.4]
  input  [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@161653.4]
  output         io_memStreams_stores_0_data_ready, // @[:@161653.4]
  input          io_memStreams_stores_0_data_valid, // @[:@161653.4]
  input  [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@161653.4]
  input          io_memStreams_stores_0_data_bits_wstrb, // @[:@161653.4]
  input          io_memStreams_stores_0_wresp_ready, // @[:@161653.4]
  output         io_memStreams_stores_0_wresp_valid, // @[:@161653.4]
  output         io_memStreams_stores_0_wresp_bits, // @[:@161653.4]
  input          io_heap_0_req_valid, // @[:@161653.4]
  input          io_heap_0_req_bits_allocDealloc, // @[:@161653.4]
  input  [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@161653.4]
  output         io_heap_0_resp_valid, // @[:@161653.4]
  output         io_heap_0_resp_bits_allocDealloc, // @[:@161653.4]
  output [63:0]  io_heap_0_resp_bits_sizeAddr // @[:@161653.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 69:28:@162124.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 69:28:@162124.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 69:28:@162124.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 69:28:@162124.4]
  wire [63:0] fringeCommon_io_argIns_1; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire [63:0] fringeCommon_io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_cmd_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_0_wresp_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_0_wresp_bits_tag; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_cmd_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire [63:0] fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_1_wresp_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_1_wresp_bits_tag; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_cmd_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire [63:0] fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_2_wresp_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_2_wresp_bits_tag; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_cmd_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire [63:0] fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_dram_3_wresp_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire [31:0] fringeCommon_io_dram_3_wresp_bits_tag; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 69:28:@162124.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 69:28:@162124.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 69:28:@162124.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 69:28:@162124.4]
  wire  AXI4LiteToRFBridge_clock; // @[FringeZynq.scala 90:31:@163030.4]
  wire  AXI4LiteToRFBridge_reset; // @[FringeZynq.scala 90:31:@163030.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_AWADDR; // @[FringeZynq.scala 90:31:@163030.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_AWPROT; // @[FringeZynq.scala 90:31:@163030.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWVALID; // @[FringeZynq.scala 90:31:@163030.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 90:31:@163030.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_ARADDR; // @[FringeZynq.scala 90:31:@163030.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_ARPROT; // @[FringeZynq.scala 90:31:@163030.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARVALID; // @[FringeZynq.scala 90:31:@163030.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 90:31:@163030.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_WDATA; // @[FringeZynq.scala 90:31:@163030.4]
  wire [3:0] AXI4LiteToRFBridge_io_S_AXI_WSTRB; // @[FringeZynq.scala 90:31:@163030.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WVALID; // @[FringeZynq.scala 90:31:@163030.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 90:31:@163030.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 90:31:@163030.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 90:31:@163030.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 90:31:@163030.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RREADY; // @[FringeZynq.scala 90:31:@163030.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 90:31:@163030.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 90:31:@163030.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BREADY; // @[FringeZynq.scala 90:31:@163030.4]
  wire [31:0] AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 90:31:@163030.4]
  wire  AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 90:31:@163030.4]
  wire [31:0] AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 90:31:@163030.4]
  wire [31:0] AXI4LiteToRFBridge_io_wdata; // @[FringeZynq.scala 90:31:@163030.4]
  wire [31:0] AXI4LiteToRFBridge_io_rdata; // @[FringeZynq.scala 90:31:@163030.4]
  wire  MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@163180.4]
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@163180.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@163180.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@163180.4]
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@163180.4]
  wire [63:0] MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@163180.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@163180.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@163336.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@163336.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@163336.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@163336.4]
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@163336.4]
  wire [63:0] MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@163336.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@163336.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@163492.4]
  wire [63:0] MAGToAXI4Bridge_2_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@163492.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@163492.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@163492.4]
  wire [511:0] MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@163492.4]
  wire [63:0] MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@163492.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@163492.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@163648.4]
  wire [63:0] MAGToAXI4Bridge_3_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@163648.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@163648.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@163648.4]
  wire [511:0] MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@163648.4]
  wire [63:0] MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@163648.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@163648.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@163648.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 69:28:@162124.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argIns_1(fringeCommon_io_argIns_1),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(fringeCommon_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(fringeCommon_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(fringeCommon_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(fringeCommon_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(fringeCommon_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(fringeCommon_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(fringeCommon_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(fringeCommon_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(fringeCommon_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(fringeCommon_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(fringeCommon_io_memStreams_stores_0_wresp_bits),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_isWr(fringeCommon_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag(fringeCommon_io_dram_0_cmd_bits_tag),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(fringeCommon_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(fringeCommon_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(fringeCommon_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(fringeCommon_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(fringeCommon_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(fringeCommon_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(fringeCommon_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(fringeCommon_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(fringeCommon_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wdata_8(fringeCommon_io_dram_0_wdata_bits_wdata_8),
    .io_dram_0_wdata_bits_wdata_9(fringeCommon_io_dram_0_wdata_bits_wdata_9),
    .io_dram_0_wdata_bits_wdata_10(fringeCommon_io_dram_0_wdata_bits_wdata_10),
    .io_dram_0_wdata_bits_wdata_11(fringeCommon_io_dram_0_wdata_bits_wdata_11),
    .io_dram_0_wdata_bits_wdata_12(fringeCommon_io_dram_0_wdata_bits_wdata_12),
    .io_dram_0_wdata_bits_wdata_13(fringeCommon_io_dram_0_wdata_bits_wdata_13),
    .io_dram_0_wdata_bits_wdata_14(fringeCommon_io_dram_0_wdata_bits_wdata_14),
    .io_dram_0_wdata_bits_wdata_15(fringeCommon_io_dram_0_wdata_bits_wdata_15),
    .io_dram_0_wdata_bits_wstrb_0(fringeCommon_io_dram_0_wdata_bits_wstrb_0),
    .io_dram_0_wdata_bits_wstrb_1(fringeCommon_io_dram_0_wdata_bits_wstrb_1),
    .io_dram_0_wdata_bits_wstrb_2(fringeCommon_io_dram_0_wdata_bits_wstrb_2),
    .io_dram_0_wdata_bits_wstrb_3(fringeCommon_io_dram_0_wdata_bits_wstrb_3),
    .io_dram_0_wdata_bits_wstrb_4(fringeCommon_io_dram_0_wdata_bits_wstrb_4),
    .io_dram_0_wdata_bits_wstrb_5(fringeCommon_io_dram_0_wdata_bits_wstrb_5),
    .io_dram_0_wdata_bits_wstrb_6(fringeCommon_io_dram_0_wdata_bits_wstrb_6),
    .io_dram_0_wdata_bits_wstrb_7(fringeCommon_io_dram_0_wdata_bits_wstrb_7),
    .io_dram_0_wdata_bits_wstrb_8(fringeCommon_io_dram_0_wdata_bits_wstrb_8),
    .io_dram_0_wdata_bits_wstrb_9(fringeCommon_io_dram_0_wdata_bits_wstrb_9),
    .io_dram_0_wdata_bits_wstrb_10(fringeCommon_io_dram_0_wdata_bits_wstrb_10),
    .io_dram_0_wdata_bits_wstrb_11(fringeCommon_io_dram_0_wdata_bits_wstrb_11),
    .io_dram_0_wdata_bits_wstrb_12(fringeCommon_io_dram_0_wdata_bits_wstrb_12),
    .io_dram_0_wdata_bits_wstrb_13(fringeCommon_io_dram_0_wdata_bits_wstrb_13),
    .io_dram_0_wdata_bits_wstrb_14(fringeCommon_io_dram_0_wdata_bits_wstrb_14),
    .io_dram_0_wdata_bits_wstrb_15(fringeCommon_io_dram_0_wdata_bits_wstrb_15),
    .io_dram_0_wdata_bits_wstrb_16(fringeCommon_io_dram_0_wdata_bits_wstrb_16),
    .io_dram_0_wdata_bits_wstrb_17(fringeCommon_io_dram_0_wdata_bits_wstrb_17),
    .io_dram_0_wdata_bits_wstrb_18(fringeCommon_io_dram_0_wdata_bits_wstrb_18),
    .io_dram_0_wdata_bits_wstrb_19(fringeCommon_io_dram_0_wdata_bits_wstrb_19),
    .io_dram_0_wdata_bits_wstrb_20(fringeCommon_io_dram_0_wdata_bits_wstrb_20),
    .io_dram_0_wdata_bits_wstrb_21(fringeCommon_io_dram_0_wdata_bits_wstrb_21),
    .io_dram_0_wdata_bits_wstrb_22(fringeCommon_io_dram_0_wdata_bits_wstrb_22),
    .io_dram_0_wdata_bits_wstrb_23(fringeCommon_io_dram_0_wdata_bits_wstrb_23),
    .io_dram_0_wdata_bits_wstrb_24(fringeCommon_io_dram_0_wdata_bits_wstrb_24),
    .io_dram_0_wdata_bits_wstrb_25(fringeCommon_io_dram_0_wdata_bits_wstrb_25),
    .io_dram_0_wdata_bits_wstrb_26(fringeCommon_io_dram_0_wdata_bits_wstrb_26),
    .io_dram_0_wdata_bits_wstrb_27(fringeCommon_io_dram_0_wdata_bits_wstrb_27),
    .io_dram_0_wdata_bits_wstrb_28(fringeCommon_io_dram_0_wdata_bits_wstrb_28),
    .io_dram_0_wdata_bits_wstrb_29(fringeCommon_io_dram_0_wdata_bits_wstrb_29),
    .io_dram_0_wdata_bits_wstrb_30(fringeCommon_io_dram_0_wdata_bits_wstrb_30),
    .io_dram_0_wdata_bits_wstrb_31(fringeCommon_io_dram_0_wdata_bits_wstrb_31),
    .io_dram_0_wdata_bits_wstrb_32(fringeCommon_io_dram_0_wdata_bits_wstrb_32),
    .io_dram_0_wdata_bits_wstrb_33(fringeCommon_io_dram_0_wdata_bits_wstrb_33),
    .io_dram_0_wdata_bits_wstrb_34(fringeCommon_io_dram_0_wdata_bits_wstrb_34),
    .io_dram_0_wdata_bits_wstrb_35(fringeCommon_io_dram_0_wdata_bits_wstrb_35),
    .io_dram_0_wdata_bits_wstrb_36(fringeCommon_io_dram_0_wdata_bits_wstrb_36),
    .io_dram_0_wdata_bits_wstrb_37(fringeCommon_io_dram_0_wdata_bits_wstrb_37),
    .io_dram_0_wdata_bits_wstrb_38(fringeCommon_io_dram_0_wdata_bits_wstrb_38),
    .io_dram_0_wdata_bits_wstrb_39(fringeCommon_io_dram_0_wdata_bits_wstrb_39),
    .io_dram_0_wdata_bits_wstrb_40(fringeCommon_io_dram_0_wdata_bits_wstrb_40),
    .io_dram_0_wdata_bits_wstrb_41(fringeCommon_io_dram_0_wdata_bits_wstrb_41),
    .io_dram_0_wdata_bits_wstrb_42(fringeCommon_io_dram_0_wdata_bits_wstrb_42),
    .io_dram_0_wdata_bits_wstrb_43(fringeCommon_io_dram_0_wdata_bits_wstrb_43),
    .io_dram_0_wdata_bits_wstrb_44(fringeCommon_io_dram_0_wdata_bits_wstrb_44),
    .io_dram_0_wdata_bits_wstrb_45(fringeCommon_io_dram_0_wdata_bits_wstrb_45),
    .io_dram_0_wdata_bits_wstrb_46(fringeCommon_io_dram_0_wdata_bits_wstrb_46),
    .io_dram_0_wdata_bits_wstrb_47(fringeCommon_io_dram_0_wdata_bits_wstrb_47),
    .io_dram_0_wdata_bits_wstrb_48(fringeCommon_io_dram_0_wdata_bits_wstrb_48),
    .io_dram_0_wdata_bits_wstrb_49(fringeCommon_io_dram_0_wdata_bits_wstrb_49),
    .io_dram_0_wdata_bits_wstrb_50(fringeCommon_io_dram_0_wdata_bits_wstrb_50),
    .io_dram_0_wdata_bits_wstrb_51(fringeCommon_io_dram_0_wdata_bits_wstrb_51),
    .io_dram_0_wdata_bits_wstrb_52(fringeCommon_io_dram_0_wdata_bits_wstrb_52),
    .io_dram_0_wdata_bits_wstrb_53(fringeCommon_io_dram_0_wdata_bits_wstrb_53),
    .io_dram_0_wdata_bits_wstrb_54(fringeCommon_io_dram_0_wdata_bits_wstrb_54),
    .io_dram_0_wdata_bits_wstrb_55(fringeCommon_io_dram_0_wdata_bits_wstrb_55),
    .io_dram_0_wdata_bits_wstrb_56(fringeCommon_io_dram_0_wdata_bits_wstrb_56),
    .io_dram_0_wdata_bits_wstrb_57(fringeCommon_io_dram_0_wdata_bits_wstrb_57),
    .io_dram_0_wdata_bits_wstrb_58(fringeCommon_io_dram_0_wdata_bits_wstrb_58),
    .io_dram_0_wdata_bits_wstrb_59(fringeCommon_io_dram_0_wdata_bits_wstrb_59),
    .io_dram_0_wdata_bits_wstrb_60(fringeCommon_io_dram_0_wdata_bits_wstrb_60),
    .io_dram_0_wdata_bits_wstrb_61(fringeCommon_io_dram_0_wdata_bits_wstrb_61),
    .io_dram_0_wdata_bits_wstrb_62(fringeCommon_io_dram_0_wdata_bits_wstrb_62),
    .io_dram_0_wdata_bits_wstrb_63(fringeCommon_io_dram_0_wdata_bits_wstrb_63),
    .io_dram_0_wdata_bits_wlast(fringeCommon_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag(fringeCommon_io_dram_0_wresp_bits_tag),
    .io_dram_1_cmd_ready(fringeCommon_io_dram_1_cmd_ready),
    .io_dram_1_cmd_valid(fringeCommon_io_dram_1_cmd_valid),
    .io_dram_1_cmd_bits_addr(fringeCommon_io_dram_1_cmd_bits_addr),
    .io_dram_1_cmd_bits_size(fringeCommon_io_dram_1_cmd_bits_size),
    .io_dram_1_cmd_bits_isWr(fringeCommon_io_dram_1_cmd_bits_isWr),
    .io_dram_1_cmd_bits_tag(fringeCommon_io_dram_1_cmd_bits_tag),
    .io_dram_1_wdata_ready(fringeCommon_io_dram_1_wdata_ready),
    .io_dram_1_wdata_valid(fringeCommon_io_dram_1_wdata_valid),
    .io_dram_1_wdata_bits_wdata_0(fringeCommon_io_dram_1_wdata_bits_wdata_0),
    .io_dram_1_wdata_bits_wdata_1(fringeCommon_io_dram_1_wdata_bits_wdata_1),
    .io_dram_1_wdata_bits_wdata_2(fringeCommon_io_dram_1_wdata_bits_wdata_2),
    .io_dram_1_wdata_bits_wdata_3(fringeCommon_io_dram_1_wdata_bits_wdata_3),
    .io_dram_1_wdata_bits_wdata_4(fringeCommon_io_dram_1_wdata_bits_wdata_4),
    .io_dram_1_wdata_bits_wdata_5(fringeCommon_io_dram_1_wdata_bits_wdata_5),
    .io_dram_1_wdata_bits_wdata_6(fringeCommon_io_dram_1_wdata_bits_wdata_6),
    .io_dram_1_wdata_bits_wdata_7(fringeCommon_io_dram_1_wdata_bits_wdata_7),
    .io_dram_1_wdata_bits_wdata_8(fringeCommon_io_dram_1_wdata_bits_wdata_8),
    .io_dram_1_wdata_bits_wdata_9(fringeCommon_io_dram_1_wdata_bits_wdata_9),
    .io_dram_1_wdata_bits_wdata_10(fringeCommon_io_dram_1_wdata_bits_wdata_10),
    .io_dram_1_wdata_bits_wdata_11(fringeCommon_io_dram_1_wdata_bits_wdata_11),
    .io_dram_1_wdata_bits_wdata_12(fringeCommon_io_dram_1_wdata_bits_wdata_12),
    .io_dram_1_wdata_bits_wdata_13(fringeCommon_io_dram_1_wdata_bits_wdata_13),
    .io_dram_1_wdata_bits_wdata_14(fringeCommon_io_dram_1_wdata_bits_wdata_14),
    .io_dram_1_wdata_bits_wdata_15(fringeCommon_io_dram_1_wdata_bits_wdata_15),
    .io_dram_1_wdata_bits_wstrb_0(fringeCommon_io_dram_1_wdata_bits_wstrb_0),
    .io_dram_1_wdata_bits_wstrb_1(fringeCommon_io_dram_1_wdata_bits_wstrb_1),
    .io_dram_1_wdata_bits_wstrb_2(fringeCommon_io_dram_1_wdata_bits_wstrb_2),
    .io_dram_1_wdata_bits_wstrb_3(fringeCommon_io_dram_1_wdata_bits_wstrb_3),
    .io_dram_1_wdata_bits_wstrb_4(fringeCommon_io_dram_1_wdata_bits_wstrb_4),
    .io_dram_1_wdata_bits_wstrb_5(fringeCommon_io_dram_1_wdata_bits_wstrb_5),
    .io_dram_1_wdata_bits_wstrb_6(fringeCommon_io_dram_1_wdata_bits_wstrb_6),
    .io_dram_1_wdata_bits_wstrb_7(fringeCommon_io_dram_1_wdata_bits_wstrb_7),
    .io_dram_1_wdata_bits_wstrb_8(fringeCommon_io_dram_1_wdata_bits_wstrb_8),
    .io_dram_1_wdata_bits_wstrb_9(fringeCommon_io_dram_1_wdata_bits_wstrb_9),
    .io_dram_1_wdata_bits_wstrb_10(fringeCommon_io_dram_1_wdata_bits_wstrb_10),
    .io_dram_1_wdata_bits_wstrb_11(fringeCommon_io_dram_1_wdata_bits_wstrb_11),
    .io_dram_1_wdata_bits_wstrb_12(fringeCommon_io_dram_1_wdata_bits_wstrb_12),
    .io_dram_1_wdata_bits_wstrb_13(fringeCommon_io_dram_1_wdata_bits_wstrb_13),
    .io_dram_1_wdata_bits_wstrb_14(fringeCommon_io_dram_1_wdata_bits_wstrb_14),
    .io_dram_1_wdata_bits_wstrb_15(fringeCommon_io_dram_1_wdata_bits_wstrb_15),
    .io_dram_1_wdata_bits_wstrb_16(fringeCommon_io_dram_1_wdata_bits_wstrb_16),
    .io_dram_1_wdata_bits_wstrb_17(fringeCommon_io_dram_1_wdata_bits_wstrb_17),
    .io_dram_1_wdata_bits_wstrb_18(fringeCommon_io_dram_1_wdata_bits_wstrb_18),
    .io_dram_1_wdata_bits_wstrb_19(fringeCommon_io_dram_1_wdata_bits_wstrb_19),
    .io_dram_1_wdata_bits_wstrb_20(fringeCommon_io_dram_1_wdata_bits_wstrb_20),
    .io_dram_1_wdata_bits_wstrb_21(fringeCommon_io_dram_1_wdata_bits_wstrb_21),
    .io_dram_1_wdata_bits_wstrb_22(fringeCommon_io_dram_1_wdata_bits_wstrb_22),
    .io_dram_1_wdata_bits_wstrb_23(fringeCommon_io_dram_1_wdata_bits_wstrb_23),
    .io_dram_1_wdata_bits_wstrb_24(fringeCommon_io_dram_1_wdata_bits_wstrb_24),
    .io_dram_1_wdata_bits_wstrb_25(fringeCommon_io_dram_1_wdata_bits_wstrb_25),
    .io_dram_1_wdata_bits_wstrb_26(fringeCommon_io_dram_1_wdata_bits_wstrb_26),
    .io_dram_1_wdata_bits_wstrb_27(fringeCommon_io_dram_1_wdata_bits_wstrb_27),
    .io_dram_1_wdata_bits_wstrb_28(fringeCommon_io_dram_1_wdata_bits_wstrb_28),
    .io_dram_1_wdata_bits_wstrb_29(fringeCommon_io_dram_1_wdata_bits_wstrb_29),
    .io_dram_1_wdata_bits_wstrb_30(fringeCommon_io_dram_1_wdata_bits_wstrb_30),
    .io_dram_1_wdata_bits_wstrb_31(fringeCommon_io_dram_1_wdata_bits_wstrb_31),
    .io_dram_1_wdata_bits_wstrb_32(fringeCommon_io_dram_1_wdata_bits_wstrb_32),
    .io_dram_1_wdata_bits_wstrb_33(fringeCommon_io_dram_1_wdata_bits_wstrb_33),
    .io_dram_1_wdata_bits_wstrb_34(fringeCommon_io_dram_1_wdata_bits_wstrb_34),
    .io_dram_1_wdata_bits_wstrb_35(fringeCommon_io_dram_1_wdata_bits_wstrb_35),
    .io_dram_1_wdata_bits_wstrb_36(fringeCommon_io_dram_1_wdata_bits_wstrb_36),
    .io_dram_1_wdata_bits_wstrb_37(fringeCommon_io_dram_1_wdata_bits_wstrb_37),
    .io_dram_1_wdata_bits_wstrb_38(fringeCommon_io_dram_1_wdata_bits_wstrb_38),
    .io_dram_1_wdata_bits_wstrb_39(fringeCommon_io_dram_1_wdata_bits_wstrb_39),
    .io_dram_1_wdata_bits_wstrb_40(fringeCommon_io_dram_1_wdata_bits_wstrb_40),
    .io_dram_1_wdata_bits_wstrb_41(fringeCommon_io_dram_1_wdata_bits_wstrb_41),
    .io_dram_1_wdata_bits_wstrb_42(fringeCommon_io_dram_1_wdata_bits_wstrb_42),
    .io_dram_1_wdata_bits_wstrb_43(fringeCommon_io_dram_1_wdata_bits_wstrb_43),
    .io_dram_1_wdata_bits_wstrb_44(fringeCommon_io_dram_1_wdata_bits_wstrb_44),
    .io_dram_1_wdata_bits_wstrb_45(fringeCommon_io_dram_1_wdata_bits_wstrb_45),
    .io_dram_1_wdata_bits_wstrb_46(fringeCommon_io_dram_1_wdata_bits_wstrb_46),
    .io_dram_1_wdata_bits_wstrb_47(fringeCommon_io_dram_1_wdata_bits_wstrb_47),
    .io_dram_1_wdata_bits_wstrb_48(fringeCommon_io_dram_1_wdata_bits_wstrb_48),
    .io_dram_1_wdata_bits_wstrb_49(fringeCommon_io_dram_1_wdata_bits_wstrb_49),
    .io_dram_1_wdata_bits_wstrb_50(fringeCommon_io_dram_1_wdata_bits_wstrb_50),
    .io_dram_1_wdata_bits_wstrb_51(fringeCommon_io_dram_1_wdata_bits_wstrb_51),
    .io_dram_1_wdata_bits_wstrb_52(fringeCommon_io_dram_1_wdata_bits_wstrb_52),
    .io_dram_1_wdata_bits_wstrb_53(fringeCommon_io_dram_1_wdata_bits_wstrb_53),
    .io_dram_1_wdata_bits_wstrb_54(fringeCommon_io_dram_1_wdata_bits_wstrb_54),
    .io_dram_1_wdata_bits_wstrb_55(fringeCommon_io_dram_1_wdata_bits_wstrb_55),
    .io_dram_1_wdata_bits_wstrb_56(fringeCommon_io_dram_1_wdata_bits_wstrb_56),
    .io_dram_1_wdata_bits_wstrb_57(fringeCommon_io_dram_1_wdata_bits_wstrb_57),
    .io_dram_1_wdata_bits_wstrb_58(fringeCommon_io_dram_1_wdata_bits_wstrb_58),
    .io_dram_1_wdata_bits_wstrb_59(fringeCommon_io_dram_1_wdata_bits_wstrb_59),
    .io_dram_1_wdata_bits_wstrb_60(fringeCommon_io_dram_1_wdata_bits_wstrb_60),
    .io_dram_1_wdata_bits_wstrb_61(fringeCommon_io_dram_1_wdata_bits_wstrb_61),
    .io_dram_1_wdata_bits_wstrb_62(fringeCommon_io_dram_1_wdata_bits_wstrb_62),
    .io_dram_1_wdata_bits_wstrb_63(fringeCommon_io_dram_1_wdata_bits_wstrb_63),
    .io_dram_1_wdata_bits_wlast(fringeCommon_io_dram_1_wdata_bits_wlast),
    .io_dram_1_rresp_ready(fringeCommon_io_dram_1_rresp_ready),
    .io_dram_1_wresp_ready(fringeCommon_io_dram_1_wresp_ready),
    .io_dram_1_wresp_valid(fringeCommon_io_dram_1_wresp_valid),
    .io_dram_1_wresp_bits_tag(fringeCommon_io_dram_1_wresp_bits_tag),
    .io_dram_2_cmd_ready(fringeCommon_io_dram_2_cmd_ready),
    .io_dram_2_cmd_valid(fringeCommon_io_dram_2_cmd_valid),
    .io_dram_2_cmd_bits_addr(fringeCommon_io_dram_2_cmd_bits_addr),
    .io_dram_2_cmd_bits_size(fringeCommon_io_dram_2_cmd_bits_size),
    .io_dram_2_cmd_bits_isWr(fringeCommon_io_dram_2_cmd_bits_isWr),
    .io_dram_2_cmd_bits_tag(fringeCommon_io_dram_2_cmd_bits_tag),
    .io_dram_2_wdata_ready(fringeCommon_io_dram_2_wdata_ready),
    .io_dram_2_wdata_valid(fringeCommon_io_dram_2_wdata_valid),
    .io_dram_2_wdata_bits_wdata_0(fringeCommon_io_dram_2_wdata_bits_wdata_0),
    .io_dram_2_wdata_bits_wdata_1(fringeCommon_io_dram_2_wdata_bits_wdata_1),
    .io_dram_2_wdata_bits_wdata_2(fringeCommon_io_dram_2_wdata_bits_wdata_2),
    .io_dram_2_wdata_bits_wdata_3(fringeCommon_io_dram_2_wdata_bits_wdata_3),
    .io_dram_2_wdata_bits_wdata_4(fringeCommon_io_dram_2_wdata_bits_wdata_4),
    .io_dram_2_wdata_bits_wdata_5(fringeCommon_io_dram_2_wdata_bits_wdata_5),
    .io_dram_2_wdata_bits_wdata_6(fringeCommon_io_dram_2_wdata_bits_wdata_6),
    .io_dram_2_wdata_bits_wdata_7(fringeCommon_io_dram_2_wdata_bits_wdata_7),
    .io_dram_2_wdata_bits_wdata_8(fringeCommon_io_dram_2_wdata_bits_wdata_8),
    .io_dram_2_wdata_bits_wdata_9(fringeCommon_io_dram_2_wdata_bits_wdata_9),
    .io_dram_2_wdata_bits_wdata_10(fringeCommon_io_dram_2_wdata_bits_wdata_10),
    .io_dram_2_wdata_bits_wdata_11(fringeCommon_io_dram_2_wdata_bits_wdata_11),
    .io_dram_2_wdata_bits_wdata_12(fringeCommon_io_dram_2_wdata_bits_wdata_12),
    .io_dram_2_wdata_bits_wdata_13(fringeCommon_io_dram_2_wdata_bits_wdata_13),
    .io_dram_2_wdata_bits_wdata_14(fringeCommon_io_dram_2_wdata_bits_wdata_14),
    .io_dram_2_wdata_bits_wdata_15(fringeCommon_io_dram_2_wdata_bits_wdata_15),
    .io_dram_2_wdata_bits_wstrb_0(fringeCommon_io_dram_2_wdata_bits_wstrb_0),
    .io_dram_2_wdata_bits_wstrb_1(fringeCommon_io_dram_2_wdata_bits_wstrb_1),
    .io_dram_2_wdata_bits_wstrb_2(fringeCommon_io_dram_2_wdata_bits_wstrb_2),
    .io_dram_2_wdata_bits_wstrb_3(fringeCommon_io_dram_2_wdata_bits_wstrb_3),
    .io_dram_2_wdata_bits_wstrb_4(fringeCommon_io_dram_2_wdata_bits_wstrb_4),
    .io_dram_2_wdata_bits_wstrb_5(fringeCommon_io_dram_2_wdata_bits_wstrb_5),
    .io_dram_2_wdata_bits_wstrb_6(fringeCommon_io_dram_2_wdata_bits_wstrb_6),
    .io_dram_2_wdata_bits_wstrb_7(fringeCommon_io_dram_2_wdata_bits_wstrb_7),
    .io_dram_2_wdata_bits_wstrb_8(fringeCommon_io_dram_2_wdata_bits_wstrb_8),
    .io_dram_2_wdata_bits_wstrb_9(fringeCommon_io_dram_2_wdata_bits_wstrb_9),
    .io_dram_2_wdata_bits_wstrb_10(fringeCommon_io_dram_2_wdata_bits_wstrb_10),
    .io_dram_2_wdata_bits_wstrb_11(fringeCommon_io_dram_2_wdata_bits_wstrb_11),
    .io_dram_2_wdata_bits_wstrb_12(fringeCommon_io_dram_2_wdata_bits_wstrb_12),
    .io_dram_2_wdata_bits_wstrb_13(fringeCommon_io_dram_2_wdata_bits_wstrb_13),
    .io_dram_2_wdata_bits_wstrb_14(fringeCommon_io_dram_2_wdata_bits_wstrb_14),
    .io_dram_2_wdata_bits_wstrb_15(fringeCommon_io_dram_2_wdata_bits_wstrb_15),
    .io_dram_2_wdata_bits_wstrb_16(fringeCommon_io_dram_2_wdata_bits_wstrb_16),
    .io_dram_2_wdata_bits_wstrb_17(fringeCommon_io_dram_2_wdata_bits_wstrb_17),
    .io_dram_2_wdata_bits_wstrb_18(fringeCommon_io_dram_2_wdata_bits_wstrb_18),
    .io_dram_2_wdata_bits_wstrb_19(fringeCommon_io_dram_2_wdata_bits_wstrb_19),
    .io_dram_2_wdata_bits_wstrb_20(fringeCommon_io_dram_2_wdata_bits_wstrb_20),
    .io_dram_2_wdata_bits_wstrb_21(fringeCommon_io_dram_2_wdata_bits_wstrb_21),
    .io_dram_2_wdata_bits_wstrb_22(fringeCommon_io_dram_2_wdata_bits_wstrb_22),
    .io_dram_2_wdata_bits_wstrb_23(fringeCommon_io_dram_2_wdata_bits_wstrb_23),
    .io_dram_2_wdata_bits_wstrb_24(fringeCommon_io_dram_2_wdata_bits_wstrb_24),
    .io_dram_2_wdata_bits_wstrb_25(fringeCommon_io_dram_2_wdata_bits_wstrb_25),
    .io_dram_2_wdata_bits_wstrb_26(fringeCommon_io_dram_2_wdata_bits_wstrb_26),
    .io_dram_2_wdata_bits_wstrb_27(fringeCommon_io_dram_2_wdata_bits_wstrb_27),
    .io_dram_2_wdata_bits_wstrb_28(fringeCommon_io_dram_2_wdata_bits_wstrb_28),
    .io_dram_2_wdata_bits_wstrb_29(fringeCommon_io_dram_2_wdata_bits_wstrb_29),
    .io_dram_2_wdata_bits_wstrb_30(fringeCommon_io_dram_2_wdata_bits_wstrb_30),
    .io_dram_2_wdata_bits_wstrb_31(fringeCommon_io_dram_2_wdata_bits_wstrb_31),
    .io_dram_2_wdata_bits_wstrb_32(fringeCommon_io_dram_2_wdata_bits_wstrb_32),
    .io_dram_2_wdata_bits_wstrb_33(fringeCommon_io_dram_2_wdata_bits_wstrb_33),
    .io_dram_2_wdata_bits_wstrb_34(fringeCommon_io_dram_2_wdata_bits_wstrb_34),
    .io_dram_2_wdata_bits_wstrb_35(fringeCommon_io_dram_2_wdata_bits_wstrb_35),
    .io_dram_2_wdata_bits_wstrb_36(fringeCommon_io_dram_2_wdata_bits_wstrb_36),
    .io_dram_2_wdata_bits_wstrb_37(fringeCommon_io_dram_2_wdata_bits_wstrb_37),
    .io_dram_2_wdata_bits_wstrb_38(fringeCommon_io_dram_2_wdata_bits_wstrb_38),
    .io_dram_2_wdata_bits_wstrb_39(fringeCommon_io_dram_2_wdata_bits_wstrb_39),
    .io_dram_2_wdata_bits_wstrb_40(fringeCommon_io_dram_2_wdata_bits_wstrb_40),
    .io_dram_2_wdata_bits_wstrb_41(fringeCommon_io_dram_2_wdata_bits_wstrb_41),
    .io_dram_2_wdata_bits_wstrb_42(fringeCommon_io_dram_2_wdata_bits_wstrb_42),
    .io_dram_2_wdata_bits_wstrb_43(fringeCommon_io_dram_2_wdata_bits_wstrb_43),
    .io_dram_2_wdata_bits_wstrb_44(fringeCommon_io_dram_2_wdata_bits_wstrb_44),
    .io_dram_2_wdata_bits_wstrb_45(fringeCommon_io_dram_2_wdata_bits_wstrb_45),
    .io_dram_2_wdata_bits_wstrb_46(fringeCommon_io_dram_2_wdata_bits_wstrb_46),
    .io_dram_2_wdata_bits_wstrb_47(fringeCommon_io_dram_2_wdata_bits_wstrb_47),
    .io_dram_2_wdata_bits_wstrb_48(fringeCommon_io_dram_2_wdata_bits_wstrb_48),
    .io_dram_2_wdata_bits_wstrb_49(fringeCommon_io_dram_2_wdata_bits_wstrb_49),
    .io_dram_2_wdata_bits_wstrb_50(fringeCommon_io_dram_2_wdata_bits_wstrb_50),
    .io_dram_2_wdata_bits_wstrb_51(fringeCommon_io_dram_2_wdata_bits_wstrb_51),
    .io_dram_2_wdata_bits_wstrb_52(fringeCommon_io_dram_2_wdata_bits_wstrb_52),
    .io_dram_2_wdata_bits_wstrb_53(fringeCommon_io_dram_2_wdata_bits_wstrb_53),
    .io_dram_2_wdata_bits_wstrb_54(fringeCommon_io_dram_2_wdata_bits_wstrb_54),
    .io_dram_2_wdata_bits_wstrb_55(fringeCommon_io_dram_2_wdata_bits_wstrb_55),
    .io_dram_2_wdata_bits_wstrb_56(fringeCommon_io_dram_2_wdata_bits_wstrb_56),
    .io_dram_2_wdata_bits_wstrb_57(fringeCommon_io_dram_2_wdata_bits_wstrb_57),
    .io_dram_2_wdata_bits_wstrb_58(fringeCommon_io_dram_2_wdata_bits_wstrb_58),
    .io_dram_2_wdata_bits_wstrb_59(fringeCommon_io_dram_2_wdata_bits_wstrb_59),
    .io_dram_2_wdata_bits_wstrb_60(fringeCommon_io_dram_2_wdata_bits_wstrb_60),
    .io_dram_2_wdata_bits_wstrb_61(fringeCommon_io_dram_2_wdata_bits_wstrb_61),
    .io_dram_2_wdata_bits_wstrb_62(fringeCommon_io_dram_2_wdata_bits_wstrb_62),
    .io_dram_2_wdata_bits_wstrb_63(fringeCommon_io_dram_2_wdata_bits_wstrb_63),
    .io_dram_2_wdata_bits_wlast(fringeCommon_io_dram_2_wdata_bits_wlast),
    .io_dram_2_rresp_ready(fringeCommon_io_dram_2_rresp_ready),
    .io_dram_2_wresp_ready(fringeCommon_io_dram_2_wresp_ready),
    .io_dram_2_wresp_valid(fringeCommon_io_dram_2_wresp_valid),
    .io_dram_2_wresp_bits_tag(fringeCommon_io_dram_2_wresp_bits_tag),
    .io_dram_3_cmd_ready(fringeCommon_io_dram_3_cmd_ready),
    .io_dram_3_cmd_valid(fringeCommon_io_dram_3_cmd_valid),
    .io_dram_3_cmd_bits_addr(fringeCommon_io_dram_3_cmd_bits_addr),
    .io_dram_3_cmd_bits_size(fringeCommon_io_dram_3_cmd_bits_size),
    .io_dram_3_cmd_bits_isWr(fringeCommon_io_dram_3_cmd_bits_isWr),
    .io_dram_3_cmd_bits_tag(fringeCommon_io_dram_3_cmd_bits_tag),
    .io_dram_3_wdata_ready(fringeCommon_io_dram_3_wdata_ready),
    .io_dram_3_wdata_valid(fringeCommon_io_dram_3_wdata_valid),
    .io_dram_3_wdata_bits_wdata_0(fringeCommon_io_dram_3_wdata_bits_wdata_0),
    .io_dram_3_wdata_bits_wdata_1(fringeCommon_io_dram_3_wdata_bits_wdata_1),
    .io_dram_3_wdata_bits_wdata_2(fringeCommon_io_dram_3_wdata_bits_wdata_2),
    .io_dram_3_wdata_bits_wdata_3(fringeCommon_io_dram_3_wdata_bits_wdata_3),
    .io_dram_3_wdata_bits_wdata_4(fringeCommon_io_dram_3_wdata_bits_wdata_4),
    .io_dram_3_wdata_bits_wdata_5(fringeCommon_io_dram_3_wdata_bits_wdata_5),
    .io_dram_3_wdata_bits_wdata_6(fringeCommon_io_dram_3_wdata_bits_wdata_6),
    .io_dram_3_wdata_bits_wdata_7(fringeCommon_io_dram_3_wdata_bits_wdata_7),
    .io_dram_3_wdata_bits_wdata_8(fringeCommon_io_dram_3_wdata_bits_wdata_8),
    .io_dram_3_wdata_bits_wdata_9(fringeCommon_io_dram_3_wdata_bits_wdata_9),
    .io_dram_3_wdata_bits_wdata_10(fringeCommon_io_dram_3_wdata_bits_wdata_10),
    .io_dram_3_wdata_bits_wdata_11(fringeCommon_io_dram_3_wdata_bits_wdata_11),
    .io_dram_3_wdata_bits_wdata_12(fringeCommon_io_dram_3_wdata_bits_wdata_12),
    .io_dram_3_wdata_bits_wdata_13(fringeCommon_io_dram_3_wdata_bits_wdata_13),
    .io_dram_3_wdata_bits_wdata_14(fringeCommon_io_dram_3_wdata_bits_wdata_14),
    .io_dram_3_wdata_bits_wdata_15(fringeCommon_io_dram_3_wdata_bits_wdata_15),
    .io_dram_3_wdata_bits_wstrb_0(fringeCommon_io_dram_3_wdata_bits_wstrb_0),
    .io_dram_3_wdata_bits_wstrb_1(fringeCommon_io_dram_3_wdata_bits_wstrb_1),
    .io_dram_3_wdata_bits_wstrb_2(fringeCommon_io_dram_3_wdata_bits_wstrb_2),
    .io_dram_3_wdata_bits_wstrb_3(fringeCommon_io_dram_3_wdata_bits_wstrb_3),
    .io_dram_3_wdata_bits_wstrb_4(fringeCommon_io_dram_3_wdata_bits_wstrb_4),
    .io_dram_3_wdata_bits_wstrb_5(fringeCommon_io_dram_3_wdata_bits_wstrb_5),
    .io_dram_3_wdata_bits_wstrb_6(fringeCommon_io_dram_3_wdata_bits_wstrb_6),
    .io_dram_3_wdata_bits_wstrb_7(fringeCommon_io_dram_3_wdata_bits_wstrb_7),
    .io_dram_3_wdata_bits_wstrb_8(fringeCommon_io_dram_3_wdata_bits_wstrb_8),
    .io_dram_3_wdata_bits_wstrb_9(fringeCommon_io_dram_3_wdata_bits_wstrb_9),
    .io_dram_3_wdata_bits_wstrb_10(fringeCommon_io_dram_3_wdata_bits_wstrb_10),
    .io_dram_3_wdata_bits_wstrb_11(fringeCommon_io_dram_3_wdata_bits_wstrb_11),
    .io_dram_3_wdata_bits_wstrb_12(fringeCommon_io_dram_3_wdata_bits_wstrb_12),
    .io_dram_3_wdata_bits_wstrb_13(fringeCommon_io_dram_3_wdata_bits_wstrb_13),
    .io_dram_3_wdata_bits_wstrb_14(fringeCommon_io_dram_3_wdata_bits_wstrb_14),
    .io_dram_3_wdata_bits_wstrb_15(fringeCommon_io_dram_3_wdata_bits_wstrb_15),
    .io_dram_3_wdata_bits_wstrb_16(fringeCommon_io_dram_3_wdata_bits_wstrb_16),
    .io_dram_3_wdata_bits_wstrb_17(fringeCommon_io_dram_3_wdata_bits_wstrb_17),
    .io_dram_3_wdata_bits_wstrb_18(fringeCommon_io_dram_3_wdata_bits_wstrb_18),
    .io_dram_3_wdata_bits_wstrb_19(fringeCommon_io_dram_3_wdata_bits_wstrb_19),
    .io_dram_3_wdata_bits_wstrb_20(fringeCommon_io_dram_3_wdata_bits_wstrb_20),
    .io_dram_3_wdata_bits_wstrb_21(fringeCommon_io_dram_3_wdata_bits_wstrb_21),
    .io_dram_3_wdata_bits_wstrb_22(fringeCommon_io_dram_3_wdata_bits_wstrb_22),
    .io_dram_3_wdata_bits_wstrb_23(fringeCommon_io_dram_3_wdata_bits_wstrb_23),
    .io_dram_3_wdata_bits_wstrb_24(fringeCommon_io_dram_3_wdata_bits_wstrb_24),
    .io_dram_3_wdata_bits_wstrb_25(fringeCommon_io_dram_3_wdata_bits_wstrb_25),
    .io_dram_3_wdata_bits_wstrb_26(fringeCommon_io_dram_3_wdata_bits_wstrb_26),
    .io_dram_3_wdata_bits_wstrb_27(fringeCommon_io_dram_3_wdata_bits_wstrb_27),
    .io_dram_3_wdata_bits_wstrb_28(fringeCommon_io_dram_3_wdata_bits_wstrb_28),
    .io_dram_3_wdata_bits_wstrb_29(fringeCommon_io_dram_3_wdata_bits_wstrb_29),
    .io_dram_3_wdata_bits_wstrb_30(fringeCommon_io_dram_3_wdata_bits_wstrb_30),
    .io_dram_3_wdata_bits_wstrb_31(fringeCommon_io_dram_3_wdata_bits_wstrb_31),
    .io_dram_3_wdata_bits_wstrb_32(fringeCommon_io_dram_3_wdata_bits_wstrb_32),
    .io_dram_3_wdata_bits_wstrb_33(fringeCommon_io_dram_3_wdata_bits_wstrb_33),
    .io_dram_3_wdata_bits_wstrb_34(fringeCommon_io_dram_3_wdata_bits_wstrb_34),
    .io_dram_3_wdata_bits_wstrb_35(fringeCommon_io_dram_3_wdata_bits_wstrb_35),
    .io_dram_3_wdata_bits_wstrb_36(fringeCommon_io_dram_3_wdata_bits_wstrb_36),
    .io_dram_3_wdata_bits_wstrb_37(fringeCommon_io_dram_3_wdata_bits_wstrb_37),
    .io_dram_3_wdata_bits_wstrb_38(fringeCommon_io_dram_3_wdata_bits_wstrb_38),
    .io_dram_3_wdata_bits_wstrb_39(fringeCommon_io_dram_3_wdata_bits_wstrb_39),
    .io_dram_3_wdata_bits_wstrb_40(fringeCommon_io_dram_3_wdata_bits_wstrb_40),
    .io_dram_3_wdata_bits_wstrb_41(fringeCommon_io_dram_3_wdata_bits_wstrb_41),
    .io_dram_3_wdata_bits_wstrb_42(fringeCommon_io_dram_3_wdata_bits_wstrb_42),
    .io_dram_3_wdata_bits_wstrb_43(fringeCommon_io_dram_3_wdata_bits_wstrb_43),
    .io_dram_3_wdata_bits_wstrb_44(fringeCommon_io_dram_3_wdata_bits_wstrb_44),
    .io_dram_3_wdata_bits_wstrb_45(fringeCommon_io_dram_3_wdata_bits_wstrb_45),
    .io_dram_3_wdata_bits_wstrb_46(fringeCommon_io_dram_3_wdata_bits_wstrb_46),
    .io_dram_3_wdata_bits_wstrb_47(fringeCommon_io_dram_3_wdata_bits_wstrb_47),
    .io_dram_3_wdata_bits_wstrb_48(fringeCommon_io_dram_3_wdata_bits_wstrb_48),
    .io_dram_3_wdata_bits_wstrb_49(fringeCommon_io_dram_3_wdata_bits_wstrb_49),
    .io_dram_3_wdata_bits_wstrb_50(fringeCommon_io_dram_3_wdata_bits_wstrb_50),
    .io_dram_3_wdata_bits_wstrb_51(fringeCommon_io_dram_3_wdata_bits_wstrb_51),
    .io_dram_3_wdata_bits_wstrb_52(fringeCommon_io_dram_3_wdata_bits_wstrb_52),
    .io_dram_3_wdata_bits_wstrb_53(fringeCommon_io_dram_3_wdata_bits_wstrb_53),
    .io_dram_3_wdata_bits_wstrb_54(fringeCommon_io_dram_3_wdata_bits_wstrb_54),
    .io_dram_3_wdata_bits_wstrb_55(fringeCommon_io_dram_3_wdata_bits_wstrb_55),
    .io_dram_3_wdata_bits_wstrb_56(fringeCommon_io_dram_3_wdata_bits_wstrb_56),
    .io_dram_3_wdata_bits_wstrb_57(fringeCommon_io_dram_3_wdata_bits_wstrb_57),
    .io_dram_3_wdata_bits_wstrb_58(fringeCommon_io_dram_3_wdata_bits_wstrb_58),
    .io_dram_3_wdata_bits_wstrb_59(fringeCommon_io_dram_3_wdata_bits_wstrb_59),
    .io_dram_3_wdata_bits_wstrb_60(fringeCommon_io_dram_3_wdata_bits_wstrb_60),
    .io_dram_3_wdata_bits_wstrb_61(fringeCommon_io_dram_3_wdata_bits_wstrb_61),
    .io_dram_3_wdata_bits_wstrb_62(fringeCommon_io_dram_3_wdata_bits_wstrb_62),
    .io_dram_3_wdata_bits_wstrb_63(fringeCommon_io_dram_3_wdata_bits_wstrb_63),
    .io_dram_3_wdata_bits_wlast(fringeCommon_io_dram_3_wdata_bits_wlast),
    .io_dram_3_rresp_ready(fringeCommon_io_dram_3_rresp_ready),
    .io_dram_3_wresp_ready(fringeCommon_io_dram_3_wresp_ready),
    .io_dram_3_wresp_valid(fringeCommon_io_dram_3_wresp_valid),
    .io_dram_3_wresp_bits_tag(fringeCommon_io_dram_3_wresp_bits_tag),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridge AXI4LiteToRFBridge ( // @[FringeZynq.scala 90:31:@163030.4]
    .clock(AXI4LiteToRFBridge_clock),
    .reset(AXI4LiteToRFBridge_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridge_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridge_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridge_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridge_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridge_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridge_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridge_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridge_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridge_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridge_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridge_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridge_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridge_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridge_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridge_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridge_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridge_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridge_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridge_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridge_io_raddr),
    .io_wen(AXI4LiteToRFBridge_io_wen),
    .io_waddr(AXI4LiteToRFBridge_io_waddr),
    .io_wdata(AXI4LiteToRFBridge_io_wdata),
    .io_rdata(AXI4LiteToRFBridge_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 131:27:@163180.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_1 ( // @[FringeZynq.scala 131:27:@163336.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_1_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_1_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_1_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_1_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_1_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_1_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_1_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_1_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_1_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_1_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_1_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_1_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_1_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_1_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_1_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_1_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_1_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_1_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_1_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_1_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_1_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_1_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_1_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_1_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_1_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_1_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_1_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_1_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_1_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_1_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_1_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_1_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_2 ( // @[FringeZynq.scala 131:27:@163492.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_2_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_2_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_2_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_2_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_2_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_2_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_2_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_2_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_2_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_2_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_2_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_2_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_2_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_2_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_2_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_2_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_2_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_2_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_2_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_2_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_2_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_2_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_2_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_2_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_2_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_2_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_2_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_2_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_2_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_2_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_2_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_2_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_3 ( // @[FringeZynq.scala 131:27:@163648.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_3_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_3_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_3_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_3_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_3_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_3_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_3_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_3_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_3_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_3_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_3_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_3_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_3_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_3_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_3_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_3_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_3_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_3_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_3_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_3_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_3_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_3_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_3_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_3_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_3_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_3_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_3_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_3_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_3_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_3_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_3_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_3_io_M_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 91:28:@163048.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 91:28:@163044.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 91:28:@163040.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 91:28:@163039.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 91:28:@163038.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 91:28:@163037.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 91:28:@163035.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 91:28:@163034.4]
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@163335.4]
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@163333.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@163332.4]
  assign io_M_AXI_0_AWVALID = MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@163325.4]
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@163323.4]
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@163321.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@163320.4]
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@163313.4]
  assign io_M_AXI_0_WDATA = MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@163311.4]
  assign io_M_AXI_0_WSTRB = MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@163310.4]
  assign io_M_AXI_0_WLAST = MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@163309.4]
  assign io_M_AXI_0_WVALID = MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@163308.4]
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@163300.4]
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@163295.4]
  assign io_M_AXI_1_AWID = MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@163491.4]
  assign io_M_AXI_1_AWADDR = MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@163489.4]
  assign io_M_AXI_1_AWLEN = MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@163488.4]
  assign io_M_AXI_1_AWVALID = MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@163481.4]
  assign io_M_AXI_1_ARID = MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@163479.4]
  assign io_M_AXI_1_ARADDR = MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@163477.4]
  assign io_M_AXI_1_ARLEN = MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@163476.4]
  assign io_M_AXI_1_ARVALID = MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@163469.4]
  assign io_M_AXI_1_WDATA = MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@163467.4]
  assign io_M_AXI_1_WSTRB = MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@163466.4]
  assign io_M_AXI_1_WLAST = MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@163465.4]
  assign io_M_AXI_1_WVALID = MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@163464.4]
  assign io_M_AXI_1_RREADY = MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@163456.4]
  assign io_M_AXI_1_BREADY = MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@163451.4]
  assign io_M_AXI_2_AWID = MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@163647.4]
  assign io_M_AXI_2_AWADDR = MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@163645.4]
  assign io_M_AXI_2_AWLEN = MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@163644.4]
  assign io_M_AXI_2_AWVALID = MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@163637.4]
  assign io_M_AXI_2_ARID = MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@163635.4]
  assign io_M_AXI_2_ARADDR = MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@163633.4]
  assign io_M_AXI_2_ARLEN = MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@163632.4]
  assign io_M_AXI_2_ARVALID = MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@163625.4]
  assign io_M_AXI_2_WDATA = MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@163623.4]
  assign io_M_AXI_2_WSTRB = MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@163622.4]
  assign io_M_AXI_2_WLAST = MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@163621.4]
  assign io_M_AXI_2_WVALID = MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@163620.4]
  assign io_M_AXI_2_RREADY = MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@163612.4]
  assign io_M_AXI_2_BREADY = MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@163607.4]
  assign io_M_AXI_3_AWID = MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@163803.4]
  assign io_M_AXI_3_AWADDR = MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@163801.4]
  assign io_M_AXI_3_AWLEN = MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@163800.4]
  assign io_M_AXI_3_AWVALID = MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@163793.4]
  assign io_M_AXI_3_ARID = MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@163791.4]
  assign io_M_AXI_3_ARADDR = MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@163789.4]
  assign io_M_AXI_3_ARLEN = MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@163788.4]
  assign io_M_AXI_3_ARVALID = MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@163781.4]
  assign io_M_AXI_3_WDATA = MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@163779.4]
  assign io_M_AXI_3_WSTRB = MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@163778.4]
  assign io_M_AXI_3_WLAST = MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@163777.4]
  assign io_M_AXI_3_WVALID = MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@163776.4]
  assign io_M_AXI_3_RREADY = MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@163768.4]
  assign io_M_AXI_3_BREADY = MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@163763.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 115:13:@163058.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 119:12:@163062.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 121:13:@163063.4]
  assign io_argIns_1 = fringeCommon_io_argIns_1; // @[FringeZynq.scala 121:13:@163064.4]
  assign io_memStreams_stores_0_cmd_ready = fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 126:17:@163151.4]
  assign io_memStreams_stores_0_data_ready = fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 126:17:@163147.4]
  assign io_memStreams_stores_0_wresp_valid = fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 126:17:@163142.4]
  assign io_memStreams_stores_0_wresp_bits = fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 126:17:@163141.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 127:11:@163176.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 127:11:@163175.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 127:11:@163174.4]
  assign fringeCommon_clock = clock; // @[:@162125.4]
  assign fringeCommon_reset = reset; // @[:@162126.4 FringeZynq.scala 117:22:@163061.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 94:27:@163052.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 95:27:@163053.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 96:27:@163054.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridge_io_wdata}; // @[FringeZynq.scala 97:27:@163055.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 116:24:@163059.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 122:27:@163066.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 122:27:@163065.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 126:17:@163150.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 126:17:@163149.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 126:17:@163148.4]
  assign fringeCommon_io_memStreams_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 126:17:@163146.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 126:17:@163145.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 126:17:@163144.4]
  assign fringeCommon_io_memStreams_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 126:17:@163143.4]
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@163294.4]
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@163287.4]
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@163184.4]
  assign fringeCommon_io_dram_0_wresp_bits_tag = MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@163183.4]
  assign fringeCommon_io_dram_1_cmd_ready = MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@163450.4]
  assign fringeCommon_io_dram_1_wdata_ready = MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@163443.4]
  assign fringeCommon_io_dram_1_wresp_valid = MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@163340.4]
  assign fringeCommon_io_dram_1_wresp_bits_tag = MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@163339.4]
  assign fringeCommon_io_dram_2_cmd_ready = MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@163606.4]
  assign fringeCommon_io_dram_2_wdata_ready = MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@163599.4]
  assign fringeCommon_io_dram_2_wresp_valid = MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@163496.4]
  assign fringeCommon_io_dram_2_wresp_bits_tag = MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@163495.4]
  assign fringeCommon_io_dram_3_cmd_ready = MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@163762.4]
  assign fringeCommon_io_dram_3_wdata_ready = MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@163755.4]
  assign fringeCommon_io_dram_3_wresp_valid = MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@163652.4]
  assign fringeCommon_io_dram_3_wresp_bits_tag = MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@163651.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 127:11:@163179.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 127:11:@163178.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 127:11:@163177.4]
  assign AXI4LiteToRFBridge_clock = clock; // @[:@163031.4]
  assign AXI4LiteToRFBridge_reset = reset; // @[:@163032.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 91:28:@163051.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 91:28:@163050.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 91:28:@163049.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 91:28:@163047.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 91:28:@163046.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 91:28:@163045.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 91:28:@163043.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 91:28:@163042.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 91:28:@163041.4]
  assign AXI4LiteToRFBridge_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 91:28:@163036.4]
  assign AXI4LiteToRFBridge_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 91:28:@163033.4]
  assign AXI4LiteToRFBridge_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 98:28:@163056.4]
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 132:21:@163293.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 132:21:@163292.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 132:21:@163291.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_isWr = fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@163289.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag = fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 132:21:@163288.4]
  assign MAGToAXI4Bridge_io_in_wdata_valid = fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 132:21:@163286.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@163270.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@163271.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@163272.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@163273.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@163274.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@163275.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@163276.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@163277.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@163278.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@163279.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@163280.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@163281.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@163282.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@163283.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@163284.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@163285.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@163206.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@163207.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@163208.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@163209.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@163210.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@163211.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@163212.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@163213.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@163214.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@163215.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@163216.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@163217.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@163218.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@163219.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@163220.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@163221.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@163222.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@163223.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@163224.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@163225.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@163226.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@163227.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@163228.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@163229.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@163230.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@163231.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@163232.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@163233.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@163234.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@163235.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@163236.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@163237.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@163238.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@163239.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@163240.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@163241.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@163242.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@163243.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@163244.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@163245.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@163246.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@163247.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@163248.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@163249.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@163250.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@163251.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@163252.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@163253.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@163254.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@163255.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@163256.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@163257.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@163258.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@163259.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@163260.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@163261.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@163262.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@163263.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@163264.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@163265.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@163266.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@163267.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@163268.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@163269.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wlast = fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@163205.4]
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 132:21:@163204.4]
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 132:21:@163185.4]
  assign MAGToAXI4Bridge_io_M_AXI_AWREADY = io_M_AXI_0_AWREADY; // @[FringeZynq.scala 133:10:@163324.4]
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY; // @[FringeZynq.scala 133:10:@163312.4]
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY; // @[FringeZynq.scala 133:10:@163307.4]
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID; // @[FringeZynq.scala 133:10:@163299.4]
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID; // @[FringeZynq.scala 133:10:@163296.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_valid = fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 132:21:@163449.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_addr = fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 132:21:@163448.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_size = fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 132:21:@163447.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_isWr = fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@163445.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_tag = fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 132:21:@163444.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_valid = fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 132:21:@163442.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@163426.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@163427.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@163428.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@163429.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@163430.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@163431.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@163432.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@163433.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@163434.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@163435.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@163436.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@163437.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@163438.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@163439.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@163440.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@163441.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@163362.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@163363.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@163364.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@163365.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@163366.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@163367.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@163368.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@163369.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@163370.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@163371.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@163372.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@163373.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@163374.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@163375.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@163376.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@163377.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@163378.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@163379.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@163380.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@163381.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@163382.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@163383.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@163384.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@163385.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@163386.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@163387.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@163388.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@163389.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@163390.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@163391.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@163392.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@163393.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@163394.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@163395.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@163396.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@163397.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@163398.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@163399.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@163400.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@163401.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@163402.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@163403.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@163404.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@163405.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@163406.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@163407.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@163408.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@163409.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@163410.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@163411.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@163412.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@163413.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@163414.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@163415.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@163416.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@163417.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@163418.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@163419.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@163420.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@163421.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@163422.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@163423.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@163424.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@163425.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wlast = fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@163361.4]
  assign MAGToAXI4Bridge_1_io_in_rresp_ready = fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 132:21:@163360.4]
  assign MAGToAXI4Bridge_1_io_in_wresp_ready = fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 132:21:@163341.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_AWREADY = io_M_AXI_1_AWREADY; // @[FringeZynq.scala 133:10:@163480.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_ARREADY = io_M_AXI_1_ARREADY; // @[FringeZynq.scala 133:10:@163468.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_WREADY = io_M_AXI_1_WREADY; // @[FringeZynq.scala 133:10:@163463.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BID = io_M_AXI_1_BID; // @[FringeZynq.scala 133:10:@163455.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BVALID = io_M_AXI_1_BVALID; // @[FringeZynq.scala 133:10:@163452.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_valid = fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 132:21:@163605.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_addr = fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 132:21:@163604.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_size = fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 132:21:@163603.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_isWr = fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@163601.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_tag = fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 132:21:@163600.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_valid = fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 132:21:@163598.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@163582.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@163583.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@163584.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@163585.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@163586.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@163587.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@163588.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@163589.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@163590.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@163591.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@163592.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@163593.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@163594.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@163595.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@163596.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@163597.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@163518.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@163519.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@163520.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@163521.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@163522.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@163523.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@163524.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@163525.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@163526.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@163527.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@163528.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@163529.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@163530.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@163531.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@163532.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@163533.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@163534.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@163535.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@163536.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@163537.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@163538.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@163539.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@163540.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@163541.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@163542.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@163543.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@163544.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@163545.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@163546.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@163547.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@163548.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@163549.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@163550.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@163551.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@163552.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@163553.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@163554.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@163555.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@163556.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@163557.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@163558.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@163559.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@163560.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@163561.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@163562.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@163563.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@163564.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@163565.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@163566.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@163567.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@163568.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@163569.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@163570.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@163571.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@163572.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@163573.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@163574.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@163575.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@163576.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@163577.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@163578.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@163579.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@163580.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@163581.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wlast = fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@163517.4]
  assign MAGToAXI4Bridge_2_io_in_rresp_ready = fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 132:21:@163516.4]
  assign MAGToAXI4Bridge_2_io_in_wresp_ready = fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 132:21:@163497.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_AWREADY = io_M_AXI_2_AWREADY; // @[FringeZynq.scala 133:10:@163636.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_ARREADY = io_M_AXI_2_ARREADY; // @[FringeZynq.scala 133:10:@163624.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_WREADY = io_M_AXI_2_WREADY; // @[FringeZynq.scala 133:10:@163619.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BID = io_M_AXI_2_BID; // @[FringeZynq.scala 133:10:@163611.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BVALID = io_M_AXI_2_BVALID; // @[FringeZynq.scala 133:10:@163608.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_valid = fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 132:21:@163761.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_addr = fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 132:21:@163760.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_size = fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 132:21:@163759.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_isWr = fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@163757.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_tag = fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 132:21:@163756.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_valid = fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 132:21:@163754.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@163738.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@163739.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@163740.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@163741.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@163742.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@163743.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@163744.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@163745.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@163746.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@163747.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@163748.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@163749.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@163750.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@163751.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@163752.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@163753.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@163674.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@163675.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@163676.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@163677.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@163678.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@163679.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@163680.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@163681.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@163682.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@163683.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@163684.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@163685.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@163686.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@163687.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@163688.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@163689.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@163690.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@163691.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@163692.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@163693.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@163694.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@163695.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@163696.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@163697.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@163698.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@163699.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@163700.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@163701.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@163702.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@163703.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@163704.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@163705.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@163706.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@163707.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@163708.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@163709.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@163710.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@163711.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@163712.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@163713.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@163714.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@163715.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@163716.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@163717.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@163718.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@163719.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@163720.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@163721.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@163722.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@163723.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@163724.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@163725.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@163726.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@163727.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@163728.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@163729.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@163730.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@163731.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@163732.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@163733.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@163734.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@163735.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@163736.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@163737.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wlast = fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@163673.4]
  assign MAGToAXI4Bridge_3_io_in_rresp_ready = fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 132:21:@163672.4]
  assign MAGToAXI4Bridge_3_io_in_wresp_ready = fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 132:21:@163653.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_AWREADY = io_M_AXI_3_AWREADY; // @[FringeZynq.scala 133:10:@163792.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_ARREADY = io_M_AXI_3_ARREADY; // @[FringeZynq.scala 133:10:@163780.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_WREADY = io_M_AXI_3_WREADY; // @[FringeZynq.scala 133:10:@163775.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BID = io_M_AXI_3_BID; // @[FringeZynq.scala 133:10:@163767.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BVALID = io_M_AXI_3_BVALID; // @[FringeZynq.scala 133:10:@163764.4]
endmodule
module SpatialIP( // @[:@163805.2]
  input          clock, // @[:@163806.4]
  input          reset, // @[:@163807.4]
  input          io_raddr, // @[:@163808.4]
  input          io_wen, // @[:@163808.4]
  input          io_waddr, // @[:@163808.4]
  input          io_wdata, // @[:@163808.4]
  output         io_rdata, // @[:@163808.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@163808.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@163808.4]
  input          io_S_AXI_AWVALID, // @[:@163808.4]
  output         io_S_AXI_AWREADY, // @[:@163808.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@163808.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@163808.4]
  input          io_S_AXI_ARVALID, // @[:@163808.4]
  output         io_S_AXI_ARREADY, // @[:@163808.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@163808.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@163808.4]
  input          io_S_AXI_WVALID, // @[:@163808.4]
  output         io_S_AXI_WREADY, // @[:@163808.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@163808.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@163808.4]
  output         io_S_AXI_RVALID, // @[:@163808.4]
  input          io_S_AXI_RREADY, // @[:@163808.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@163808.4]
  output         io_S_AXI_BVALID, // @[:@163808.4]
  input          io_S_AXI_BREADY, // @[:@163808.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@163808.4]
  output [31:0]  io_M_AXI_0_AWUSER, // @[:@163808.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@163808.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@163808.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@163808.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@163808.4]
  output         io_M_AXI_0_AWLOCK, // @[:@163808.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@163808.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@163808.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@163808.4]
  output         io_M_AXI_0_AWVALID, // @[:@163808.4]
  input          io_M_AXI_0_AWREADY, // @[:@163808.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@163808.4]
  output [31:0]  io_M_AXI_0_ARUSER, // @[:@163808.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@163808.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@163808.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@163808.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@163808.4]
  output         io_M_AXI_0_ARLOCK, // @[:@163808.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@163808.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@163808.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@163808.4]
  output         io_M_AXI_0_ARVALID, // @[:@163808.4]
  input          io_M_AXI_0_ARREADY, // @[:@163808.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@163808.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@163808.4]
  output         io_M_AXI_0_WLAST, // @[:@163808.4]
  output         io_M_AXI_0_WVALID, // @[:@163808.4]
  input          io_M_AXI_0_WREADY, // @[:@163808.4]
  input  [31:0]  io_M_AXI_0_RID, // @[:@163808.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@163808.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@163808.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@163808.4]
  input          io_M_AXI_0_RLAST, // @[:@163808.4]
  input          io_M_AXI_0_RVALID, // @[:@163808.4]
  output         io_M_AXI_0_RREADY, // @[:@163808.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@163808.4]
  input  [31:0]  io_M_AXI_0_BUSER, // @[:@163808.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@163808.4]
  input          io_M_AXI_0_BVALID, // @[:@163808.4]
  output         io_M_AXI_0_BREADY, // @[:@163808.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@163808.4]
  output [31:0]  io_M_AXI_1_AWUSER, // @[:@163808.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@163808.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@163808.4]
  output [2:0]   io_M_AXI_1_AWSIZE, // @[:@163808.4]
  output [1:0]   io_M_AXI_1_AWBURST, // @[:@163808.4]
  output         io_M_AXI_1_AWLOCK, // @[:@163808.4]
  output [3:0]   io_M_AXI_1_AWCACHE, // @[:@163808.4]
  output [2:0]   io_M_AXI_1_AWPROT, // @[:@163808.4]
  output [3:0]   io_M_AXI_1_AWQOS, // @[:@163808.4]
  output         io_M_AXI_1_AWVALID, // @[:@163808.4]
  input          io_M_AXI_1_AWREADY, // @[:@163808.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@163808.4]
  output [31:0]  io_M_AXI_1_ARUSER, // @[:@163808.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@163808.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@163808.4]
  output [2:0]   io_M_AXI_1_ARSIZE, // @[:@163808.4]
  output [1:0]   io_M_AXI_1_ARBURST, // @[:@163808.4]
  output         io_M_AXI_1_ARLOCK, // @[:@163808.4]
  output [3:0]   io_M_AXI_1_ARCACHE, // @[:@163808.4]
  output [2:0]   io_M_AXI_1_ARPROT, // @[:@163808.4]
  output [3:0]   io_M_AXI_1_ARQOS, // @[:@163808.4]
  output         io_M_AXI_1_ARVALID, // @[:@163808.4]
  input          io_M_AXI_1_ARREADY, // @[:@163808.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@163808.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@163808.4]
  output         io_M_AXI_1_WLAST, // @[:@163808.4]
  output         io_M_AXI_1_WVALID, // @[:@163808.4]
  input          io_M_AXI_1_WREADY, // @[:@163808.4]
  input  [31:0]  io_M_AXI_1_RID, // @[:@163808.4]
  input  [31:0]  io_M_AXI_1_RUSER, // @[:@163808.4]
  input  [511:0] io_M_AXI_1_RDATA, // @[:@163808.4]
  input  [1:0]   io_M_AXI_1_RRESP, // @[:@163808.4]
  input          io_M_AXI_1_RLAST, // @[:@163808.4]
  input          io_M_AXI_1_RVALID, // @[:@163808.4]
  output         io_M_AXI_1_RREADY, // @[:@163808.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@163808.4]
  input  [31:0]  io_M_AXI_1_BUSER, // @[:@163808.4]
  input  [1:0]   io_M_AXI_1_BRESP, // @[:@163808.4]
  input          io_M_AXI_1_BVALID, // @[:@163808.4]
  output         io_M_AXI_1_BREADY, // @[:@163808.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@163808.4]
  output [31:0]  io_M_AXI_2_AWUSER, // @[:@163808.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@163808.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@163808.4]
  output [2:0]   io_M_AXI_2_AWSIZE, // @[:@163808.4]
  output [1:0]   io_M_AXI_2_AWBURST, // @[:@163808.4]
  output         io_M_AXI_2_AWLOCK, // @[:@163808.4]
  output [3:0]   io_M_AXI_2_AWCACHE, // @[:@163808.4]
  output [2:0]   io_M_AXI_2_AWPROT, // @[:@163808.4]
  output [3:0]   io_M_AXI_2_AWQOS, // @[:@163808.4]
  output         io_M_AXI_2_AWVALID, // @[:@163808.4]
  input          io_M_AXI_2_AWREADY, // @[:@163808.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@163808.4]
  output [31:0]  io_M_AXI_2_ARUSER, // @[:@163808.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@163808.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@163808.4]
  output [2:0]   io_M_AXI_2_ARSIZE, // @[:@163808.4]
  output [1:0]   io_M_AXI_2_ARBURST, // @[:@163808.4]
  output         io_M_AXI_2_ARLOCK, // @[:@163808.4]
  output [3:0]   io_M_AXI_2_ARCACHE, // @[:@163808.4]
  output [2:0]   io_M_AXI_2_ARPROT, // @[:@163808.4]
  output [3:0]   io_M_AXI_2_ARQOS, // @[:@163808.4]
  output         io_M_AXI_2_ARVALID, // @[:@163808.4]
  input          io_M_AXI_2_ARREADY, // @[:@163808.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@163808.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@163808.4]
  output         io_M_AXI_2_WLAST, // @[:@163808.4]
  output         io_M_AXI_2_WVALID, // @[:@163808.4]
  input          io_M_AXI_2_WREADY, // @[:@163808.4]
  input  [31:0]  io_M_AXI_2_RID, // @[:@163808.4]
  input  [31:0]  io_M_AXI_2_RUSER, // @[:@163808.4]
  input  [511:0] io_M_AXI_2_RDATA, // @[:@163808.4]
  input  [1:0]   io_M_AXI_2_RRESP, // @[:@163808.4]
  input          io_M_AXI_2_RLAST, // @[:@163808.4]
  input          io_M_AXI_2_RVALID, // @[:@163808.4]
  output         io_M_AXI_2_RREADY, // @[:@163808.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@163808.4]
  input  [31:0]  io_M_AXI_2_BUSER, // @[:@163808.4]
  input  [1:0]   io_M_AXI_2_BRESP, // @[:@163808.4]
  input          io_M_AXI_2_BVALID, // @[:@163808.4]
  output         io_M_AXI_2_BREADY, // @[:@163808.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@163808.4]
  output [31:0]  io_M_AXI_3_AWUSER, // @[:@163808.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@163808.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@163808.4]
  output [2:0]   io_M_AXI_3_AWSIZE, // @[:@163808.4]
  output [1:0]   io_M_AXI_3_AWBURST, // @[:@163808.4]
  output         io_M_AXI_3_AWLOCK, // @[:@163808.4]
  output [3:0]   io_M_AXI_3_AWCACHE, // @[:@163808.4]
  output [2:0]   io_M_AXI_3_AWPROT, // @[:@163808.4]
  output [3:0]   io_M_AXI_3_AWQOS, // @[:@163808.4]
  output         io_M_AXI_3_AWVALID, // @[:@163808.4]
  input          io_M_AXI_3_AWREADY, // @[:@163808.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@163808.4]
  output [31:0]  io_M_AXI_3_ARUSER, // @[:@163808.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@163808.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@163808.4]
  output [2:0]   io_M_AXI_3_ARSIZE, // @[:@163808.4]
  output [1:0]   io_M_AXI_3_ARBURST, // @[:@163808.4]
  output         io_M_AXI_3_ARLOCK, // @[:@163808.4]
  output [3:0]   io_M_AXI_3_ARCACHE, // @[:@163808.4]
  output [2:0]   io_M_AXI_3_ARPROT, // @[:@163808.4]
  output [3:0]   io_M_AXI_3_ARQOS, // @[:@163808.4]
  output         io_M_AXI_3_ARVALID, // @[:@163808.4]
  input          io_M_AXI_3_ARREADY, // @[:@163808.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@163808.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@163808.4]
  output         io_M_AXI_3_WLAST, // @[:@163808.4]
  output         io_M_AXI_3_WVALID, // @[:@163808.4]
  input          io_M_AXI_3_WREADY, // @[:@163808.4]
  input  [31:0]  io_M_AXI_3_RID, // @[:@163808.4]
  input  [31:0]  io_M_AXI_3_RUSER, // @[:@163808.4]
  input  [511:0] io_M_AXI_3_RDATA, // @[:@163808.4]
  input  [1:0]   io_M_AXI_3_RRESP, // @[:@163808.4]
  input          io_M_AXI_3_RLAST, // @[:@163808.4]
  input          io_M_AXI_3_RVALID, // @[:@163808.4]
  output         io_M_AXI_3_RREADY, // @[:@163808.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@163808.4]
  input  [31:0]  io_M_AXI_3_BUSER, // @[:@163808.4]
  input  [1:0]   io_M_AXI_3_BRESP, // @[:@163808.4]
  input          io_M_AXI_3_BVALID, // @[:@163808.4]
  output         io_M_AXI_3_BREADY, // @[:@163808.4]
  input          io_TOP_AXI_AWID, // @[:@163808.4]
  input          io_TOP_AXI_AWUSER, // @[:@163808.4]
  input  [31:0]  io_TOP_AXI_AWADDR, // @[:@163808.4]
  input  [7:0]   io_TOP_AXI_AWLEN, // @[:@163808.4]
  input  [2:0]   io_TOP_AXI_AWSIZE, // @[:@163808.4]
  input  [1:0]   io_TOP_AXI_AWBURST, // @[:@163808.4]
  input          io_TOP_AXI_AWLOCK, // @[:@163808.4]
  input  [3:0]   io_TOP_AXI_AWCACHE, // @[:@163808.4]
  input  [2:0]   io_TOP_AXI_AWPROT, // @[:@163808.4]
  input  [3:0]   io_TOP_AXI_AWQOS, // @[:@163808.4]
  input          io_TOP_AXI_AWVALID, // @[:@163808.4]
  input          io_TOP_AXI_AWREADY, // @[:@163808.4]
  input          io_TOP_AXI_ARID, // @[:@163808.4]
  input          io_TOP_AXI_ARUSER, // @[:@163808.4]
  input  [31:0]  io_TOP_AXI_ARADDR, // @[:@163808.4]
  input  [7:0]   io_TOP_AXI_ARLEN, // @[:@163808.4]
  input  [2:0]   io_TOP_AXI_ARSIZE, // @[:@163808.4]
  input  [1:0]   io_TOP_AXI_ARBURST, // @[:@163808.4]
  input          io_TOP_AXI_ARLOCK, // @[:@163808.4]
  input  [3:0]   io_TOP_AXI_ARCACHE, // @[:@163808.4]
  input  [2:0]   io_TOP_AXI_ARPROT, // @[:@163808.4]
  input  [3:0]   io_TOP_AXI_ARQOS, // @[:@163808.4]
  input          io_TOP_AXI_ARVALID, // @[:@163808.4]
  input          io_TOP_AXI_ARREADY, // @[:@163808.4]
  input  [31:0]  io_TOP_AXI_WDATA, // @[:@163808.4]
  input  [63:0]  io_TOP_AXI_WSTRB, // @[:@163808.4]
  input          io_TOP_AXI_WLAST, // @[:@163808.4]
  input          io_TOP_AXI_WVALID, // @[:@163808.4]
  input          io_TOP_AXI_WREADY, // @[:@163808.4]
  input          io_TOP_AXI_RID, // @[:@163808.4]
  input          io_TOP_AXI_RUSER, // @[:@163808.4]
  input  [31:0]  io_TOP_AXI_RDATA, // @[:@163808.4]
  input  [1:0]   io_TOP_AXI_RRESP, // @[:@163808.4]
  input          io_TOP_AXI_RLAST, // @[:@163808.4]
  input          io_TOP_AXI_RVALID, // @[:@163808.4]
  input          io_TOP_AXI_RREADY, // @[:@163808.4]
  input          io_TOP_AXI_BID, // @[:@163808.4]
  input          io_TOP_AXI_BUSER, // @[:@163808.4]
  input  [1:0]   io_TOP_AXI_BRESP, // @[:@163808.4]
  input          io_TOP_AXI_BVALID, // @[:@163808.4]
  input          io_TOP_AXI_BREADY, // @[:@163808.4]
  input          io_DWIDTH_AXI_AWID, // @[:@163808.4]
  input          io_DWIDTH_AXI_AWUSER, // @[:@163808.4]
  input  [31:0]  io_DWIDTH_AXI_AWADDR, // @[:@163808.4]
  input  [7:0]   io_DWIDTH_AXI_AWLEN, // @[:@163808.4]
  input  [2:0]   io_DWIDTH_AXI_AWSIZE, // @[:@163808.4]
  input  [1:0]   io_DWIDTH_AXI_AWBURST, // @[:@163808.4]
  input          io_DWIDTH_AXI_AWLOCK, // @[:@163808.4]
  input  [3:0]   io_DWIDTH_AXI_AWCACHE, // @[:@163808.4]
  input  [2:0]   io_DWIDTH_AXI_AWPROT, // @[:@163808.4]
  input  [3:0]   io_DWIDTH_AXI_AWQOS, // @[:@163808.4]
  input          io_DWIDTH_AXI_AWVALID, // @[:@163808.4]
  input          io_DWIDTH_AXI_AWREADY, // @[:@163808.4]
  input          io_DWIDTH_AXI_ARID, // @[:@163808.4]
  input          io_DWIDTH_AXI_ARUSER, // @[:@163808.4]
  input  [31:0]  io_DWIDTH_AXI_ARADDR, // @[:@163808.4]
  input  [7:0]   io_DWIDTH_AXI_ARLEN, // @[:@163808.4]
  input  [2:0]   io_DWIDTH_AXI_ARSIZE, // @[:@163808.4]
  input  [1:0]   io_DWIDTH_AXI_ARBURST, // @[:@163808.4]
  input          io_DWIDTH_AXI_ARLOCK, // @[:@163808.4]
  input  [3:0]   io_DWIDTH_AXI_ARCACHE, // @[:@163808.4]
  input  [2:0]   io_DWIDTH_AXI_ARPROT, // @[:@163808.4]
  input  [3:0]   io_DWIDTH_AXI_ARQOS, // @[:@163808.4]
  input          io_DWIDTH_AXI_ARVALID, // @[:@163808.4]
  input          io_DWIDTH_AXI_ARREADY, // @[:@163808.4]
  input  [31:0]  io_DWIDTH_AXI_WDATA, // @[:@163808.4]
  input  [63:0]  io_DWIDTH_AXI_WSTRB, // @[:@163808.4]
  input          io_DWIDTH_AXI_WLAST, // @[:@163808.4]
  input          io_DWIDTH_AXI_WVALID, // @[:@163808.4]
  input          io_DWIDTH_AXI_WREADY, // @[:@163808.4]
  input          io_DWIDTH_AXI_RID, // @[:@163808.4]
  input          io_DWIDTH_AXI_RUSER, // @[:@163808.4]
  input  [31:0]  io_DWIDTH_AXI_RDATA, // @[:@163808.4]
  input  [1:0]   io_DWIDTH_AXI_RRESP, // @[:@163808.4]
  input          io_DWIDTH_AXI_RLAST, // @[:@163808.4]
  input          io_DWIDTH_AXI_RVALID, // @[:@163808.4]
  input          io_DWIDTH_AXI_RREADY, // @[:@163808.4]
  input          io_DWIDTH_AXI_BID, // @[:@163808.4]
  input          io_DWIDTH_AXI_BUSER, // @[:@163808.4]
  input  [1:0]   io_DWIDTH_AXI_BRESP, // @[:@163808.4]
  input          io_DWIDTH_AXI_BVALID, // @[:@163808.4]
  input          io_DWIDTH_AXI_BREADY, // @[:@163808.4]
  input          io_PROTOCOL_AXI_AWID, // @[:@163808.4]
  input          io_PROTOCOL_AXI_AWUSER, // @[:@163808.4]
  input  [31:0]  io_PROTOCOL_AXI_AWADDR, // @[:@163808.4]
  input  [7:0]   io_PROTOCOL_AXI_AWLEN, // @[:@163808.4]
  input  [2:0]   io_PROTOCOL_AXI_AWSIZE, // @[:@163808.4]
  input  [1:0]   io_PROTOCOL_AXI_AWBURST, // @[:@163808.4]
  input          io_PROTOCOL_AXI_AWLOCK, // @[:@163808.4]
  input  [3:0]   io_PROTOCOL_AXI_AWCACHE, // @[:@163808.4]
  input  [2:0]   io_PROTOCOL_AXI_AWPROT, // @[:@163808.4]
  input  [3:0]   io_PROTOCOL_AXI_AWQOS, // @[:@163808.4]
  input          io_PROTOCOL_AXI_AWVALID, // @[:@163808.4]
  input          io_PROTOCOL_AXI_AWREADY, // @[:@163808.4]
  input          io_PROTOCOL_AXI_ARID, // @[:@163808.4]
  input          io_PROTOCOL_AXI_ARUSER, // @[:@163808.4]
  input  [31:0]  io_PROTOCOL_AXI_ARADDR, // @[:@163808.4]
  input  [7:0]   io_PROTOCOL_AXI_ARLEN, // @[:@163808.4]
  input  [2:0]   io_PROTOCOL_AXI_ARSIZE, // @[:@163808.4]
  input  [1:0]   io_PROTOCOL_AXI_ARBURST, // @[:@163808.4]
  input          io_PROTOCOL_AXI_ARLOCK, // @[:@163808.4]
  input  [3:0]   io_PROTOCOL_AXI_ARCACHE, // @[:@163808.4]
  input  [2:0]   io_PROTOCOL_AXI_ARPROT, // @[:@163808.4]
  input  [3:0]   io_PROTOCOL_AXI_ARQOS, // @[:@163808.4]
  input          io_PROTOCOL_AXI_ARVALID, // @[:@163808.4]
  input          io_PROTOCOL_AXI_ARREADY, // @[:@163808.4]
  input  [31:0]  io_PROTOCOL_AXI_WDATA, // @[:@163808.4]
  input  [63:0]  io_PROTOCOL_AXI_WSTRB, // @[:@163808.4]
  input          io_PROTOCOL_AXI_WLAST, // @[:@163808.4]
  input          io_PROTOCOL_AXI_WVALID, // @[:@163808.4]
  input          io_PROTOCOL_AXI_WREADY, // @[:@163808.4]
  input          io_PROTOCOL_AXI_RID, // @[:@163808.4]
  input          io_PROTOCOL_AXI_RUSER, // @[:@163808.4]
  input  [31:0]  io_PROTOCOL_AXI_RDATA, // @[:@163808.4]
  input  [1:0]   io_PROTOCOL_AXI_RRESP, // @[:@163808.4]
  input          io_PROTOCOL_AXI_RLAST, // @[:@163808.4]
  input          io_PROTOCOL_AXI_RVALID, // @[:@163808.4]
  input          io_PROTOCOL_AXI_RREADY, // @[:@163808.4]
  input          io_PROTOCOL_AXI_BID, // @[:@163808.4]
  input          io_PROTOCOL_AXI_BUSER, // @[:@163808.4]
  input  [1:0]   io_PROTOCOL_AXI_BRESP, // @[:@163808.4]
  input          io_PROTOCOL_AXI_BVALID, // @[:@163808.4]
  input          io_PROTOCOL_AXI_BREADY, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_AWID, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_AWUSER, // @[:@163808.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_AWADDR, // @[:@163808.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_AWLEN, // @[:@163808.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWSIZE, // @[:@163808.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_AWBURST, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_AWLOCK, // @[:@163808.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWCACHE, // @[:@163808.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWPROT, // @[:@163808.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWQOS, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_AWVALID, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_AWREADY, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_ARID, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_ARUSER, // @[:@163808.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_ARADDR, // @[:@163808.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_ARLEN, // @[:@163808.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARSIZE, // @[:@163808.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_ARBURST, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_ARLOCK, // @[:@163808.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARCACHE, // @[:@163808.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARPROT, // @[:@163808.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARQOS, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_ARVALID, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_ARREADY, // @[:@163808.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_WDATA, // @[:@163808.4]
  input  [63:0]  io_CLOCKCONVERT_AXI_WSTRB, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_WLAST, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_WVALID, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_WREADY, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_RID, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_RUSER, // @[:@163808.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_RDATA, // @[:@163808.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_RRESP, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_RLAST, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_RVALID, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_RREADY, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_BID, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_BUSER, // @[:@163808.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_BRESP, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_BVALID, // @[:@163808.4]
  input          io_CLOCKCONVERT_AXI_BREADY // @[:@163808.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@163810.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@163810.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@163810.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@163810.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@163810.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@163810.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@163810.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@163810.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@163810.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@163810.4]
  wire  FringeZynq_clock; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_reset; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[Zynq.scala 18:24:@163952.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[Zynq.scala 18:24:@163952.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[Zynq.scala 18:24:@163952.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 18:24:@163952.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 18:24:@163952.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_0_AWREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 18:24:@163952.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_0_ARREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [511:0] FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 18:24:@163952.4]
  wire [63:0] FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_0_WREADY; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_0_BID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_0_BVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 18:24:@163952.4]
  wire [7:0] FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_1_AWREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 18:24:@163952.4]
  wire [7:0] FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_1_ARREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [511:0] FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 18:24:@163952.4]
  wire [63:0] FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_1_WREADY; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_1_BID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_1_BVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 18:24:@163952.4]
  wire [7:0] FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_2_AWREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 18:24:@163952.4]
  wire [7:0] FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_2_ARREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [511:0] FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 18:24:@163952.4]
  wire [63:0] FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_2_WREADY; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_2_BID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_2_BVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 18:24:@163952.4]
  wire [7:0] FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_3_AWREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 18:24:@163952.4]
  wire [7:0] FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_3_ARREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [511:0] FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 18:24:@163952.4]
  wire [63:0] FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_3_WREADY; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_M_AXI_3_BID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_3_BVALID; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_enable; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_done; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_reset; // @[Zynq.scala 18:24:@163952.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[Zynq.scala 18:24:@163952.4]
  wire [63:0] FringeZynq_io_argIns_1; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[Zynq.scala 18:24:@163952.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 18:24:@163952.4]
  wire [63:0] FringeZynq_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_memStreams_stores_0_data_valid; // @[Zynq.scala 18:24:@163952.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 18:24:@163952.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 18:24:@163952.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 18:24:@163952.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 18:24:@163952.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@163810.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  FringeZynq FringeZynq ( // @[Zynq.scala 18:24:@163952.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWID(FringeZynq_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeZynq_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_AWVALID(FringeZynq_io_M_AXI_0_AWVALID),
    .io_M_AXI_0_AWREADY(FringeZynq_io_M_AXI_0_AWREADY),
    .io_M_AXI_0_ARID(FringeZynq_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeZynq_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeZynq_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeZynq_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WDATA(FringeZynq_io_M_AXI_0_WDATA),
    .io_M_AXI_0_WSTRB(FringeZynq_io_M_AXI_0_WSTRB),
    .io_M_AXI_0_WLAST(FringeZynq_io_M_AXI_0_WLAST),
    .io_M_AXI_0_WVALID(FringeZynq_io_M_AXI_0_WVALID),
    .io_M_AXI_0_WREADY(FringeZynq_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RREADY(FringeZynq_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeZynq_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeZynq_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeZynq_io_M_AXI_0_BREADY),
    .io_M_AXI_1_AWID(FringeZynq_io_M_AXI_1_AWID),
    .io_M_AXI_1_AWADDR(FringeZynq_io_M_AXI_1_AWADDR),
    .io_M_AXI_1_AWLEN(FringeZynq_io_M_AXI_1_AWLEN),
    .io_M_AXI_1_AWVALID(FringeZynq_io_M_AXI_1_AWVALID),
    .io_M_AXI_1_AWREADY(FringeZynq_io_M_AXI_1_AWREADY),
    .io_M_AXI_1_ARID(FringeZynq_io_M_AXI_1_ARID),
    .io_M_AXI_1_ARADDR(FringeZynq_io_M_AXI_1_ARADDR),
    .io_M_AXI_1_ARLEN(FringeZynq_io_M_AXI_1_ARLEN),
    .io_M_AXI_1_ARVALID(FringeZynq_io_M_AXI_1_ARVALID),
    .io_M_AXI_1_ARREADY(FringeZynq_io_M_AXI_1_ARREADY),
    .io_M_AXI_1_WDATA(FringeZynq_io_M_AXI_1_WDATA),
    .io_M_AXI_1_WSTRB(FringeZynq_io_M_AXI_1_WSTRB),
    .io_M_AXI_1_WLAST(FringeZynq_io_M_AXI_1_WLAST),
    .io_M_AXI_1_WVALID(FringeZynq_io_M_AXI_1_WVALID),
    .io_M_AXI_1_WREADY(FringeZynq_io_M_AXI_1_WREADY),
    .io_M_AXI_1_RREADY(FringeZynq_io_M_AXI_1_RREADY),
    .io_M_AXI_1_BID(FringeZynq_io_M_AXI_1_BID),
    .io_M_AXI_1_BVALID(FringeZynq_io_M_AXI_1_BVALID),
    .io_M_AXI_1_BREADY(FringeZynq_io_M_AXI_1_BREADY),
    .io_M_AXI_2_AWID(FringeZynq_io_M_AXI_2_AWID),
    .io_M_AXI_2_AWADDR(FringeZynq_io_M_AXI_2_AWADDR),
    .io_M_AXI_2_AWLEN(FringeZynq_io_M_AXI_2_AWLEN),
    .io_M_AXI_2_AWVALID(FringeZynq_io_M_AXI_2_AWVALID),
    .io_M_AXI_2_AWREADY(FringeZynq_io_M_AXI_2_AWREADY),
    .io_M_AXI_2_ARID(FringeZynq_io_M_AXI_2_ARID),
    .io_M_AXI_2_ARADDR(FringeZynq_io_M_AXI_2_ARADDR),
    .io_M_AXI_2_ARLEN(FringeZynq_io_M_AXI_2_ARLEN),
    .io_M_AXI_2_ARVALID(FringeZynq_io_M_AXI_2_ARVALID),
    .io_M_AXI_2_ARREADY(FringeZynq_io_M_AXI_2_ARREADY),
    .io_M_AXI_2_WDATA(FringeZynq_io_M_AXI_2_WDATA),
    .io_M_AXI_2_WSTRB(FringeZynq_io_M_AXI_2_WSTRB),
    .io_M_AXI_2_WLAST(FringeZynq_io_M_AXI_2_WLAST),
    .io_M_AXI_2_WVALID(FringeZynq_io_M_AXI_2_WVALID),
    .io_M_AXI_2_WREADY(FringeZynq_io_M_AXI_2_WREADY),
    .io_M_AXI_2_RREADY(FringeZynq_io_M_AXI_2_RREADY),
    .io_M_AXI_2_BID(FringeZynq_io_M_AXI_2_BID),
    .io_M_AXI_2_BVALID(FringeZynq_io_M_AXI_2_BVALID),
    .io_M_AXI_2_BREADY(FringeZynq_io_M_AXI_2_BREADY),
    .io_M_AXI_3_AWID(FringeZynq_io_M_AXI_3_AWID),
    .io_M_AXI_3_AWADDR(FringeZynq_io_M_AXI_3_AWADDR),
    .io_M_AXI_3_AWLEN(FringeZynq_io_M_AXI_3_AWLEN),
    .io_M_AXI_3_AWVALID(FringeZynq_io_M_AXI_3_AWVALID),
    .io_M_AXI_3_AWREADY(FringeZynq_io_M_AXI_3_AWREADY),
    .io_M_AXI_3_ARID(FringeZynq_io_M_AXI_3_ARID),
    .io_M_AXI_3_ARADDR(FringeZynq_io_M_AXI_3_ARADDR),
    .io_M_AXI_3_ARLEN(FringeZynq_io_M_AXI_3_ARLEN),
    .io_M_AXI_3_ARVALID(FringeZynq_io_M_AXI_3_ARVALID),
    .io_M_AXI_3_ARREADY(FringeZynq_io_M_AXI_3_ARREADY),
    .io_M_AXI_3_WDATA(FringeZynq_io_M_AXI_3_WDATA),
    .io_M_AXI_3_WSTRB(FringeZynq_io_M_AXI_3_WSTRB),
    .io_M_AXI_3_WLAST(FringeZynq_io_M_AXI_3_WLAST),
    .io_M_AXI_3_WVALID(FringeZynq_io_M_AXI_3_WVALID),
    .io_M_AXI_3_WREADY(FringeZynq_io_M_AXI_3_WREADY),
    .io_M_AXI_3_RREADY(FringeZynq_io_M_AXI_3_RREADY),
    .io_M_AXI_3_BID(FringeZynq_io_M_AXI_3_BID),
    .io_M_AXI_3_BVALID(FringeZynq_io_M_AXI_3_BVALID),
    .io_M_AXI_3_BREADY(FringeZynq_io_M_AXI_3_BREADY),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argIns_1(FringeZynq_io_argIns_1),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(FringeZynq_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(FringeZynq_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(FringeZynq_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(FringeZynq_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(FringeZynq_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(FringeZynq_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(FringeZynq_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(FringeZynq_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(FringeZynq_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(FringeZynq_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(FringeZynq_io_memStreams_stores_0_wresp_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 21:21:@163970.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 21:21:@163966.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 21:21:@163962.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 21:21:@163961.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 21:21:@163960.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 21:21:@163959.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 21:21:@163957.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 21:21:@163956.4]
  assign io_M_AXI_0_AWID = FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 24:14:@164014.4]
  assign io_M_AXI_0_AWUSER = 32'h0; // @[Zynq.scala 24:14:@164013.4]
  assign io_M_AXI_0_AWADDR = FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 24:14:@164012.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 24:14:@164011.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@164010.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[Zynq.scala 24:14:@164009.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@164008.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@164007.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[Zynq.scala 24:14:@164006.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[Zynq.scala 24:14:@164005.4]
  assign io_M_AXI_0_AWVALID = FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 24:14:@164004.4]
  assign io_M_AXI_0_ARID = FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 24:14:@164002.4]
  assign io_M_AXI_0_ARUSER = 32'h0; // @[Zynq.scala 24:14:@164001.4]
  assign io_M_AXI_0_ARADDR = FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 24:14:@164000.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 24:14:@163999.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@163998.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[Zynq.scala 24:14:@163997.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@163996.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@163995.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[Zynq.scala 24:14:@163994.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[Zynq.scala 24:14:@163993.4]
  assign io_M_AXI_0_ARVALID = FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 24:14:@163992.4]
  assign io_M_AXI_0_WDATA = FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 24:14:@163990.4]
  assign io_M_AXI_0_WSTRB = FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 24:14:@163989.4]
  assign io_M_AXI_0_WLAST = FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 24:14:@163988.4]
  assign io_M_AXI_0_WVALID = FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 24:14:@163987.4]
  assign io_M_AXI_0_RREADY = FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 24:14:@163979.4]
  assign io_M_AXI_0_BREADY = FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 24:14:@163974.4]
  assign io_M_AXI_1_AWID = FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 24:14:@164055.4]
  assign io_M_AXI_1_AWUSER = 32'h0; // @[Zynq.scala 24:14:@164054.4]
  assign io_M_AXI_1_AWADDR = FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 24:14:@164053.4]
  assign io_M_AXI_1_AWLEN = FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 24:14:@164052.4]
  assign io_M_AXI_1_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@164051.4]
  assign io_M_AXI_1_AWBURST = 2'h1; // @[Zynq.scala 24:14:@164050.4]
  assign io_M_AXI_1_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@164049.4]
  assign io_M_AXI_1_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@164048.4]
  assign io_M_AXI_1_AWPROT = 3'h0; // @[Zynq.scala 24:14:@164047.4]
  assign io_M_AXI_1_AWQOS = 4'h0; // @[Zynq.scala 24:14:@164046.4]
  assign io_M_AXI_1_AWVALID = FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 24:14:@164045.4]
  assign io_M_AXI_1_ARID = FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 24:14:@164043.4]
  assign io_M_AXI_1_ARUSER = 32'h0; // @[Zynq.scala 24:14:@164042.4]
  assign io_M_AXI_1_ARADDR = FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 24:14:@164041.4]
  assign io_M_AXI_1_ARLEN = FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 24:14:@164040.4]
  assign io_M_AXI_1_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@164039.4]
  assign io_M_AXI_1_ARBURST = 2'h1; // @[Zynq.scala 24:14:@164038.4]
  assign io_M_AXI_1_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@164037.4]
  assign io_M_AXI_1_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@164036.4]
  assign io_M_AXI_1_ARPROT = 3'h0; // @[Zynq.scala 24:14:@164035.4]
  assign io_M_AXI_1_ARQOS = 4'h0; // @[Zynq.scala 24:14:@164034.4]
  assign io_M_AXI_1_ARVALID = FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 24:14:@164033.4]
  assign io_M_AXI_1_WDATA = FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 24:14:@164031.4]
  assign io_M_AXI_1_WSTRB = FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 24:14:@164030.4]
  assign io_M_AXI_1_WLAST = FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 24:14:@164029.4]
  assign io_M_AXI_1_WVALID = FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 24:14:@164028.4]
  assign io_M_AXI_1_RREADY = FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 24:14:@164020.4]
  assign io_M_AXI_1_BREADY = FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 24:14:@164015.4]
  assign io_M_AXI_2_AWID = FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 24:14:@164096.4]
  assign io_M_AXI_2_AWUSER = 32'h0; // @[Zynq.scala 24:14:@164095.4]
  assign io_M_AXI_2_AWADDR = FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 24:14:@164094.4]
  assign io_M_AXI_2_AWLEN = FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 24:14:@164093.4]
  assign io_M_AXI_2_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@164092.4]
  assign io_M_AXI_2_AWBURST = 2'h1; // @[Zynq.scala 24:14:@164091.4]
  assign io_M_AXI_2_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@164090.4]
  assign io_M_AXI_2_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@164089.4]
  assign io_M_AXI_2_AWPROT = 3'h0; // @[Zynq.scala 24:14:@164088.4]
  assign io_M_AXI_2_AWQOS = 4'h0; // @[Zynq.scala 24:14:@164087.4]
  assign io_M_AXI_2_AWVALID = FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 24:14:@164086.4]
  assign io_M_AXI_2_ARID = FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 24:14:@164084.4]
  assign io_M_AXI_2_ARUSER = 32'h0; // @[Zynq.scala 24:14:@164083.4]
  assign io_M_AXI_2_ARADDR = FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 24:14:@164082.4]
  assign io_M_AXI_2_ARLEN = FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 24:14:@164081.4]
  assign io_M_AXI_2_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@164080.4]
  assign io_M_AXI_2_ARBURST = 2'h1; // @[Zynq.scala 24:14:@164079.4]
  assign io_M_AXI_2_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@164078.4]
  assign io_M_AXI_2_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@164077.4]
  assign io_M_AXI_2_ARPROT = 3'h0; // @[Zynq.scala 24:14:@164076.4]
  assign io_M_AXI_2_ARQOS = 4'h0; // @[Zynq.scala 24:14:@164075.4]
  assign io_M_AXI_2_ARVALID = FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 24:14:@164074.4]
  assign io_M_AXI_2_WDATA = FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 24:14:@164072.4]
  assign io_M_AXI_2_WSTRB = FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 24:14:@164071.4]
  assign io_M_AXI_2_WLAST = FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 24:14:@164070.4]
  assign io_M_AXI_2_WVALID = FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 24:14:@164069.4]
  assign io_M_AXI_2_RREADY = FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 24:14:@164061.4]
  assign io_M_AXI_2_BREADY = FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 24:14:@164056.4]
  assign io_M_AXI_3_AWID = FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 24:14:@164137.4]
  assign io_M_AXI_3_AWUSER = 32'h0; // @[Zynq.scala 24:14:@164136.4]
  assign io_M_AXI_3_AWADDR = FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 24:14:@164135.4]
  assign io_M_AXI_3_AWLEN = FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 24:14:@164134.4]
  assign io_M_AXI_3_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@164133.4]
  assign io_M_AXI_3_AWBURST = 2'h1; // @[Zynq.scala 24:14:@164132.4]
  assign io_M_AXI_3_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@164131.4]
  assign io_M_AXI_3_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@164130.4]
  assign io_M_AXI_3_AWPROT = 3'h0; // @[Zynq.scala 24:14:@164129.4]
  assign io_M_AXI_3_AWQOS = 4'h0; // @[Zynq.scala 24:14:@164128.4]
  assign io_M_AXI_3_AWVALID = FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 24:14:@164127.4]
  assign io_M_AXI_3_ARID = FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 24:14:@164125.4]
  assign io_M_AXI_3_ARUSER = 32'h0; // @[Zynq.scala 24:14:@164124.4]
  assign io_M_AXI_3_ARADDR = FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 24:14:@164123.4]
  assign io_M_AXI_3_ARLEN = FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 24:14:@164122.4]
  assign io_M_AXI_3_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@164121.4]
  assign io_M_AXI_3_ARBURST = 2'h1; // @[Zynq.scala 24:14:@164120.4]
  assign io_M_AXI_3_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@164119.4]
  assign io_M_AXI_3_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@164118.4]
  assign io_M_AXI_3_ARPROT = 3'h0; // @[Zynq.scala 24:14:@164117.4]
  assign io_M_AXI_3_ARQOS = 4'h0; // @[Zynq.scala 24:14:@164116.4]
  assign io_M_AXI_3_ARVALID = FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 24:14:@164115.4]
  assign io_M_AXI_3_WDATA = FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 24:14:@164113.4]
  assign io_M_AXI_3_WSTRB = FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 24:14:@164112.4]
  assign io_M_AXI_3_WLAST = FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 24:14:@164111.4]
  assign io_M_AXI_3_WVALID = FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 24:14:@164110.4]
  assign io_M_AXI_3_RREADY = FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 24:14:@164102.4]
  assign io_M_AXI_3_BREADY = FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 24:14:@164097.4]
  assign accel_clock = clock; // @[:@163811.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@163812.4 Zynq.scala 54:17:@164426.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[Zynq.scala 51:21:@164421.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@164414.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@164409.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[Zynq.scala 49:26:@164393.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[Zynq.scala 49:26:@164394.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[Zynq.scala 49:26:@164395.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[Zynq.scala 49:26:@164396.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[Zynq.scala 49:26:@164397.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[Zynq.scala 49:26:@164398.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[Zynq.scala 49:26:@164399.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[Zynq.scala 49:26:@164400.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[Zynq.scala 49:26:@164401.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[Zynq.scala 49:26:@164402.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[Zynq.scala 49:26:@164403.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[Zynq.scala 49:26:@164404.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[Zynq.scala 49:26:@164405.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[Zynq.scala 49:26:@164406.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[Zynq.scala 49:26:@164407.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[Zynq.scala 49:26:@164408.4]
  assign accel_io_memStreams_stores_0_cmd_ready = FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 49:26:@164392.4]
  assign accel_io_memStreams_stores_0_data_ready = FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 49:26:@164388.4]
  assign accel_io_memStreams_stores_0_wresp_valid = FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 49:26:@164383.4]
  assign accel_io_memStreams_stores_0_wresp_bits = FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 49:26:@164382.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@164381.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@164362.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[Zynq.scala 49:26:@164346.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[Zynq.scala 49:26:@164347.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[Zynq.scala 49:26:@164348.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[Zynq.scala 49:26:@164349.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[Zynq.scala 49:26:@164350.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[Zynq.scala 49:26:@164351.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[Zynq.scala 49:26:@164352.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[Zynq.scala 49:26:@164353.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[Zynq.scala 49:26:@164354.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[Zynq.scala 49:26:@164355.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[Zynq.scala 49:26:@164356.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[Zynq.scala 49:26:@164357.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[Zynq.scala 49:26:@164358.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[Zynq.scala 49:26:@164359.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[Zynq.scala 49:26:@164360.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[Zynq.scala 49:26:@164361.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@164345.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[Zynq.scala 49:26:@164310.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[Zynq.scala 49:26:@164309.4]
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 50:20:@164417.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 50:20:@164416.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 50:20:@164415.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[Zynq.scala 34:21:@164303.4]
  assign accel_io_argIns_1 = FringeZynq_io_argIns_1; // @[Zynq.scala 34:21:@164304.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[Zynq.scala 40:24:@164307.4]
  assign FringeZynq_clock = clock; // @[:@163953.4]
  assign FringeZynq_reset = reset == 1'h0; // @[:@163954.4 Zynq.scala 53:18:@164425.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[Zynq.scala 21:21:@163973.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[Zynq.scala 21:21:@163972.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[Zynq.scala 21:21:@163971.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[Zynq.scala 21:21:@163969.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[Zynq.scala 21:21:@163968.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[Zynq.scala 21:21:@163967.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[Zynq.scala 21:21:@163965.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[Zynq.scala 21:21:@163964.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[Zynq.scala 21:21:@163963.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[Zynq.scala 21:21:@163958.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[Zynq.scala 21:21:@163955.4]
  assign FringeZynq_io_M_AXI_0_AWREADY = io_M_AXI_0_AWREADY; // @[Zynq.scala 24:14:@164003.4]
  assign FringeZynq_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY; // @[Zynq.scala 24:14:@163991.4]
  assign FringeZynq_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY; // @[Zynq.scala 24:14:@163986.4]
  assign FringeZynq_io_M_AXI_0_BID = io_M_AXI_0_BID; // @[Zynq.scala 24:14:@163978.4]
  assign FringeZynq_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID; // @[Zynq.scala 24:14:@163975.4]
  assign FringeZynq_io_M_AXI_1_AWREADY = io_M_AXI_1_AWREADY; // @[Zynq.scala 24:14:@164044.4]
  assign FringeZynq_io_M_AXI_1_ARREADY = io_M_AXI_1_ARREADY; // @[Zynq.scala 24:14:@164032.4]
  assign FringeZynq_io_M_AXI_1_WREADY = io_M_AXI_1_WREADY; // @[Zynq.scala 24:14:@164027.4]
  assign FringeZynq_io_M_AXI_1_BID = io_M_AXI_1_BID; // @[Zynq.scala 24:14:@164019.4]
  assign FringeZynq_io_M_AXI_1_BVALID = io_M_AXI_1_BVALID; // @[Zynq.scala 24:14:@164016.4]
  assign FringeZynq_io_M_AXI_2_AWREADY = io_M_AXI_2_AWREADY; // @[Zynq.scala 24:14:@164085.4]
  assign FringeZynq_io_M_AXI_2_ARREADY = io_M_AXI_2_ARREADY; // @[Zynq.scala 24:14:@164073.4]
  assign FringeZynq_io_M_AXI_2_WREADY = io_M_AXI_2_WREADY; // @[Zynq.scala 24:14:@164068.4]
  assign FringeZynq_io_M_AXI_2_BID = io_M_AXI_2_BID; // @[Zynq.scala 24:14:@164060.4]
  assign FringeZynq_io_M_AXI_2_BVALID = io_M_AXI_2_BVALID; // @[Zynq.scala 24:14:@164057.4]
  assign FringeZynq_io_M_AXI_3_AWREADY = io_M_AXI_3_AWREADY; // @[Zynq.scala 24:14:@164126.4]
  assign FringeZynq_io_M_AXI_3_ARREADY = io_M_AXI_3_ARREADY; // @[Zynq.scala 24:14:@164114.4]
  assign FringeZynq_io_M_AXI_3_WREADY = io_M_AXI_3_WREADY; // @[Zynq.scala 24:14:@164109.4]
  assign FringeZynq_io_M_AXI_3_BID = io_M_AXI_3_BID; // @[Zynq.scala 24:14:@164101.4]
  assign FringeZynq_io_M_AXI_3_BVALID = io_M_AXI_3_BVALID; // @[Zynq.scala 24:14:@164098.4]
  assign FringeZynq_io_done = accel_io_done; // @[Zynq.scala 52:20:@164422.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[Zynq.scala 37:26:@164306.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[Zynq.scala 36:25:@164305.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_valid = accel_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 49:26:@164391.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_addr = accel_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 49:26:@164390.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_size = accel_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 49:26:@164389.4]
  assign FringeZynq_io_memStreams_stores_0_data_valid = accel_io_memStreams_stores_0_data_valid; // @[Zynq.scala 49:26:@164387.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wdata_0 = accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 49:26:@164386.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wstrb = accel_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 49:26:@164385.4]
  assign FringeZynq_io_memStreams_stores_0_wresp_ready = accel_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 49:26:@164384.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[Zynq.scala 50:20:@164420.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 50:20:@164419.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 50:20:@164418.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module SRAMVerilogDualRead
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr0,
    input [AWIDTH-1:0] raddr1,
    input [AWIDTH-1:0] waddr,
    input raddrEn0,
    input raddrEn1,
    input waddrEn,
    input wen,
    input backpressure0,
    input backpressure1,
    input [DWIDTH-1:0] wdata,
    output reg [DWIDTH-1:0] rdata0,
    output reg [DWIDTH-1:0] rdata1
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk)
    begin
            if (wen)
            begin
                mem[waddr] <= wdata;
            end
            if (backpressure0) rdata0 <= mem[raddr0];
    end


    always @(posedge clk)
    begin
        if (backpressure1) rdata1 <= mem[raddr1];
    end
endmodule




