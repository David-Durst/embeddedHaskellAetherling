module FIFO(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  input  [15:0] I_3,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3
);
  reg [15:0] _T__0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [15:0] _T__1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg [15:0] _T__2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg [15:0] _T__3; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_4;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0 = _T__0; // @[FIFO.scala 14:7]
  assign O_1 = _T__1; // @[FIFO.scala 14:7]
  assign O_2 = _T__2; // @[FIFO.scala 14:7]
  assign O_3 = _T__3; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0 <= I_0;
    _T__1 <= I_1;
    _T__2 <= I_2;
    _T__3 <= I_3;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module NestedCounters(
  input   CE,
  output  valid
);
  assign valid = CE; // @[NestedCounters.scala 65:13]
endmodule
module NestedCounters_1(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 53:31]
  wire  NestedCounters_valid; // @[NestedCounters.scala 53:31]
  NestedCounters NestedCounters ( // @[NestedCounters.scala 53:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 56:11]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 57:22]
endmodule
module NestedCountersWithNumValid(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 20:44]
  wire  NestedCounters_valid; // @[NestedCounters.scala 20:44]
  NestedCounters_1 NestedCounters ( // @[NestedCounters.scala 20:44]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 22:9]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 21:27]
endmodule
module RAM_ST(
  input         clock,
  input         RE,
  input  [8:0]  RADDR,
  output [15:0] RDATA_0,
  output [15:0] RDATA_1,
  output [15:0] RDATA_2,
  output [15:0] RDATA_3,
  input         WE,
  input  [8:0]  WADDR,
  input  [15:0] WDATA_0,
  input  [15:0] WDATA_1,
  input  [15:0] WDATA_2,
  input  [15:0] WDATA_3
);
  wire  write_elem_counter_CE; // @[RAM_ST.scala 20:34]
  wire  write_elem_counter_valid; // @[RAM_ST.scala 20:34]
  wire  read_elem_counter_CE; // @[RAM_ST.scala 21:33]
  wire  read_elem_counter_valid; // @[RAM_ST.scala 21:33]
  reg [63:0] ram [0:479]; // @[RAM_ST.scala 29:24]
  reg [63:0] _RAND_0;
  wire [63:0] ram__T_11_data; // @[RAM_ST.scala 29:24]
  wire [8:0] ram__T_11_addr; // @[RAM_ST.scala 29:24]
  reg [63:0] _RAND_1;
  wire [63:0] ram__T_5_data; // @[RAM_ST.scala 29:24]
  wire [8:0] ram__T_5_addr; // @[RAM_ST.scala 29:24]
  wire  ram__T_5_mask; // @[RAM_ST.scala 29:24]
  wire  ram__T_5_en; // @[RAM_ST.scala 29:24]
  reg  ram__T_11_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [8:0] ram__T_11_addr_pipe_0;
  reg [31:0] _RAND_3;
  wire [8:0] _GEN_1; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_2; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_3; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_4; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_5; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_6; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_7; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_8; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_9; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_10; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_11; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_12; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_13; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_14; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_15; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_16; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_17; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_18; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_19; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_20; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_21; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_22; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_23; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_24; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_25; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_26; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_27; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_28; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_29; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_30; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_31; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_32; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_33; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_34; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_35; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_36; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_37; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_38; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_39; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_40; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_41; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_42; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_43; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_44; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_45; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_46; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_47; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_48; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_49; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_50; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_51; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_52; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_53; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_54; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_55; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_56; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_57; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_58; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_59; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_60; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_61; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_62; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_63; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_64; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_65; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_66; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_67; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_68; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_69; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_70; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_71; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_72; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_73; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_74; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_75; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_76; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_77; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_78; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_79; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_80; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_81; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_82; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_83; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_84; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_85; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_86; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_87; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_88; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_89; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_90; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_91; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_92; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_93; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_94; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_95; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_96; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_97; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_98; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_99; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_100; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_101; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_102; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_103; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_104; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_105; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_106; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_107; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_108; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_109; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_110; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_111; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_112; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_113; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_114; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_115; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_116; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_117; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_118; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_119; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_120; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_121; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_122; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_123; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_124; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_125; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_126; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_127; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_128; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_129; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_130; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_131; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_132; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_133; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_134; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_135; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_136; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_137; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_138; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_139; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_140; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_141; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_142; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_143; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_144; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_145; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_146; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_147; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_148; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_149; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_150; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_151; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_152; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_153; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_154; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_155; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_156; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_157; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_158; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_159; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_160; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_161; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_162; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_163; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_164; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_165; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_166; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_167; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_168; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_169; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_170; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_171; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_172; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_173; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_174; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_175; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_176; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_177; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_178; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_179; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_180; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_181; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_182; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_183; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_184; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_185; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_186; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_187; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_188; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_189; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_190; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_191; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_192; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_193; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_194; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_195; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_196; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_197; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_198; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_199; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_200; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_201; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_202; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_203; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_204; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_205; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_206; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_207; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_208; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_209; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_210; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_211; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_212; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_213; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_214; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_215; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_216; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_217; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_218; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_219; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_220; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_221; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_222; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_223; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_224; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_225; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_226; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_227; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_228; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_229; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_230; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_231; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_232; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_233; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_234; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_235; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_236; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_237; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_238; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_239; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_240; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_241; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_242; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_243; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_244; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_245; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_246; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_247; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_248; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_249; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_250; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_251; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_252; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_253; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_254; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_255; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_256; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_257; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_258; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_259; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_260; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_261; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_262; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_263; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_264; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_265; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_266; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_267; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_268; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_269; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_270; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_271; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_272; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_273; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_274; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_275; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_276; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_277; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_278; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_279; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_280; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_281; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_282; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_283; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_284; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_285; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_286; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_287; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_288; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_289; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_290; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_291; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_292; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_293; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_294; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_295; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_296; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_297; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_298; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_299; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_300; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_301; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_302; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_303; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_304; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_305; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_306; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_307; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_308; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_309; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_310; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_311; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_312; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_313; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_314; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_315; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_316; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_317; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_318; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_319; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_320; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_321; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_322; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_323; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_324; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_325; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_326; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_327; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_328; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_329; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_330; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_331; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_332; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_333; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_334; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_335; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_336; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_337; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_338; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_339; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_340; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_341; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_342; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_343; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_344; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_345; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_346; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_347; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_348; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_349; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_350; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_351; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_352; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_353; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_354; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_355; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_356; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_357; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_358; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_359; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_360; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_361; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_362; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_363; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_364; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_365; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_366; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_367; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_368; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_369; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_370; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_371; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_372; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_373; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_374; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_375; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_376; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_377; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_378; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_379; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_380; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_381; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_382; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_383; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_384; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_385; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_386; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_387; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_388; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_389; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_390; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_391; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_392; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_393; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_394; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_395; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_396; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_397; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_398; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_399; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_400; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_401; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_402; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_403; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_404; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_405; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_406; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_407; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_408; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_409; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_410; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_411; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_412; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_413; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_414; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_415; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_416; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_417; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_418; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_419; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_420; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_421; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_422; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_423; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_424; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_425; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_426; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_427; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_428; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_429; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_430; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_431; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_432; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_433; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_434; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_435; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_436; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_437; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_438; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_439; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_440; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_441; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_442; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_443; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_444; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_445; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_446; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_447; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_448; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_449; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_450; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_451; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_452; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_453; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_454; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_455; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_456; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_457; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_458; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_459; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_460; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_461; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_462; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_463; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_464; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_465; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_466; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_467; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_468; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_469; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_470; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_471; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_472; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_473; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_474; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_475; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_476; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_477; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_478; // @[RAM_ST.scala 31:71]
  wire [8:0] _GEN_479; // @[RAM_ST.scala 31:71]
  wire [9:0] _T; // @[RAM_ST.scala 31:71]
  wire [31:0] _T_2; // @[RAM_ST.scala 31:115]
  wire [31:0] _T_3; // @[RAM_ST.scala 31:115]
  wire [8:0] _GEN_486; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_487; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_488; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_489; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_490; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_491; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_492; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_493; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_494; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_495; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_496; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_497; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_498; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_499; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_500; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_501; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_502; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_503; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_504; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_505; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_506; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_507; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_508; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_509; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_510; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_511; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_512; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_513; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_514; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_515; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_516; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_517; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_518; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_519; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_520; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_521; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_522; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_523; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_524; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_525; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_526; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_527; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_528; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_529; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_530; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_531; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_532; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_533; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_534; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_535; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_536; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_537; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_538; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_539; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_540; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_541; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_542; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_543; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_544; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_545; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_546; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_547; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_548; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_549; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_550; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_551; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_552; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_553; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_554; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_555; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_556; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_557; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_558; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_559; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_560; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_561; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_562; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_563; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_564; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_565; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_566; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_567; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_568; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_569; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_570; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_571; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_572; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_573; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_574; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_575; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_576; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_577; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_578; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_579; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_580; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_581; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_582; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_583; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_584; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_585; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_586; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_587; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_588; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_589; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_590; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_591; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_592; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_593; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_594; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_595; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_596; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_597; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_598; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_599; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_600; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_601; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_602; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_603; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_604; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_605; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_606; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_607; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_608; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_609; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_610; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_611; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_612; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_613; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_614; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_615; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_616; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_617; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_618; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_619; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_620; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_621; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_622; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_623; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_624; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_625; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_626; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_627; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_628; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_629; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_630; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_631; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_632; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_633; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_634; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_635; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_636; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_637; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_638; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_639; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_640; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_641; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_642; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_643; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_644; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_645; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_646; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_647; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_648; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_649; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_650; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_651; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_652; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_653; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_654; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_655; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_656; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_657; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_658; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_659; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_660; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_661; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_662; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_663; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_664; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_665; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_666; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_667; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_668; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_669; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_670; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_671; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_672; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_673; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_674; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_675; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_676; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_677; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_678; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_679; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_680; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_681; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_682; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_683; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_684; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_685; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_686; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_687; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_688; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_689; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_690; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_691; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_692; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_693; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_694; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_695; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_696; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_697; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_698; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_699; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_700; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_701; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_702; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_703; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_704; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_705; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_706; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_707; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_708; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_709; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_710; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_711; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_712; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_713; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_714; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_715; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_716; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_717; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_718; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_719; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_720; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_721; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_722; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_723; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_724; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_725; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_726; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_727; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_728; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_729; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_730; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_731; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_732; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_733; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_734; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_735; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_736; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_737; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_738; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_739; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_740; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_741; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_742; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_743; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_744; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_745; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_746; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_747; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_748; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_749; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_750; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_751; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_752; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_753; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_754; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_755; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_756; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_757; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_758; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_759; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_760; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_761; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_762; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_763; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_764; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_765; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_766; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_767; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_768; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_769; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_770; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_771; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_772; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_773; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_774; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_775; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_776; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_777; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_778; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_779; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_780; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_781; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_782; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_783; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_784; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_785; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_786; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_787; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_788; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_789; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_790; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_791; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_792; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_793; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_794; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_795; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_796; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_797; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_798; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_799; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_800; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_801; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_802; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_803; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_804; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_805; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_806; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_807; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_808; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_809; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_810; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_811; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_812; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_813; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_814; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_815; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_816; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_817; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_818; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_819; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_820; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_821; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_822; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_823; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_824; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_825; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_826; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_827; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_828; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_829; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_830; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_831; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_832; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_833; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_834; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_835; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_836; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_837; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_838; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_839; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_840; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_841; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_842; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_843; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_844; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_845; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_846; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_847; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_848; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_849; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_850; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_851; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_852; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_853; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_854; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_855; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_856; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_857; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_858; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_859; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_860; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_861; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_862; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_863; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_864; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_865; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_866; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_867; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_868; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_869; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_870; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_871; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_872; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_873; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_874; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_875; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_876; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_877; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_878; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_879; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_880; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_881; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_882; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_883; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_884; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_885; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_886; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_887; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_888; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_889; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_890; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_891; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_892; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_893; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_894; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_895; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_896; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_897; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_898; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_899; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_900; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_901; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_902; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_903; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_904; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_905; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_906; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_907; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_908; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_909; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_910; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_911; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_912; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_913; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_914; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_915; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_916; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_917; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_918; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_919; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_920; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_921; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_922; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_923; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_924; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_925; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_926; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_927; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_928; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_929; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_930; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_931; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_932; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_933; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_934; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_935; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_936; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_937; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_938; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_939; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_940; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_941; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_942; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_943; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_944; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_945; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_946; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_947; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_948; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_949; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_950; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_951; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_952; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_953; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_954; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_955; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_956; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_957; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_958; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_959; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_960; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_961; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_962; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_963; // @[RAM_ST.scala 32:46]
  wire [8:0] _GEN_964; // @[RAM_ST.scala 32:46]
  wire [9:0] _T_6; // @[RAM_ST.scala 32:46]
  wire [63:0] _T_13;
  NestedCountersWithNumValid write_elem_counter ( // @[RAM_ST.scala 20:34]
    .CE(write_elem_counter_CE),
    .valid(write_elem_counter_valid)
  );
  NestedCountersWithNumValid read_elem_counter ( // @[RAM_ST.scala 21:33]
    .CE(read_elem_counter_CE),
    .valid(read_elem_counter_valid)
  );
  assign ram__T_11_addr = ram__T_11_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_11_data = ram[ram__T_11_addr]; // @[RAM_ST.scala 29:24]
  `else
  assign ram__T_11_data = ram__T_11_addr >= 9'h1e0 ? _RAND_1[63:0] : ram[ram__T_11_addr]; // @[RAM_ST.scala 29:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_5_data = {_T_3,_T_2};
  assign ram__T_5_addr = _T[8:0];
  assign ram__T_5_mask = 1'h1;
  assign ram__T_5_en = write_elem_counter_valid;
  assign _GEN_1 = 9'h1 == WADDR ? 9'h1 : 9'h0; // @[RAM_ST.scala 31:71]
  assign _GEN_2 = 9'h2 == WADDR ? 9'h2 : _GEN_1; // @[RAM_ST.scala 31:71]
  assign _GEN_3 = 9'h3 == WADDR ? 9'h3 : _GEN_2; // @[RAM_ST.scala 31:71]
  assign _GEN_4 = 9'h4 == WADDR ? 9'h4 : _GEN_3; // @[RAM_ST.scala 31:71]
  assign _GEN_5 = 9'h5 == WADDR ? 9'h5 : _GEN_4; // @[RAM_ST.scala 31:71]
  assign _GEN_6 = 9'h6 == WADDR ? 9'h6 : _GEN_5; // @[RAM_ST.scala 31:71]
  assign _GEN_7 = 9'h7 == WADDR ? 9'h7 : _GEN_6; // @[RAM_ST.scala 31:71]
  assign _GEN_8 = 9'h8 == WADDR ? 9'h8 : _GEN_7; // @[RAM_ST.scala 31:71]
  assign _GEN_9 = 9'h9 == WADDR ? 9'h9 : _GEN_8; // @[RAM_ST.scala 31:71]
  assign _GEN_10 = 9'ha == WADDR ? 9'ha : _GEN_9; // @[RAM_ST.scala 31:71]
  assign _GEN_11 = 9'hb == WADDR ? 9'hb : _GEN_10; // @[RAM_ST.scala 31:71]
  assign _GEN_12 = 9'hc == WADDR ? 9'hc : _GEN_11; // @[RAM_ST.scala 31:71]
  assign _GEN_13 = 9'hd == WADDR ? 9'hd : _GEN_12; // @[RAM_ST.scala 31:71]
  assign _GEN_14 = 9'he == WADDR ? 9'he : _GEN_13; // @[RAM_ST.scala 31:71]
  assign _GEN_15 = 9'hf == WADDR ? 9'hf : _GEN_14; // @[RAM_ST.scala 31:71]
  assign _GEN_16 = 9'h10 == WADDR ? 9'h10 : _GEN_15; // @[RAM_ST.scala 31:71]
  assign _GEN_17 = 9'h11 == WADDR ? 9'h11 : _GEN_16; // @[RAM_ST.scala 31:71]
  assign _GEN_18 = 9'h12 == WADDR ? 9'h12 : _GEN_17; // @[RAM_ST.scala 31:71]
  assign _GEN_19 = 9'h13 == WADDR ? 9'h13 : _GEN_18; // @[RAM_ST.scala 31:71]
  assign _GEN_20 = 9'h14 == WADDR ? 9'h14 : _GEN_19; // @[RAM_ST.scala 31:71]
  assign _GEN_21 = 9'h15 == WADDR ? 9'h15 : _GEN_20; // @[RAM_ST.scala 31:71]
  assign _GEN_22 = 9'h16 == WADDR ? 9'h16 : _GEN_21; // @[RAM_ST.scala 31:71]
  assign _GEN_23 = 9'h17 == WADDR ? 9'h17 : _GEN_22; // @[RAM_ST.scala 31:71]
  assign _GEN_24 = 9'h18 == WADDR ? 9'h18 : _GEN_23; // @[RAM_ST.scala 31:71]
  assign _GEN_25 = 9'h19 == WADDR ? 9'h19 : _GEN_24; // @[RAM_ST.scala 31:71]
  assign _GEN_26 = 9'h1a == WADDR ? 9'h1a : _GEN_25; // @[RAM_ST.scala 31:71]
  assign _GEN_27 = 9'h1b == WADDR ? 9'h1b : _GEN_26; // @[RAM_ST.scala 31:71]
  assign _GEN_28 = 9'h1c == WADDR ? 9'h1c : _GEN_27; // @[RAM_ST.scala 31:71]
  assign _GEN_29 = 9'h1d == WADDR ? 9'h1d : _GEN_28; // @[RAM_ST.scala 31:71]
  assign _GEN_30 = 9'h1e == WADDR ? 9'h1e : _GEN_29; // @[RAM_ST.scala 31:71]
  assign _GEN_31 = 9'h1f == WADDR ? 9'h1f : _GEN_30; // @[RAM_ST.scala 31:71]
  assign _GEN_32 = 9'h20 == WADDR ? 9'h20 : _GEN_31; // @[RAM_ST.scala 31:71]
  assign _GEN_33 = 9'h21 == WADDR ? 9'h21 : _GEN_32; // @[RAM_ST.scala 31:71]
  assign _GEN_34 = 9'h22 == WADDR ? 9'h22 : _GEN_33; // @[RAM_ST.scala 31:71]
  assign _GEN_35 = 9'h23 == WADDR ? 9'h23 : _GEN_34; // @[RAM_ST.scala 31:71]
  assign _GEN_36 = 9'h24 == WADDR ? 9'h24 : _GEN_35; // @[RAM_ST.scala 31:71]
  assign _GEN_37 = 9'h25 == WADDR ? 9'h25 : _GEN_36; // @[RAM_ST.scala 31:71]
  assign _GEN_38 = 9'h26 == WADDR ? 9'h26 : _GEN_37; // @[RAM_ST.scala 31:71]
  assign _GEN_39 = 9'h27 == WADDR ? 9'h27 : _GEN_38; // @[RAM_ST.scala 31:71]
  assign _GEN_40 = 9'h28 == WADDR ? 9'h28 : _GEN_39; // @[RAM_ST.scala 31:71]
  assign _GEN_41 = 9'h29 == WADDR ? 9'h29 : _GEN_40; // @[RAM_ST.scala 31:71]
  assign _GEN_42 = 9'h2a == WADDR ? 9'h2a : _GEN_41; // @[RAM_ST.scala 31:71]
  assign _GEN_43 = 9'h2b == WADDR ? 9'h2b : _GEN_42; // @[RAM_ST.scala 31:71]
  assign _GEN_44 = 9'h2c == WADDR ? 9'h2c : _GEN_43; // @[RAM_ST.scala 31:71]
  assign _GEN_45 = 9'h2d == WADDR ? 9'h2d : _GEN_44; // @[RAM_ST.scala 31:71]
  assign _GEN_46 = 9'h2e == WADDR ? 9'h2e : _GEN_45; // @[RAM_ST.scala 31:71]
  assign _GEN_47 = 9'h2f == WADDR ? 9'h2f : _GEN_46; // @[RAM_ST.scala 31:71]
  assign _GEN_48 = 9'h30 == WADDR ? 9'h30 : _GEN_47; // @[RAM_ST.scala 31:71]
  assign _GEN_49 = 9'h31 == WADDR ? 9'h31 : _GEN_48; // @[RAM_ST.scala 31:71]
  assign _GEN_50 = 9'h32 == WADDR ? 9'h32 : _GEN_49; // @[RAM_ST.scala 31:71]
  assign _GEN_51 = 9'h33 == WADDR ? 9'h33 : _GEN_50; // @[RAM_ST.scala 31:71]
  assign _GEN_52 = 9'h34 == WADDR ? 9'h34 : _GEN_51; // @[RAM_ST.scala 31:71]
  assign _GEN_53 = 9'h35 == WADDR ? 9'h35 : _GEN_52; // @[RAM_ST.scala 31:71]
  assign _GEN_54 = 9'h36 == WADDR ? 9'h36 : _GEN_53; // @[RAM_ST.scala 31:71]
  assign _GEN_55 = 9'h37 == WADDR ? 9'h37 : _GEN_54; // @[RAM_ST.scala 31:71]
  assign _GEN_56 = 9'h38 == WADDR ? 9'h38 : _GEN_55; // @[RAM_ST.scala 31:71]
  assign _GEN_57 = 9'h39 == WADDR ? 9'h39 : _GEN_56; // @[RAM_ST.scala 31:71]
  assign _GEN_58 = 9'h3a == WADDR ? 9'h3a : _GEN_57; // @[RAM_ST.scala 31:71]
  assign _GEN_59 = 9'h3b == WADDR ? 9'h3b : _GEN_58; // @[RAM_ST.scala 31:71]
  assign _GEN_60 = 9'h3c == WADDR ? 9'h3c : _GEN_59; // @[RAM_ST.scala 31:71]
  assign _GEN_61 = 9'h3d == WADDR ? 9'h3d : _GEN_60; // @[RAM_ST.scala 31:71]
  assign _GEN_62 = 9'h3e == WADDR ? 9'h3e : _GEN_61; // @[RAM_ST.scala 31:71]
  assign _GEN_63 = 9'h3f == WADDR ? 9'h3f : _GEN_62; // @[RAM_ST.scala 31:71]
  assign _GEN_64 = 9'h40 == WADDR ? 9'h40 : _GEN_63; // @[RAM_ST.scala 31:71]
  assign _GEN_65 = 9'h41 == WADDR ? 9'h41 : _GEN_64; // @[RAM_ST.scala 31:71]
  assign _GEN_66 = 9'h42 == WADDR ? 9'h42 : _GEN_65; // @[RAM_ST.scala 31:71]
  assign _GEN_67 = 9'h43 == WADDR ? 9'h43 : _GEN_66; // @[RAM_ST.scala 31:71]
  assign _GEN_68 = 9'h44 == WADDR ? 9'h44 : _GEN_67; // @[RAM_ST.scala 31:71]
  assign _GEN_69 = 9'h45 == WADDR ? 9'h45 : _GEN_68; // @[RAM_ST.scala 31:71]
  assign _GEN_70 = 9'h46 == WADDR ? 9'h46 : _GEN_69; // @[RAM_ST.scala 31:71]
  assign _GEN_71 = 9'h47 == WADDR ? 9'h47 : _GEN_70; // @[RAM_ST.scala 31:71]
  assign _GEN_72 = 9'h48 == WADDR ? 9'h48 : _GEN_71; // @[RAM_ST.scala 31:71]
  assign _GEN_73 = 9'h49 == WADDR ? 9'h49 : _GEN_72; // @[RAM_ST.scala 31:71]
  assign _GEN_74 = 9'h4a == WADDR ? 9'h4a : _GEN_73; // @[RAM_ST.scala 31:71]
  assign _GEN_75 = 9'h4b == WADDR ? 9'h4b : _GEN_74; // @[RAM_ST.scala 31:71]
  assign _GEN_76 = 9'h4c == WADDR ? 9'h4c : _GEN_75; // @[RAM_ST.scala 31:71]
  assign _GEN_77 = 9'h4d == WADDR ? 9'h4d : _GEN_76; // @[RAM_ST.scala 31:71]
  assign _GEN_78 = 9'h4e == WADDR ? 9'h4e : _GEN_77; // @[RAM_ST.scala 31:71]
  assign _GEN_79 = 9'h4f == WADDR ? 9'h4f : _GEN_78; // @[RAM_ST.scala 31:71]
  assign _GEN_80 = 9'h50 == WADDR ? 9'h50 : _GEN_79; // @[RAM_ST.scala 31:71]
  assign _GEN_81 = 9'h51 == WADDR ? 9'h51 : _GEN_80; // @[RAM_ST.scala 31:71]
  assign _GEN_82 = 9'h52 == WADDR ? 9'h52 : _GEN_81; // @[RAM_ST.scala 31:71]
  assign _GEN_83 = 9'h53 == WADDR ? 9'h53 : _GEN_82; // @[RAM_ST.scala 31:71]
  assign _GEN_84 = 9'h54 == WADDR ? 9'h54 : _GEN_83; // @[RAM_ST.scala 31:71]
  assign _GEN_85 = 9'h55 == WADDR ? 9'h55 : _GEN_84; // @[RAM_ST.scala 31:71]
  assign _GEN_86 = 9'h56 == WADDR ? 9'h56 : _GEN_85; // @[RAM_ST.scala 31:71]
  assign _GEN_87 = 9'h57 == WADDR ? 9'h57 : _GEN_86; // @[RAM_ST.scala 31:71]
  assign _GEN_88 = 9'h58 == WADDR ? 9'h58 : _GEN_87; // @[RAM_ST.scala 31:71]
  assign _GEN_89 = 9'h59 == WADDR ? 9'h59 : _GEN_88; // @[RAM_ST.scala 31:71]
  assign _GEN_90 = 9'h5a == WADDR ? 9'h5a : _GEN_89; // @[RAM_ST.scala 31:71]
  assign _GEN_91 = 9'h5b == WADDR ? 9'h5b : _GEN_90; // @[RAM_ST.scala 31:71]
  assign _GEN_92 = 9'h5c == WADDR ? 9'h5c : _GEN_91; // @[RAM_ST.scala 31:71]
  assign _GEN_93 = 9'h5d == WADDR ? 9'h5d : _GEN_92; // @[RAM_ST.scala 31:71]
  assign _GEN_94 = 9'h5e == WADDR ? 9'h5e : _GEN_93; // @[RAM_ST.scala 31:71]
  assign _GEN_95 = 9'h5f == WADDR ? 9'h5f : _GEN_94; // @[RAM_ST.scala 31:71]
  assign _GEN_96 = 9'h60 == WADDR ? 9'h60 : _GEN_95; // @[RAM_ST.scala 31:71]
  assign _GEN_97 = 9'h61 == WADDR ? 9'h61 : _GEN_96; // @[RAM_ST.scala 31:71]
  assign _GEN_98 = 9'h62 == WADDR ? 9'h62 : _GEN_97; // @[RAM_ST.scala 31:71]
  assign _GEN_99 = 9'h63 == WADDR ? 9'h63 : _GEN_98; // @[RAM_ST.scala 31:71]
  assign _GEN_100 = 9'h64 == WADDR ? 9'h64 : _GEN_99; // @[RAM_ST.scala 31:71]
  assign _GEN_101 = 9'h65 == WADDR ? 9'h65 : _GEN_100; // @[RAM_ST.scala 31:71]
  assign _GEN_102 = 9'h66 == WADDR ? 9'h66 : _GEN_101; // @[RAM_ST.scala 31:71]
  assign _GEN_103 = 9'h67 == WADDR ? 9'h67 : _GEN_102; // @[RAM_ST.scala 31:71]
  assign _GEN_104 = 9'h68 == WADDR ? 9'h68 : _GEN_103; // @[RAM_ST.scala 31:71]
  assign _GEN_105 = 9'h69 == WADDR ? 9'h69 : _GEN_104; // @[RAM_ST.scala 31:71]
  assign _GEN_106 = 9'h6a == WADDR ? 9'h6a : _GEN_105; // @[RAM_ST.scala 31:71]
  assign _GEN_107 = 9'h6b == WADDR ? 9'h6b : _GEN_106; // @[RAM_ST.scala 31:71]
  assign _GEN_108 = 9'h6c == WADDR ? 9'h6c : _GEN_107; // @[RAM_ST.scala 31:71]
  assign _GEN_109 = 9'h6d == WADDR ? 9'h6d : _GEN_108; // @[RAM_ST.scala 31:71]
  assign _GEN_110 = 9'h6e == WADDR ? 9'h6e : _GEN_109; // @[RAM_ST.scala 31:71]
  assign _GEN_111 = 9'h6f == WADDR ? 9'h6f : _GEN_110; // @[RAM_ST.scala 31:71]
  assign _GEN_112 = 9'h70 == WADDR ? 9'h70 : _GEN_111; // @[RAM_ST.scala 31:71]
  assign _GEN_113 = 9'h71 == WADDR ? 9'h71 : _GEN_112; // @[RAM_ST.scala 31:71]
  assign _GEN_114 = 9'h72 == WADDR ? 9'h72 : _GEN_113; // @[RAM_ST.scala 31:71]
  assign _GEN_115 = 9'h73 == WADDR ? 9'h73 : _GEN_114; // @[RAM_ST.scala 31:71]
  assign _GEN_116 = 9'h74 == WADDR ? 9'h74 : _GEN_115; // @[RAM_ST.scala 31:71]
  assign _GEN_117 = 9'h75 == WADDR ? 9'h75 : _GEN_116; // @[RAM_ST.scala 31:71]
  assign _GEN_118 = 9'h76 == WADDR ? 9'h76 : _GEN_117; // @[RAM_ST.scala 31:71]
  assign _GEN_119 = 9'h77 == WADDR ? 9'h77 : _GEN_118; // @[RAM_ST.scala 31:71]
  assign _GEN_120 = 9'h78 == WADDR ? 9'h78 : _GEN_119; // @[RAM_ST.scala 31:71]
  assign _GEN_121 = 9'h79 == WADDR ? 9'h79 : _GEN_120; // @[RAM_ST.scala 31:71]
  assign _GEN_122 = 9'h7a == WADDR ? 9'h7a : _GEN_121; // @[RAM_ST.scala 31:71]
  assign _GEN_123 = 9'h7b == WADDR ? 9'h7b : _GEN_122; // @[RAM_ST.scala 31:71]
  assign _GEN_124 = 9'h7c == WADDR ? 9'h7c : _GEN_123; // @[RAM_ST.scala 31:71]
  assign _GEN_125 = 9'h7d == WADDR ? 9'h7d : _GEN_124; // @[RAM_ST.scala 31:71]
  assign _GEN_126 = 9'h7e == WADDR ? 9'h7e : _GEN_125; // @[RAM_ST.scala 31:71]
  assign _GEN_127 = 9'h7f == WADDR ? 9'h7f : _GEN_126; // @[RAM_ST.scala 31:71]
  assign _GEN_128 = 9'h80 == WADDR ? 9'h80 : _GEN_127; // @[RAM_ST.scala 31:71]
  assign _GEN_129 = 9'h81 == WADDR ? 9'h81 : _GEN_128; // @[RAM_ST.scala 31:71]
  assign _GEN_130 = 9'h82 == WADDR ? 9'h82 : _GEN_129; // @[RAM_ST.scala 31:71]
  assign _GEN_131 = 9'h83 == WADDR ? 9'h83 : _GEN_130; // @[RAM_ST.scala 31:71]
  assign _GEN_132 = 9'h84 == WADDR ? 9'h84 : _GEN_131; // @[RAM_ST.scala 31:71]
  assign _GEN_133 = 9'h85 == WADDR ? 9'h85 : _GEN_132; // @[RAM_ST.scala 31:71]
  assign _GEN_134 = 9'h86 == WADDR ? 9'h86 : _GEN_133; // @[RAM_ST.scala 31:71]
  assign _GEN_135 = 9'h87 == WADDR ? 9'h87 : _GEN_134; // @[RAM_ST.scala 31:71]
  assign _GEN_136 = 9'h88 == WADDR ? 9'h88 : _GEN_135; // @[RAM_ST.scala 31:71]
  assign _GEN_137 = 9'h89 == WADDR ? 9'h89 : _GEN_136; // @[RAM_ST.scala 31:71]
  assign _GEN_138 = 9'h8a == WADDR ? 9'h8a : _GEN_137; // @[RAM_ST.scala 31:71]
  assign _GEN_139 = 9'h8b == WADDR ? 9'h8b : _GEN_138; // @[RAM_ST.scala 31:71]
  assign _GEN_140 = 9'h8c == WADDR ? 9'h8c : _GEN_139; // @[RAM_ST.scala 31:71]
  assign _GEN_141 = 9'h8d == WADDR ? 9'h8d : _GEN_140; // @[RAM_ST.scala 31:71]
  assign _GEN_142 = 9'h8e == WADDR ? 9'h8e : _GEN_141; // @[RAM_ST.scala 31:71]
  assign _GEN_143 = 9'h8f == WADDR ? 9'h8f : _GEN_142; // @[RAM_ST.scala 31:71]
  assign _GEN_144 = 9'h90 == WADDR ? 9'h90 : _GEN_143; // @[RAM_ST.scala 31:71]
  assign _GEN_145 = 9'h91 == WADDR ? 9'h91 : _GEN_144; // @[RAM_ST.scala 31:71]
  assign _GEN_146 = 9'h92 == WADDR ? 9'h92 : _GEN_145; // @[RAM_ST.scala 31:71]
  assign _GEN_147 = 9'h93 == WADDR ? 9'h93 : _GEN_146; // @[RAM_ST.scala 31:71]
  assign _GEN_148 = 9'h94 == WADDR ? 9'h94 : _GEN_147; // @[RAM_ST.scala 31:71]
  assign _GEN_149 = 9'h95 == WADDR ? 9'h95 : _GEN_148; // @[RAM_ST.scala 31:71]
  assign _GEN_150 = 9'h96 == WADDR ? 9'h96 : _GEN_149; // @[RAM_ST.scala 31:71]
  assign _GEN_151 = 9'h97 == WADDR ? 9'h97 : _GEN_150; // @[RAM_ST.scala 31:71]
  assign _GEN_152 = 9'h98 == WADDR ? 9'h98 : _GEN_151; // @[RAM_ST.scala 31:71]
  assign _GEN_153 = 9'h99 == WADDR ? 9'h99 : _GEN_152; // @[RAM_ST.scala 31:71]
  assign _GEN_154 = 9'h9a == WADDR ? 9'h9a : _GEN_153; // @[RAM_ST.scala 31:71]
  assign _GEN_155 = 9'h9b == WADDR ? 9'h9b : _GEN_154; // @[RAM_ST.scala 31:71]
  assign _GEN_156 = 9'h9c == WADDR ? 9'h9c : _GEN_155; // @[RAM_ST.scala 31:71]
  assign _GEN_157 = 9'h9d == WADDR ? 9'h9d : _GEN_156; // @[RAM_ST.scala 31:71]
  assign _GEN_158 = 9'h9e == WADDR ? 9'h9e : _GEN_157; // @[RAM_ST.scala 31:71]
  assign _GEN_159 = 9'h9f == WADDR ? 9'h9f : _GEN_158; // @[RAM_ST.scala 31:71]
  assign _GEN_160 = 9'ha0 == WADDR ? 9'ha0 : _GEN_159; // @[RAM_ST.scala 31:71]
  assign _GEN_161 = 9'ha1 == WADDR ? 9'ha1 : _GEN_160; // @[RAM_ST.scala 31:71]
  assign _GEN_162 = 9'ha2 == WADDR ? 9'ha2 : _GEN_161; // @[RAM_ST.scala 31:71]
  assign _GEN_163 = 9'ha3 == WADDR ? 9'ha3 : _GEN_162; // @[RAM_ST.scala 31:71]
  assign _GEN_164 = 9'ha4 == WADDR ? 9'ha4 : _GEN_163; // @[RAM_ST.scala 31:71]
  assign _GEN_165 = 9'ha5 == WADDR ? 9'ha5 : _GEN_164; // @[RAM_ST.scala 31:71]
  assign _GEN_166 = 9'ha6 == WADDR ? 9'ha6 : _GEN_165; // @[RAM_ST.scala 31:71]
  assign _GEN_167 = 9'ha7 == WADDR ? 9'ha7 : _GEN_166; // @[RAM_ST.scala 31:71]
  assign _GEN_168 = 9'ha8 == WADDR ? 9'ha8 : _GEN_167; // @[RAM_ST.scala 31:71]
  assign _GEN_169 = 9'ha9 == WADDR ? 9'ha9 : _GEN_168; // @[RAM_ST.scala 31:71]
  assign _GEN_170 = 9'haa == WADDR ? 9'haa : _GEN_169; // @[RAM_ST.scala 31:71]
  assign _GEN_171 = 9'hab == WADDR ? 9'hab : _GEN_170; // @[RAM_ST.scala 31:71]
  assign _GEN_172 = 9'hac == WADDR ? 9'hac : _GEN_171; // @[RAM_ST.scala 31:71]
  assign _GEN_173 = 9'had == WADDR ? 9'had : _GEN_172; // @[RAM_ST.scala 31:71]
  assign _GEN_174 = 9'hae == WADDR ? 9'hae : _GEN_173; // @[RAM_ST.scala 31:71]
  assign _GEN_175 = 9'haf == WADDR ? 9'haf : _GEN_174; // @[RAM_ST.scala 31:71]
  assign _GEN_176 = 9'hb0 == WADDR ? 9'hb0 : _GEN_175; // @[RAM_ST.scala 31:71]
  assign _GEN_177 = 9'hb1 == WADDR ? 9'hb1 : _GEN_176; // @[RAM_ST.scala 31:71]
  assign _GEN_178 = 9'hb2 == WADDR ? 9'hb2 : _GEN_177; // @[RAM_ST.scala 31:71]
  assign _GEN_179 = 9'hb3 == WADDR ? 9'hb3 : _GEN_178; // @[RAM_ST.scala 31:71]
  assign _GEN_180 = 9'hb4 == WADDR ? 9'hb4 : _GEN_179; // @[RAM_ST.scala 31:71]
  assign _GEN_181 = 9'hb5 == WADDR ? 9'hb5 : _GEN_180; // @[RAM_ST.scala 31:71]
  assign _GEN_182 = 9'hb6 == WADDR ? 9'hb6 : _GEN_181; // @[RAM_ST.scala 31:71]
  assign _GEN_183 = 9'hb7 == WADDR ? 9'hb7 : _GEN_182; // @[RAM_ST.scala 31:71]
  assign _GEN_184 = 9'hb8 == WADDR ? 9'hb8 : _GEN_183; // @[RAM_ST.scala 31:71]
  assign _GEN_185 = 9'hb9 == WADDR ? 9'hb9 : _GEN_184; // @[RAM_ST.scala 31:71]
  assign _GEN_186 = 9'hba == WADDR ? 9'hba : _GEN_185; // @[RAM_ST.scala 31:71]
  assign _GEN_187 = 9'hbb == WADDR ? 9'hbb : _GEN_186; // @[RAM_ST.scala 31:71]
  assign _GEN_188 = 9'hbc == WADDR ? 9'hbc : _GEN_187; // @[RAM_ST.scala 31:71]
  assign _GEN_189 = 9'hbd == WADDR ? 9'hbd : _GEN_188; // @[RAM_ST.scala 31:71]
  assign _GEN_190 = 9'hbe == WADDR ? 9'hbe : _GEN_189; // @[RAM_ST.scala 31:71]
  assign _GEN_191 = 9'hbf == WADDR ? 9'hbf : _GEN_190; // @[RAM_ST.scala 31:71]
  assign _GEN_192 = 9'hc0 == WADDR ? 9'hc0 : _GEN_191; // @[RAM_ST.scala 31:71]
  assign _GEN_193 = 9'hc1 == WADDR ? 9'hc1 : _GEN_192; // @[RAM_ST.scala 31:71]
  assign _GEN_194 = 9'hc2 == WADDR ? 9'hc2 : _GEN_193; // @[RAM_ST.scala 31:71]
  assign _GEN_195 = 9'hc3 == WADDR ? 9'hc3 : _GEN_194; // @[RAM_ST.scala 31:71]
  assign _GEN_196 = 9'hc4 == WADDR ? 9'hc4 : _GEN_195; // @[RAM_ST.scala 31:71]
  assign _GEN_197 = 9'hc5 == WADDR ? 9'hc5 : _GEN_196; // @[RAM_ST.scala 31:71]
  assign _GEN_198 = 9'hc6 == WADDR ? 9'hc6 : _GEN_197; // @[RAM_ST.scala 31:71]
  assign _GEN_199 = 9'hc7 == WADDR ? 9'hc7 : _GEN_198; // @[RAM_ST.scala 31:71]
  assign _GEN_200 = 9'hc8 == WADDR ? 9'hc8 : _GEN_199; // @[RAM_ST.scala 31:71]
  assign _GEN_201 = 9'hc9 == WADDR ? 9'hc9 : _GEN_200; // @[RAM_ST.scala 31:71]
  assign _GEN_202 = 9'hca == WADDR ? 9'hca : _GEN_201; // @[RAM_ST.scala 31:71]
  assign _GEN_203 = 9'hcb == WADDR ? 9'hcb : _GEN_202; // @[RAM_ST.scala 31:71]
  assign _GEN_204 = 9'hcc == WADDR ? 9'hcc : _GEN_203; // @[RAM_ST.scala 31:71]
  assign _GEN_205 = 9'hcd == WADDR ? 9'hcd : _GEN_204; // @[RAM_ST.scala 31:71]
  assign _GEN_206 = 9'hce == WADDR ? 9'hce : _GEN_205; // @[RAM_ST.scala 31:71]
  assign _GEN_207 = 9'hcf == WADDR ? 9'hcf : _GEN_206; // @[RAM_ST.scala 31:71]
  assign _GEN_208 = 9'hd0 == WADDR ? 9'hd0 : _GEN_207; // @[RAM_ST.scala 31:71]
  assign _GEN_209 = 9'hd1 == WADDR ? 9'hd1 : _GEN_208; // @[RAM_ST.scala 31:71]
  assign _GEN_210 = 9'hd2 == WADDR ? 9'hd2 : _GEN_209; // @[RAM_ST.scala 31:71]
  assign _GEN_211 = 9'hd3 == WADDR ? 9'hd3 : _GEN_210; // @[RAM_ST.scala 31:71]
  assign _GEN_212 = 9'hd4 == WADDR ? 9'hd4 : _GEN_211; // @[RAM_ST.scala 31:71]
  assign _GEN_213 = 9'hd5 == WADDR ? 9'hd5 : _GEN_212; // @[RAM_ST.scala 31:71]
  assign _GEN_214 = 9'hd6 == WADDR ? 9'hd6 : _GEN_213; // @[RAM_ST.scala 31:71]
  assign _GEN_215 = 9'hd7 == WADDR ? 9'hd7 : _GEN_214; // @[RAM_ST.scala 31:71]
  assign _GEN_216 = 9'hd8 == WADDR ? 9'hd8 : _GEN_215; // @[RAM_ST.scala 31:71]
  assign _GEN_217 = 9'hd9 == WADDR ? 9'hd9 : _GEN_216; // @[RAM_ST.scala 31:71]
  assign _GEN_218 = 9'hda == WADDR ? 9'hda : _GEN_217; // @[RAM_ST.scala 31:71]
  assign _GEN_219 = 9'hdb == WADDR ? 9'hdb : _GEN_218; // @[RAM_ST.scala 31:71]
  assign _GEN_220 = 9'hdc == WADDR ? 9'hdc : _GEN_219; // @[RAM_ST.scala 31:71]
  assign _GEN_221 = 9'hdd == WADDR ? 9'hdd : _GEN_220; // @[RAM_ST.scala 31:71]
  assign _GEN_222 = 9'hde == WADDR ? 9'hde : _GEN_221; // @[RAM_ST.scala 31:71]
  assign _GEN_223 = 9'hdf == WADDR ? 9'hdf : _GEN_222; // @[RAM_ST.scala 31:71]
  assign _GEN_224 = 9'he0 == WADDR ? 9'he0 : _GEN_223; // @[RAM_ST.scala 31:71]
  assign _GEN_225 = 9'he1 == WADDR ? 9'he1 : _GEN_224; // @[RAM_ST.scala 31:71]
  assign _GEN_226 = 9'he2 == WADDR ? 9'he2 : _GEN_225; // @[RAM_ST.scala 31:71]
  assign _GEN_227 = 9'he3 == WADDR ? 9'he3 : _GEN_226; // @[RAM_ST.scala 31:71]
  assign _GEN_228 = 9'he4 == WADDR ? 9'he4 : _GEN_227; // @[RAM_ST.scala 31:71]
  assign _GEN_229 = 9'he5 == WADDR ? 9'he5 : _GEN_228; // @[RAM_ST.scala 31:71]
  assign _GEN_230 = 9'he6 == WADDR ? 9'he6 : _GEN_229; // @[RAM_ST.scala 31:71]
  assign _GEN_231 = 9'he7 == WADDR ? 9'he7 : _GEN_230; // @[RAM_ST.scala 31:71]
  assign _GEN_232 = 9'he8 == WADDR ? 9'he8 : _GEN_231; // @[RAM_ST.scala 31:71]
  assign _GEN_233 = 9'he9 == WADDR ? 9'he9 : _GEN_232; // @[RAM_ST.scala 31:71]
  assign _GEN_234 = 9'hea == WADDR ? 9'hea : _GEN_233; // @[RAM_ST.scala 31:71]
  assign _GEN_235 = 9'heb == WADDR ? 9'heb : _GEN_234; // @[RAM_ST.scala 31:71]
  assign _GEN_236 = 9'hec == WADDR ? 9'hec : _GEN_235; // @[RAM_ST.scala 31:71]
  assign _GEN_237 = 9'hed == WADDR ? 9'hed : _GEN_236; // @[RAM_ST.scala 31:71]
  assign _GEN_238 = 9'hee == WADDR ? 9'hee : _GEN_237; // @[RAM_ST.scala 31:71]
  assign _GEN_239 = 9'hef == WADDR ? 9'hef : _GEN_238; // @[RAM_ST.scala 31:71]
  assign _GEN_240 = 9'hf0 == WADDR ? 9'hf0 : _GEN_239; // @[RAM_ST.scala 31:71]
  assign _GEN_241 = 9'hf1 == WADDR ? 9'hf1 : _GEN_240; // @[RAM_ST.scala 31:71]
  assign _GEN_242 = 9'hf2 == WADDR ? 9'hf2 : _GEN_241; // @[RAM_ST.scala 31:71]
  assign _GEN_243 = 9'hf3 == WADDR ? 9'hf3 : _GEN_242; // @[RAM_ST.scala 31:71]
  assign _GEN_244 = 9'hf4 == WADDR ? 9'hf4 : _GEN_243; // @[RAM_ST.scala 31:71]
  assign _GEN_245 = 9'hf5 == WADDR ? 9'hf5 : _GEN_244; // @[RAM_ST.scala 31:71]
  assign _GEN_246 = 9'hf6 == WADDR ? 9'hf6 : _GEN_245; // @[RAM_ST.scala 31:71]
  assign _GEN_247 = 9'hf7 == WADDR ? 9'hf7 : _GEN_246; // @[RAM_ST.scala 31:71]
  assign _GEN_248 = 9'hf8 == WADDR ? 9'hf8 : _GEN_247; // @[RAM_ST.scala 31:71]
  assign _GEN_249 = 9'hf9 == WADDR ? 9'hf9 : _GEN_248; // @[RAM_ST.scala 31:71]
  assign _GEN_250 = 9'hfa == WADDR ? 9'hfa : _GEN_249; // @[RAM_ST.scala 31:71]
  assign _GEN_251 = 9'hfb == WADDR ? 9'hfb : _GEN_250; // @[RAM_ST.scala 31:71]
  assign _GEN_252 = 9'hfc == WADDR ? 9'hfc : _GEN_251; // @[RAM_ST.scala 31:71]
  assign _GEN_253 = 9'hfd == WADDR ? 9'hfd : _GEN_252; // @[RAM_ST.scala 31:71]
  assign _GEN_254 = 9'hfe == WADDR ? 9'hfe : _GEN_253; // @[RAM_ST.scala 31:71]
  assign _GEN_255 = 9'hff == WADDR ? 9'hff : _GEN_254; // @[RAM_ST.scala 31:71]
  assign _GEN_256 = 9'h100 == WADDR ? 9'h100 : _GEN_255; // @[RAM_ST.scala 31:71]
  assign _GEN_257 = 9'h101 == WADDR ? 9'h101 : _GEN_256; // @[RAM_ST.scala 31:71]
  assign _GEN_258 = 9'h102 == WADDR ? 9'h102 : _GEN_257; // @[RAM_ST.scala 31:71]
  assign _GEN_259 = 9'h103 == WADDR ? 9'h103 : _GEN_258; // @[RAM_ST.scala 31:71]
  assign _GEN_260 = 9'h104 == WADDR ? 9'h104 : _GEN_259; // @[RAM_ST.scala 31:71]
  assign _GEN_261 = 9'h105 == WADDR ? 9'h105 : _GEN_260; // @[RAM_ST.scala 31:71]
  assign _GEN_262 = 9'h106 == WADDR ? 9'h106 : _GEN_261; // @[RAM_ST.scala 31:71]
  assign _GEN_263 = 9'h107 == WADDR ? 9'h107 : _GEN_262; // @[RAM_ST.scala 31:71]
  assign _GEN_264 = 9'h108 == WADDR ? 9'h108 : _GEN_263; // @[RAM_ST.scala 31:71]
  assign _GEN_265 = 9'h109 == WADDR ? 9'h109 : _GEN_264; // @[RAM_ST.scala 31:71]
  assign _GEN_266 = 9'h10a == WADDR ? 9'h10a : _GEN_265; // @[RAM_ST.scala 31:71]
  assign _GEN_267 = 9'h10b == WADDR ? 9'h10b : _GEN_266; // @[RAM_ST.scala 31:71]
  assign _GEN_268 = 9'h10c == WADDR ? 9'h10c : _GEN_267; // @[RAM_ST.scala 31:71]
  assign _GEN_269 = 9'h10d == WADDR ? 9'h10d : _GEN_268; // @[RAM_ST.scala 31:71]
  assign _GEN_270 = 9'h10e == WADDR ? 9'h10e : _GEN_269; // @[RAM_ST.scala 31:71]
  assign _GEN_271 = 9'h10f == WADDR ? 9'h10f : _GEN_270; // @[RAM_ST.scala 31:71]
  assign _GEN_272 = 9'h110 == WADDR ? 9'h110 : _GEN_271; // @[RAM_ST.scala 31:71]
  assign _GEN_273 = 9'h111 == WADDR ? 9'h111 : _GEN_272; // @[RAM_ST.scala 31:71]
  assign _GEN_274 = 9'h112 == WADDR ? 9'h112 : _GEN_273; // @[RAM_ST.scala 31:71]
  assign _GEN_275 = 9'h113 == WADDR ? 9'h113 : _GEN_274; // @[RAM_ST.scala 31:71]
  assign _GEN_276 = 9'h114 == WADDR ? 9'h114 : _GEN_275; // @[RAM_ST.scala 31:71]
  assign _GEN_277 = 9'h115 == WADDR ? 9'h115 : _GEN_276; // @[RAM_ST.scala 31:71]
  assign _GEN_278 = 9'h116 == WADDR ? 9'h116 : _GEN_277; // @[RAM_ST.scala 31:71]
  assign _GEN_279 = 9'h117 == WADDR ? 9'h117 : _GEN_278; // @[RAM_ST.scala 31:71]
  assign _GEN_280 = 9'h118 == WADDR ? 9'h118 : _GEN_279; // @[RAM_ST.scala 31:71]
  assign _GEN_281 = 9'h119 == WADDR ? 9'h119 : _GEN_280; // @[RAM_ST.scala 31:71]
  assign _GEN_282 = 9'h11a == WADDR ? 9'h11a : _GEN_281; // @[RAM_ST.scala 31:71]
  assign _GEN_283 = 9'h11b == WADDR ? 9'h11b : _GEN_282; // @[RAM_ST.scala 31:71]
  assign _GEN_284 = 9'h11c == WADDR ? 9'h11c : _GEN_283; // @[RAM_ST.scala 31:71]
  assign _GEN_285 = 9'h11d == WADDR ? 9'h11d : _GEN_284; // @[RAM_ST.scala 31:71]
  assign _GEN_286 = 9'h11e == WADDR ? 9'h11e : _GEN_285; // @[RAM_ST.scala 31:71]
  assign _GEN_287 = 9'h11f == WADDR ? 9'h11f : _GEN_286; // @[RAM_ST.scala 31:71]
  assign _GEN_288 = 9'h120 == WADDR ? 9'h120 : _GEN_287; // @[RAM_ST.scala 31:71]
  assign _GEN_289 = 9'h121 == WADDR ? 9'h121 : _GEN_288; // @[RAM_ST.scala 31:71]
  assign _GEN_290 = 9'h122 == WADDR ? 9'h122 : _GEN_289; // @[RAM_ST.scala 31:71]
  assign _GEN_291 = 9'h123 == WADDR ? 9'h123 : _GEN_290; // @[RAM_ST.scala 31:71]
  assign _GEN_292 = 9'h124 == WADDR ? 9'h124 : _GEN_291; // @[RAM_ST.scala 31:71]
  assign _GEN_293 = 9'h125 == WADDR ? 9'h125 : _GEN_292; // @[RAM_ST.scala 31:71]
  assign _GEN_294 = 9'h126 == WADDR ? 9'h126 : _GEN_293; // @[RAM_ST.scala 31:71]
  assign _GEN_295 = 9'h127 == WADDR ? 9'h127 : _GEN_294; // @[RAM_ST.scala 31:71]
  assign _GEN_296 = 9'h128 == WADDR ? 9'h128 : _GEN_295; // @[RAM_ST.scala 31:71]
  assign _GEN_297 = 9'h129 == WADDR ? 9'h129 : _GEN_296; // @[RAM_ST.scala 31:71]
  assign _GEN_298 = 9'h12a == WADDR ? 9'h12a : _GEN_297; // @[RAM_ST.scala 31:71]
  assign _GEN_299 = 9'h12b == WADDR ? 9'h12b : _GEN_298; // @[RAM_ST.scala 31:71]
  assign _GEN_300 = 9'h12c == WADDR ? 9'h12c : _GEN_299; // @[RAM_ST.scala 31:71]
  assign _GEN_301 = 9'h12d == WADDR ? 9'h12d : _GEN_300; // @[RAM_ST.scala 31:71]
  assign _GEN_302 = 9'h12e == WADDR ? 9'h12e : _GEN_301; // @[RAM_ST.scala 31:71]
  assign _GEN_303 = 9'h12f == WADDR ? 9'h12f : _GEN_302; // @[RAM_ST.scala 31:71]
  assign _GEN_304 = 9'h130 == WADDR ? 9'h130 : _GEN_303; // @[RAM_ST.scala 31:71]
  assign _GEN_305 = 9'h131 == WADDR ? 9'h131 : _GEN_304; // @[RAM_ST.scala 31:71]
  assign _GEN_306 = 9'h132 == WADDR ? 9'h132 : _GEN_305; // @[RAM_ST.scala 31:71]
  assign _GEN_307 = 9'h133 == WADDR ? 9'h133 : _GEN_306; // @[RAM_ST.scala 31:71]
  assign _GEN_308 = 9'h134 == WADDR ? 9'h134 : _GEN_307; // @[RAM_ST.scala 31:71]
  assign _GEN_309 = 9'h135 == WADDR ? 9'h135 : _GEN_308; // @[RAM_ST.scala 31:71]
  assign _GEN_310 = 9'h136 == WADDR ? 9'h136 : _GEN_309; // @[RAM_ST.scala 31:71]
  assign _GEN_311 = 9'h137 == WADDR ? 9'h137 : _GEN_310; // @[RAM_ST.scala 31:71]
  assign _GEN_312 = 9'h138 == WADDR ? 9'h138 : _GEN_311; // @[RAM_ST.scala 31:71]
  assign _GEN_313 = 9'h139 == WADDR ? 9'h139 : _GEN_312; // @[RAM_ST.scala 31:71]
  assign _GEN_314 = 9'h13a == WADDR ? 9'h13a : _GEN_313; // @[RAM_ST.scala 31:71]
  assign _GEN_315 = 9'h13b == WADDR ? 9'h13b : _GEN_314; // @[RAM_ST.scala 31:71]
  assign _GEN_316 = 9'h13c == WADDR ? 9'h13c : _GEN_315; // @[RAM_ST.scala 31:71]
  assign _GEN_317 = 9'h13d == WADDR ? 9'h13d : _GEN_316; // @[RAM_ST.scala 31:71]
  assign _GEN_318 = 9'h13e == WADDR ? 9'h13e : _GEN_317; // @[RAM_ST.scala 31:71]
  assign _GEN_319 = 9'h13f == WADDR ? 9'h13f : _GEN_318; // @[RAM_ST.scala 31:71]
  assign _GEN_320 = 9'h140 == WADDR ? 9'h140 : _GEN_319; // @[RAM_ST.scala 31:71]
  assign _GEN_321 = 9'h141 == WADDR ? 9'h141 : _GEN_320; // @[RAM_ST.scala 31:71]
  assign _GEN_322 = 9'h142 == WADDR ? 9'h142 : _GEN_321; // @[RAM_ST.scala 31:71]
  assign _GEN_323 = 9'h143 == WADDR ? 9'h143 : _GEN_322; // @[RAM_ST.scala 31:71]
  assign _GEN_324 = 9'h144 == WADDR ? 9'h144 : _GEN_323; // @[RAM_ST.scala 31:71]
  assign _GEN_325 = 9'h145 == WADDR ? 9'h145 : _GEN_324; // @[RAM_ST.scala 31:71]
  assign _GEN_326 = 9'h146 == WADDR ? 9'h146 : _GEN_325; // @[RAM_ST.scala 31:71]
  assign _GEN_327 = 9'h147 == WADDR ? 9'h147 : _GEN_326; // @[RAM_ST.scala 31:71]
  assign _GEN_328 = 9'h148 == WADDR ? 9'h148 : _GEN_327; // @[RAM_ST.scala 31:71]
  assign _GEN_329 = 9'h149 == WADDR ? 9'h149 : _GEN_328; // @[RAM_ST.scala 31:71]
  assign _GEN_330 = 9'h14a == WADDR ? 9'h14a : _GEN_329; // @[RAM_ST.scala 31:71]
  assign _GEN_331 = 9'h14b == WADDR ? 9'h14b : _GEN_330; // @[RAM_ST.scala 31:71]
  assign _GEN_332 = 9'h14c == WADDR ? 9'h14c : _GEN_331; // @[RAM_ST.scala 31:71]
  assign _GEN_333 = 9'h14d == WADDR ? 9'h14d : _GEN_332; // @[RAM_ST.scala 31:71]
  assign _GEN_334 = 9'h14e == WADDR ? 9'h14e : _GEN_333; // @[RAM_ST.scala 31:71]
  assign _GEN_335 = 9'h14f == WADDR ? 9'h14f : _GEN_334; // @[RAM_ST.scala 31:71]
  assign _GEN_336 = 9'h150 == WADDR ? 9'h150 : _GEN_335; // @[RAM_ST.scala 31:71]
  assign _GEN_337 = 9'h151 == WADDR ? 9'h151 : _GEN_336; // @[RAM_ST.scala 31:71]
  assign _GEN_338 = 9'h152 == WADDR ? 9'h152 : _GEN_337; // @[RAM_ST.scala 31:71]
  assign _GEN_339 = 9'h153 == WADDR ? 9'h153 : _GEN_338; // @[RAM_ST.scala 31:71]
  assign _GEN_340 = 9'h154 == WADDR ? 9'h154 : _GEN_339; // @[RAM_ST.scala 31:71]
  assign _GEN_341 = 9'h155 == WADDR ? 9'h155 : _GEN_340; // @[RAM_ST.scala 31:71]
  assign _GEN_342 = 9'h156 == WADDR ? 9'h156 : _GEN_341; // @[RAM_ST.scala 31:71]
  assign _GEN_343 = 9'h157 == WADDR ? 9'h157 : _GEN_342; // @[RAM_ST.scala 31:71]
  assign _GEN_344 = 9'h158 == WADDR ? 9'h158 : _GEN_343; // @[RAM_ST.scala 31:71]
  assign _GEN_345 = 9'h159 == WADDR ? 9'h159 : _GEN_344; // @[RAM_ST.scala 31:71]
  assign _GEN_346 = 9'h15a == WADDR ? 9'h15a : _GEN_345; // @[RAM_ST.scala 31:71]
  assign _GEN_347 = 9'h15b == WADDR ? 9'h15b : _GEN_346; // @[RAM_ST.scala 31:71]
  assign _GEN_348 = 9'h15c == WADDR ? 9'h15c : _GEN_347; // @[RAM_ST.scala 31:71]
  assign _GEN_349 = 9'h15d == WADDR ? 9'h15d : _GEN_348; // @[RAM_ST.scala 31:71]
  assign _GEN_350 = 9'h15e == WADDR ? 9'h15e : _GEN_349; // @[RAM_ST.scala 31:71]
  assign _GEN_351 = 9'h15f == WADDR ? 9'h15f : _GEN_350; // @[RAM_ST.scala 31:71]
  assign _GEN_352 = 9'h160 == WADDR ? 9'h160 : _GEN_351; // @[RAM_ST.scala 31:71]
  assign _GEN_353 = 9'h161 == WADDR ? 9'h161 : _GEN_352; // @[RAM_ST.scala 31:71]
  assign _GEN_354 = 9'h162 == WADDR ? 9'h162 : _GEN_353; // @[RAM_ST.scala 31:71]
  assign _GEN_355 = 9'h163 == WADDR ? 9'h163 : _GEN_354; // @[RAM_ST.scala 31:71]
  assign _GEN_356 = 9'h164 == WADDR ? 9'h164 : _GEN_355; // @[RAM_ST.scala 31:71]
  assign _GEN_357 = 9'h165 == WADDR ? 9'h165 : _GEN_356; // @[RAM_ST.scala 31:71]
  assign _GEN_358 = 9'h166 == WADDR ? 9'h166 : _GEN_357; // @[RAM_ST.scala 31:71]
  assign _GEN_359 = 9'h167 == WADDR ? 9'h167 : _GEN_358; // @[RAM_ST.scala 31:71]
  assign _GEN_360 = 9'h168 == WADDR ? 9'h168 : _GEN_359; // @[RAM_ST.scala 31:71]
  assign _GEN_361 = 9'h169 == WADDR ? 9'h169 : _GEN_360; // @[RAM_ST.scala 31:71]
  assign _GEN_362 = 9'h16a == WADDR ? 9'h16a : _GEN_361; // @[RAM_ST.scala 31:71]
  assign _GEN_363 = 9'h16b == WADDR ? 9'h16b : _GEN_362; // @[RAM_ST.scala 31:71]
  assign _GEN_364 = 9'h16c == WADDR ? 9'h16c : _GEN_363; // @[RAM_ST.scala 31:71]
  assign _GEN_365 = 9'h16d == WADDR ? 9'h16d : _GEN_364; // @[RAM_ST.scala 31:71]
  assign _GEN_366 = 9'h16e == WADDR ? 9'h16e : _GEN_365; // @[RAM_ST.scala 31:71]
  assign _GEN_367 = 9'h16f == WADDR ? 9'h16f : _GEN_366; // @[RAM_ST.scala 31:71]
  assign _GEN_368 = 9'h170 == WADDR ? 9'h170 : _GEN_367; // @[RAM_ST.scala 31:71]
  assign _GEN_369 = 9'h171 == WADDR ? 9'h171 : _GEN_368; // @[RAM_ST.scala 31:71]
  assign _GEN_370 = 9'h172 == WADDR ? 9'h172 : _GEN_369; // @[RAM_ST.scala 31:71]
  assign _GEN_371 = 9'h173 == WADDR ? 9'h173 : _GEN_370; // @[RAM_ST.scala 31:71]
  assign _GEN_372 = 9'h174 == WADDR ? 9'h174 : _GEN_371; // @[RAM_ST.scala 31:71]
  assign _GEN_373 = 9'h175 == WADDR ? 9'h175 : _GEN_372; // @[RAM_ST.scala 31:71]
  assign _GEN_374 = 9'h176 == WADDR ? 9'h176 : _GEN_373; // @[RAM_ST.scala 31:71]
  assign _GEN_375 = 9'h177 == WADDR ? 9'h177 : _GEN_374; // @[RAM_ST.scala 31:71]
  assign _GEN_376 = 9'h178 == WADDR ? 9'h178 : _GEN_375; // @[RAM_ST.scala 31:71]
  assign _GEN_377 = 9'h179 == WADDR ? 9'h179 : _GEN_376; // @[RAM_ST.scala 31:71]
  assign _GEN_378 = 9'h17a == WADDR ? 9'h17a : _GEN_377; // @[RAM_ST.scala 31:71]
  assign _GEN_379 = 9'h17b == WADDR ? 9'h17b : _GEN_378; // @[RAM_ST.scala 31:71]
  assign _GEN_380 = 9'h17c == WADDR ? 9'h17c : _GEN_379; // @[RAM_ST.scala 31:71]
  assign _GEN_381 = 9'h17d == WADDR ? 9'h17d : _GEN_380; // @[RAM_ST.scala 31:71]
  assign _GEN_382 = 9'h17e == WADDR ? 9'h17e : _GEN_381; // @[RAM_ST.scala 31:71]
  assign _GEN_383 = 9'h17f == WADDR ? 9'h17f : _GEN_382; // @[RAM_ST.scala 31:71]
  assign _GEN_384 = 9'h180 == WADDR ? 9'h180 : _GEN_383; // @[RAM_ST.scala 31:71]
  assign _GEN_385 = 9'h181 == WADDR ? 9'h181 : _GEN_384; // @[RAM_ST.scala 31:71]
  assign _GEN_386 = 9'h182 == WADDR ? 9'h182 : _GEN_385; // @[RAM_ST.scala 31:71]
  assign _GEN_387 = 9'h183 == WADDR ? 9'h183 : _GEN_386; // @[RAM_ST.scala 31:71]
  assign _GEN_388 = 9'h184 == WADDR ? 9'h184 : _GEN_387; // @[RAM_ST.scala 31:71]
  assign _GEN_389 = 9'h185 == WADDR ? 9'h185 : _GEN_388; // @[RAM_ST.scala 31:71]
  assign _GEN_390 = 9'h186 == WADDR ? 9'h186 : _GEN_389; // @[RAM_ST.scala 31:71]
  assign _GEN_391 = 9'h187 == WADDR ? 9'h187 : _GEN_390; // @[RAM_ST.scala 31:71]
  assign _GEN_392 = 9'h188 == WADDR ? 9'h188 : _GEN_391; // @[RAM_ST.scala 31:71]
  assign _GEN_393 = 9'h189 == WADDR ? 9'h189 : _GEN_392; // @[RAM_ST.scala 31:71]
  assign _GEN_394 = 9'h18a == WADDR ? 9'h18a : _GEN_393; // @[RAM_ST.scala 31:71]
  assign _GEN_395 = 9'h18b == WADDR ? 9'h18b : _GEN_394; // @[RAM_ST.scala 31:71]
  assign _GEN_396 = 9'h18c == WADDR ? 9'h18c : _GEN_395; // @[RAM_ST.scala 31:71]
  assign _GEN_397 = 9'h18d == WADDR ? 9'h18d : _GEN_396; // @[RAM_ST.scala 31:71]
  assign _GEN_398 = 9'h18e == WADDR ? 9'h18e : _GEN_397; // @[RAM_ST.scala 31:71]
  assign _GEN_399 = 9'h18f == WADDR ? 9'h18f : _GEN_398; // @[RAM_ST.scala 31:71]
  assign _GEN_400 = 9'h190 == WADDR ? 9'h190 : _GEN_399; // @[RAM_ST.scala 31:71]
  assign _GEN_401 = 9'h191 == WADDR ? 9'h191 : _GEN_400; // @[RAM_ST.scala 31:71]
  assign _GEN_402 = 9'h192 == WADDR ? 9'h192 : _GEN_401; // @[RAM_ST.scala 31:71]
  assign _GEN_403 = 9'h193 == WADDR ? 9'h193 : _GEN_402; // @[RAM_ST.scala 31:71]
  assign _GEN_404 = 9'h194 == WADDR ? 9'h194 : _GEN_403; // @[RAM_ST.scala 31:71]
  assign _GEN_405 = 9'h195 == WADDR ? 9'h195 : _GEN_404; // @[RAM_ST.scala 31:71]
  assign _GEN_406 = 9'h196 == WADDR ? 9'h196 : _GEN_405; // @[RAM_ST.scala 31:71]
  assign _GEN_407 = 9'h197 == WADDR ? 9'h197 : _GEN_406; // @[RAM_ST.scala 31:71]
  assign _GEN_408 = 9'h198 == WADDR ? 9'h198 : _GEN_407; // @[RAM_ST.scala 31:71]
  assign _GEN_409 = 9'h199 == WADDR ? 9'h199 : _GEN_408; // @[RAM_ST.scala 31:71]
  assign _GEN_410 = 9'h19a == WADDR ? 9'h19a : _GEN_409; // @[RAM_ST.scala 31:71]
  assign _GEN_411 = 9'h19b == WADDR ? 9'h19b : _GEN_410; // @[RAM_ST.scala 31:71]
  assign _GEN_412 = 9'h19c == WADDR ? 9'h19c : _GEN_411; // @[RAM_ST.scala 31:71]
  assign _GEN_413 = 9'h19d == WADDR ? 9'h19d : _GEN_412; // @[RAM_ST.scala 31:71]
  assign _GEN_414 = 9'h19e == WADDR ? 9'h19e : _GEN_413; // @[RAM_ST.scala 31:71]
  assign _GEN_415 = 9'h19f == WADDR ? 9'h19f : _GEN_414; // @[RAM_ST.scala 31:71]
  assign _GEN_416 = 9'h1a0 == WADDR ? 9'h1a0 : _GEN_415; // @[RAM_ST.scala 31:71]
  assign _GEN_417 = 9'h1a1 == WADDR ? 9'h1a1 : _GEN_416; // @[RAM_ST.scala 31:71]
  assign _GEN_418 = 9'h1a2 == WADDR ? 9'h1a2 : _GEN_417; // @[RAM_ST.scala 31:71]
  assign _GEN_419 = 9'h1a3 == WADDR ? 9'h1a3 : _GEN_418; // @[RAM_ST.scala 31:71]
  assign _GEN_420 = 9'h1a4 == WADDR ? 9'h1a4 : _GEN_419; // @[RAM_ST.scala 31:71]
  assign _GEN_421 = 9'h1a5 == WADDR ? 9'h1a5 : _GEN_420; // @[RAM_ST.scala 31:71]
  assign _GEN_422 = 9'h1a6 == WADDR ? 9'h1a6 : _GEN_421; // @[RAM_ST.scala 31:71]
  assign _GEN_423 = 9'h1a7 == WADDR ? 9'h1a7 : _GEN_422; // @[RAM_ST.scala 31:71]
  assign _GEN_424 = 9'h1a8 == WADDR ? 9'h1a8 : _GEN_423; // @[RAM_ST.scala 31:71]
  assign _GEN_425 = 9'h1a9 == WADDR ? 9'h1a9 : _GEN_424; // @[RAM_ST.scala 31:71]
  assign _GEN_426 = 9'h1aa == WADDR ? 9'h1aa : _GEN_425; // @[RAM_ST.scala 31:71]
  assign _GEN_427 = 9'h1ab == WADDR ? 9'h1ab : _GEN_426; // @[RAM_ST.scala 31:71]
  assign _GEN_428 = 9'h1ac == WADDR ? 9'h1ac : _GEN_427; // @[RAM_ST.scala 31:71]
  assign _GEN_429 = 9'h1ad == WADDR ? 9'h1ad : _GEN_428; // @[RAM_ST.scala 31:71]
  assign _GEN_430 = 9'h1ae == WADDR ? 9'h1ae : _GEN_429; // @[RAM_ST.scala 31:71]
  assign _GEN_431 = 9'h1af == WADDR ? 9'h1af : _GEN_430; // @[RAM_ST.scala 31:71]
  assign _GEN_432 = 9'h1b0 == WADDR ? 9'h1b0 : _GEN_431; // @[RAM_ST.scala 31:71]
  assign _GEN_433 = 9'h1b1 == WADDR ? 9'h1b1 : _GEN_432; // @[RAM_ST.scala 31:71]
  assign _GEN_434 = 9'h1b2 == WADDR ? 9'h1b2 : _GEN_433; // @[RAM_ST.scala 31:71]
  assign _GEN_435 = 9'h1b3 == WADDR ? 9'h1b3 : _GEN_434; // @[RAM_ST.scala 31:71]
  assign _GEN_436 = 9'h1b4 == WADDR ? 9'h1b4 : _GEN_435; // @[RAM_ST.scala 31:71]
  assign _GEN_437 = 9'h1b5 == WADDR ? 9'h1b5 : _GEN_436; // @[RAM_ST.scala 31:71]
  assign _GEN_438 = 9'h1b6 == WADDR ? 9'h1b6 : _GEN_437; // @[RAM_ST.scala 31:71]
  assign _GEN_439 = 9'h1b7 == WADDR ? 9'h1b7 : _GEN_438; // @[RAM_ST.scala 31:71]
  assign _GEN_440 = 9'h1b8 == WADDR ? 9'h1b8 : _GEN_439; // @[RAM_ST.scala 31:71]
  assign _GEN_441 = 9'h1b9 == WADDR ? 9'h1b9 : _GEN_440; // @[RAM_ST.scala 31:71]
  assign _GEN_442 = 9'h1ba == WADDR ? 9'h1ba : _GEN_441; // @[RAM_ST.scala 31:71]
  assign _GEN_443 = 9'h1bb == WADDR ? 9'h1bb : _GEN_442; // @[RAM_ST.scala 31:71]
  assign _GEN_444 = 9'h1bc == WADDR ? 9'h1bc : _GEN_443; // @[RAM_ST.scala 31:71]
  assign _GEN_445 = 9'h1bd == WADDR ? 9'h1bd : _GEN_444; // @[RAM_ST.scala 31:71]
  assign _GEN_446 = 9'h1be == WADDR ? 9'h1be : _GEN_445; // @[RAM_ST.scala 31:71]
  assign _GEN_447 = 9'h1bf == WADDR ? 9'h1bf : _GEN_446; // @[RAM_ST.scala 31:71]
  assign _GEN_448 = 9'h1c0 == WADDR ? 9'h1c0 : _GEN_447; // @[RAM_ST.scala 31:71]
  assign _GEN_449 = 9'h1c1 == WADDR ? 9'h1c1 : _GEN_448; // @[RAM_ST.scala 31:71]
  assign _GEN_450 = 9'h1c2 == WADDR ? 9'h1c2 : _GEN_449; // @[RAM_ST.scala 31:71]
  assign _GEN_451 = 9'h1c3 == WADDR ? 9'h1c3 : _GEN_450; // @[RAM_ST.scala 31:71]
  assign _GEN_452 = 9'h1c4 == WADDR ? 9'h1c4 : _GEN_451; // @[RAM_ST.scala 31:71]
  assign _GEN_453 = 9'h1c5 == WADDR ? 9'h1c5 : _GEN_452; // @[RAM_ST.scala 31:71]
  assign _GEN_454 = 9'h1c6 == WADDR ? 9'h1c6 : _GEN_453; // @[RAM_ST.scala 31:71]
  assign _GEN_455 = 9'h1c7 == WADDR ? 9'h1c7 : _GEN_454; // @[RAM_ST.scala 31:71]
  assign _GEN_456 = 9'h1c8 == WADDR ? 9'h1c8 : _GEN_455; // @[RAM_ST.scala 31:71]
  assign _GEN_457 = 9'h1c9 == WADDR ? 9'h1c9 : _GEN_456; // @[RAM_ST.scala 31:71]
  assign _GEN_458 = 9'h1ca == WADDR ? 9'h1ca : _GEN_457; // @[RAM_ST.scala 31:71]
  assign _GEN_459 = 9'h1cb == WADDR ? 9'h1cb : _GEN_458; // @[RAM_ST.scala 31:71]
  assign _GEN_460 = 9'h1cc == WADDR ? 9'h1cc : _GEN_459; // @[RAM_ST.scala 31:71]
  assign _GEN_461 = 9'h1cd == WADDR ? 9'h1cd : _GEN_460; // @[RAM_ST.scala 31:71]
  assign _GEN_462 = 9'h1ce == WADDR ? 9'h1ce : _GEN_461; // @[RAM_ST.scala 31:71]
  assign _GEN_463 = 9'h1cf == WADDR ? 9'h1cf : _GEN_462; // @[RAM_ST.scala 31:71]
  assign _GEN_464 = 9'h1d0 == WADDR ? 9'h1d0 : _GEN_463; // @[RAM_ST.scala 31:71]
  assign _GEN_465 = 9'h1d1 == WADDR ? 9'h1d1 : _GEN_464; // @[RAM_ST.scala 31:71]
  assign _GEN_466 = 9'h1d2 == WADDR ? 9'h1d2 : _GEN_465; // @[RAM_ST.scala 31:71]
  assign _GEN_467 = 9'h1d3 == WADDR ? 9'h1d3 : _GEN_466; // @[RAM_ST.scala 31:71]
  assign _GEN_468 = 9'h1d4 == WADDR ? 9'h1d4 : _GEN_467; // @[RAM_ST.scala 31:71]
  assign _GEN_469 = 9'h1d5 == WADDR ? 9'h1d5 : _GEN_468; // @[RAM_ST.scala 31:71]
  assign _GEN_470 = 9'h1d6 == WADDR ? 9'h1d6 : _GEN_469; // @[RAM_ST.scala 31:71]
  assign _GEN_471 = 9'h1d7 == WADDR ? 9'h1d7 : _GEN_470; // @[RAM_ST.scala 31:71]
  assign _GEN_472 = 9'h1d8 == WADDR ? 9'h1d8 : _GEN_471; // @[RAM_ST.scala 31:71]
  assign _GEN_473 = 9'h1d9 == WADDR ? 9'h1d9 : _GEN_472; // @[RAM_ST.scala 31:71]
  assign _GEN_474 = 9'h1da == WADDR ? 9'h1da : _GEN_473; // @[RAM_ST.scala 31:71]
  assign _GEN_475 = 9'h1db == WADDR ? 9'h1db : _GEN_474; // @[RAM_ST.scala 31:71]
  assign _GEN_476 = 9'h1dc == WADDR ? 9'h1dc : _GEN_475; // @[RAM_ST.scala 31:71]
  assign _GEN_477 = 9'h1dd == WADDR ? 9'h1dd : _GEN_476; // @[RAM_ST.scala 31:71]
  assign _GEN_478 = 9'h1de == WADDR ? 9'h1de : _GEN_477; // @[RAM_ST.scala 31:71]
  assign _GEN_479 = 9'h1df == WADDR ? 9'h1df : _GEN_478; // @[RAM_ST.scala 31:71]
  assign _T = {{1'd0}, _GEN_479}; // @[RAM_ST.scala 31:71]
  assign _T_2 = {WDATA_1,WDATA_0}; // @[RAM_ST.scala 31:115]
  assign _T_3 = {WDATA_3,WDATA_2}; // @[RAM_ST.scala 31:115]
  assign _GEN_486 = 9'h1 == RADDR ? 9'h1 : 9'h0; // @[RAM_ST.scala 32:46]
  assign _GEN_487 = 9'h2 == RADDR ? 9'h2 : _GEN_486; // @[RAM_ST.scala 32:46]
  assign _GEN_488 = 9'h3 == RADDR ? 9'h3 : _GEN_487; // @[RAM_ST.scala 32:46]
  assign _GEN_489 = 9'h4 == RADDR ? 9'h4 : _GEN_488; // @[RAM_ST.scala 32:46]
  assign _GEN_490 = 9'h5 == RADDR ? 9'h5 : _GEN_489; // @[RAM_ST.scala 32:46]
  assign _GEN_491 = 9'h6 == RADDR ? 9'h6 : _GEN_490; // @[RAM_ST.scala 32:46]
  assign _GEN_492 = 9'h7 == RADDR ? 9'h7 : _GEN_491; // @[RAM_ST.scala 32:46]
  assign _GEN_493 = 9'h8 == RADDR ? 9'h8 : _GEN_492; // @[RAM_ST.scala 32:46]
  assign _GEN_494 = 9'h9 == RADDR ? 9'h9 : _GEN_493; // @[RAM_ST.scala 32:46]
  assign _GEN_495 = 9'ha == RADDR ? 9'ha : _GEN_494; // @[RAM_ST.scala 32:46]
  assign _GEN_496 = 9'hb == RADDR ? 9'hb : _GEN_495; // @[RAM_ST.scala 32:46]
  assign _GEN_497 = 9'hc == RADDR ? 9'hc : _GEN_496; // @[RAM_ST.scala 32:46]
  assign _GEN_498 = 9'hd == RADDR ? 9'hd : _GEN_497; // @[RAM_ST.scala 32:46]
  assign _GEN_499 = 9'he == RADDR ? 9'he : _GEN_498; // @[RAM_ST.scala 32:46]
  assign _GEN_500 = 9'hf == RADDR ? 9'hf : _GEN_499; // @[RAM_ST.scala 32:46]
  assign _GEN_501 = 9'h10 == RADDR ? 9'h10 : _GEN_500; // @[RAM_ST.scala 32:46]
  assign _GEN_502 = 9'h11 == RADDR ? 9'h11 : _GEN_501; // @[RAM_ST.scala 32:46]
  assign _GEN_503 = 9'h12 == RADDR ? 9'h12 : _GEN_502; // @[RAM_ST.scala 32:46]
  assign _GEN_504 = 9'h13 == RADDR ? 9'h13 : _GEN_503; // @[RAM_ST.scala 32:46]
  assign _GEN_505 = 9'h14 == RADDR ? 9'h14 : _GEN_504; // @[RAM_ST.scala 32:46]
  assign _GEN_506 = 9'h15 == RADDR ? 9'h15 : _GEN_505; // @[RAM_ST.scala 32:46]
  assign _GEN_507 = 9'h16 == RADDR ? 9'h16 : _GEN_506; // @[RAM_ST.scala 32:46]
  assign _GEN_508 = 9'h17 == RADDR ? 9'h17 : _GEN_507; // @[RAM_ST.scala 32:46]
  assign _GEN_509 = 9'h18 == RADDR ? 9'h18 : _GEN_508; // @[RAM_ST.scala 32:46]
  assign _GEN_510 = 9'h19 == RADDR ? 9'h19 : _GEN_509; // @[RAM_ST.scala 32:46]
  assign _GEN_511 = 9'h1a == RADDR ? 9'h1a : _GEN_510; // @[RAM_ST.scala 32:46]
  assign _GEN_512 = 9'h1b == RADDR ? 9'h1b : _GEN_511; // @[RAM_ST.scala 32:46]
  assign _GEN_513 = 9'h1c == RADDR ? 9'h1c : _GEN_512; // @[RAM_ST.scala 32:46]
  assign _GEN_514 = 9'h1d == RADDR ? 9'h1d : _GEN_513; // @[RAM_ST.scala 32:46]
  assign _GEN_515 = 9'h1e == RADDR ? 9'h1e : _GEN_514; // @[RAM_ST.scala 32:46]
  assign _GEN_516 = 9'h1f == RADDR ? 9'h1f : _GEN_515; // @[RAM_ST.scala 32:46]
  assign _GEN_517 = 9'h20 == RADDR ? 9'h20 : _GEN_516; // @[RAM_ST.scala 32:46]
  assign _GEN_518 = 9'h21 == RADDR ? 9'h21 : _GEN_517; // @[RAM_ST.scala 32:46]
  assign _GEN_519 = 9'h22 == RADDR ? 9'h22 : _GEN_518; // @[RAM_ST.scala 32:46]
  assign _GEN_520 = 9'h23 == RADDR ? 9'h23 : _GEN_519; // @[RAM_ST.scala 32:46]
  assign _GEN_521 = 9'h24 == RADDR ? 9'h24 : _GEN_520; // @[RAM_ST.scala 32:46]
  assign _GEN_522 = 9'h25 == RADDR ? 9'h25 : _GEN_521; // @[RAM_ST.scala 32:46]
  assign _GEN_523 = 9'h26 == RADDR ? 9'h26 : _GEN_522; // @[RAM_ST.scala 32:46]
  assign _GEN_524 = 9'h27 == RADDR ? 9'h27 : _GEN_523; // @[RAM_ST.scala 32:46]
  assign _GEN_525 = 9'h28 == RADDR ? 9'h28 : _GEN_524; // @[RAM_ST.scala 32:46]
  assign _GEN_526 = 9'h29 == RADDR ? 9'h29 : _GEN_525; // @[RAM_ST.scala 32:46]
  assign _GEN_527 = 9'h2a == RADDR ? 9'h2a : _GEN_526; // @[RAM_ST.scala 32:46]
  assign _GEN_528 = 9'h2b == RADDR ? 9'h2b : _GEN_527; // @[RAM_ST.scala 32:46]
  assign _GEN_529 = 9'h2c == RADDR ? 9'h2c : _GEN_528; // @[RAM_ST.scala 32:46]
  assign _GEN_530 = 9'h2d == RADDR ? 9'h2d : _GEN_529; // @[RAM_ST.scala 32:46]
  assign _GEN_531 = 9'h2e == RADDR ? 9'h2e : _GEN_530; // @[RAM_ST.scala 32:46]
  assign _GEN_532 = 9'h2f == RADDR ? 9'h2f : _GEN_531; // @[RAM_ST.scala 32:46]
  assign _GEN_533 = 9'h30 == RADDR ? 9'h30 : _GEN_532; // @[RAM_ST.scala 32:46]
  assign _GEN_534 = 9'h31 == RADDR ? 9'h31 : _GEN_533; // @[RAM_ST.scala 32:46]
  assign _GEN_535 = 9'h32 == RADDR ? 9'h32 : _GEN_534; // @[RAM_ST.scala 32:46]
  assign _GEN_536 = 9'h33 == RADDR ? 9'h33 : _GEN_535; // @[RAM_ST.scala 32:46]
  assign _GEN_537 = 9'h34 == RADDR ? 9'h34 : _GEN_536; // @[RAM_ST.scala 32:46]
  assign _GEN_538 = 9'h35 == RADDR ? 9'h35 : _GEN_537; // @[RAM_ST.scala 32:46]
  assign _GEN_539 = 9'h36 == RADDR ? 9'h36 : _GEN_538; // @[RAM_ST.scala 32:46]
  assign _GEN_540 = 9'h37 == RADDR ? 9'h37 : _GEN_539; // @[RAM_ST.scala 32:46]
  assign _GEN_541 = 9'h38 == RADDR ? 9'h38 : _GEN_540; // @[RAM_ST.scala 32:46]
  assign _GEN_542 = 9'h39 == RADDR ? 9'h39 : _GEN_541; // @[RAM_ST.scala 32:46]
  assign _GEN_543 = 9'h3a == RADDR ? 9'h3a : _GEN_542; // @[RAM_ST.scala 32:46]
  assign _GEN_544 = 9'h3b == RADDR ? 9'h3b : _GEN_543; // @[RAM_ST.scala 32:46]
  assign _GEN_545 = 9'h3c == RADDR ? 9'h3c : _GEN_544; // @[RAM_ST.scala 32:46]
  assign _GEN_546 = 9'h3d == RADDR ? 9'h3d : _GEN_545; // @[RAM_ST.scala 32:46]
  assign _GEN_547 = 9'h3e == RADDR ? 9'h3e : _GEN_546; // @[RAM_ST.scala 32:46]
  assign _GEN_548 = 9'h3f == RADDR ? 9'h3f : _GEN_547; // @[RAM_ST.scala 32:46]
  assign _GEN_549 = 9'h40 == RADDR ? 9'h40 : _GEN_548; // @[RAM_ST.scala 32:46]
  assign _GEN_550 = 9'h41 == RADDR ? 9'h41 : _GEN_549; // @[RAM_ST.scala 32:46]
  assign _GEN_551 = 9'h42 == RADDR ? 9'h42 : _GEN_550; // @[RAM_ST.scala 32:46]
  assign _GEN_552 = 9'h43 == RADDR ? 9'h43 : _GEN_551; // @[RAM_ST.scala 32:46]
  assign _GEN_553 = 9'h44 == RADDR ? 9'h44 : _GEN_552; // @[RAM_ST.scala 32:46]
  assign _GEN_554 = 9'h45 == RADDR ? 9'h45 : _GEN_553; // @[RAM_ST.scala 32:46]
  assign _GEN_555 = 9'h46 == RADDR ? 9'h46 : _GEN_554; // @[RAM_ST.scala 32:46]
  assign _GEN_556 = 9'h47 == RADDR ? 9'h47 : _GEN_555; // @[RAM_ST.scala 32:46]
  assign _GEN_557 = 9'h48 == RADDR ? 9'h48 : _GEN_556; // @[RAM_ST.scala 32:46]
  assign _GEN_558 = 9'h49 == RADDR ? 9'h49 : _GEN_557; // @[RAM_ST.scala 32:46]
  assign _GEN_559 = 9'h4a == RADDR ? 9'h4a : _GEN_558; // @[RAM_ST.scala 32:46]
  assign _GEN_560 = 9'h4b == RADDR ? 9'h4b : _GEN_559; // @[RAM_ST.scala 32:46]
  assign _GEN_561 = 9'h4c == RADDR ? 9'h4c : _GEN_560; // @[RAM_ST.scala 32:46]
  assign _GEN_562 = 9'h4d == RADDR ? 9'h4d : _GEN_561; // @[RAM_ST.scala 32:46]
  assign _GEN_563 = 9'h4e == RADDR ? 9'h4e : _GEN_562; // @[RAM_ST.scala 32:46]
  assign _GEN_564 = 9'h4f == RADDR ? 9'h4f : _GEN_563; // @[RAM_ST.scala 32:46]
  assign _GEN_565 = 9'h50 == RADDR ? 9'h50 : _GEN_564; // @[RAM_ST.scala 32:46]
  assign _GEN_566 = 9'h51 == RADDR ? 9'h51 : _GEN_565; // @[RAM_ST.scala 32:46]
  assign _GEN_567 = 9'h52 == RADDR ? 9'h52 : _GEN_566; // @[RAM_ST.scala 32:46]
  assign _GEN_568 = 9'h53 == RADDR ? 9'h53 : _GEN_567; // @[RAM_ST.scala 32:46]
  assign _GEN_569 = 9'h54 == RADDR ? 9'h54 : _GEN_568; // @[RAM_ST.scala 32:46]
  assign _GEN_570 = 9'h55 == RADDR ? 9'h55 : _GEN_569; // @[RAM_ST.scala 32:46]
  assign _GEN_571 = 9'h56 == RADDR ? 9'h56 : _GEN_570; // @[RAM_ST.scala 32:46]
  assign _GEN_572 = 9'h57 == RADDR ? 9'h57 : _GEN_571; // @[RAM_ST.scala 32:46]
  assign _GEN_573 = 9'h58 == RADDR ? 9'h58 : _GEN_572; // @[RAM_ST.scala 32:46]
  assign _GEN_574 = 9'h59 == RADDR ? 9'h59 : _GEN_573; // @[RAM_ST.scala 32:46]
  assign _GEN_575 = 9'h5a == RADDR ? 9'h5a : _GEN_574; // @[RAM_ST.scala 32:46]
  assign _GEN_576 = 9'h5b == RADDR ? 9'h5b : _GEN_575; // @[RAM_ST.scala 32:46]
  assign _GEN_577 = 9'h5c == RADDR ? 9'h5c : _GEN_576; // @[RAM_ST.scala 32:46]
  assign _GEN_578 = 9'h5d == RADDR ? 9'h5d : _GEN_577; // @[RAM_ST.scala 32:46]
  assign _GEN_579 = 9'h5e == RADDR ? 9'h5e : _GEN_578; // @[RAM_ST.scala 32:46]
  assign _GEN_580 = 9'h5f == RADDR ? 9'h5f : _GEN_579; // @[RAM_ST.scala 32:46]
  assign _GEN_581 = 9'h60 == RADDR ? 9'h60 : _GEN_580; // @[RAM_ST.scala 32:46]
  assign _GEN_582 = 9'h61 == RADDR ? 9'h61 : _GEN_581; // @[RAM_ST.scala 32:46]
  assign _GEN_583 = 9'h62 == RADDR ? 9'h62 : _GEN_582; // @[RAM_ST.scala 32:46]
  assign _GEN_584 = 9'h63 == RADDR ? 9'h63 : _GEN_583; // @[RAM_ST.scala 32:46]
  assign _GEN_585 = 9'h64 == RADDR ? 9'h64 : _GEN_584; // @[RAM_ST.scala 32:46]
  assign _GEN_586 = 9'h65 == RADDR ? 9'h65 : _GEN_585; // @[RAM_ST.scala 32:46]
  assign _GEN_587 = 9'h66 == RADDR ? 9'h66 : _GEN_586; // @[RAM_ST.scala 32:46]
  assign _GEN_588 = 9'h67 == RADDR ? 9'h67 : _GEN_587; // @[RAM_ST.scala 32:46]
  assign _GEN_589 = 9'h68 == RADDR ? 9'h68 : _GEN_588; // @[RAM_ST.scala 32:46]
  assign _GEN_590 = 9'h69 == RADDR ? 9'h69 : _GEN_589; // @[RAM_ST.scala 32:46]
  assign _GEN_591 = 9'h6a == RADDR ? 9'h6a : _GEN_590; // @[RAM_ST.scala 32:46]
  assign _GEN_592 = 9'h6b == RADDR ? 9'h6b : _GEN_591; // @[RAM_ST.scala 32:46]
  assign _GEN_593 = 9'h6c == RADDR ? 9'h6c : _GEN_592; // @[RAM_ST.scala 32:46]
  assign _GEN_594 = 9'h6d == RADDR ? 9'h6d : _GEN_593; // @[RAM_ST.scala 32:46]
  assign _GEN_595 = 9'h6e == RADDR ? 9'h6e : _GEN_594; // @[RAM_ST.scala 32:46]
  assign _GEN_596 = 9'h6f == RADDR ? 9'h6f : _GEN_595; // @[RAM_ST.scala 32:46]
  assign _GEN_597 = 9'h70 == RADDR ? 9'h70 : _GEN_596; // @[RAM_ST.scala 32:46]
  assign _GEN_598 = 9'h71 == RADDR ? 9'h71 : _GEN_597; // @[RAM_ST.scala 32:46]
  assign _GEN_599 = 9'h72 == RADDR ? 9'h72 : _GEN_598; // @[RAM_ST.scala 32:46]
  assign _GEN_600 = 9'h73 == RADDR ? 9'h73 : _GEN_599; // @[RAM_ST.scala 32:46]
  assign _GEN_601 = 9'h74 == RADDR ? 9'h74 : _GEN_600; // @[RAM_ST.scala 32:46]
  assign _GEN_602 = 9'h75 == RADDR ? 9'h75 : _GEN_601; // @[RAM_ST.scala 32:46]
  assign _GEN_603 = 9'h76 == RADDR ? 9'h76 : _GEN_602; // @[RAM_ST.scala 32:46]
  assign _GEN_604 = 9'h77 == RADDR ? 9'h77 : _GEN_603; // @[RAM_ST.scala 32:46]
  assign _GEN_605 = 9'h78 == RADDR ? 9'h78 : _GEN_604; // @[RAM_ST.scala 32:46]
  assign _GEN_606 = 9'h79 == RADDR ? 9'h79 : _GEN_605; // @[RAM_ST.scala 32:46]
  assign _GEN_607 = 9'h7a == RADDR ? 9'h7a : _GEN_606; // @[RAM_ST.scala 32:46]
  assign _GEN_608 = 9'h7b == RADDR ? 9'h7b : _GEN_607; // @[RAM_ST.scala 32:46]
  assign _GEN_609 = 9'h7c == RADDR ? 9'h7c : _GEN_608; // @[RAM_ST.scala 32:46]
  assign _GEN_610 = 9'h7d == RADDR ? 9'h7d : _GEN_609; // @[RAM_ST.scala 32:46]
  assign _GEN_611 = 9'h7e == RADDR ? 9'h7e : _GEN_610; // @[RAM_ST.scala 32:46]
  assign _GEN_612 = 9'h7f == RADDR ? 9'h7f : _GEN_611; // @[RAM_ST.scala 32:46]
  assign _GEN_613 = 9'h80 == RADDR ? 9'h80 : _GEN_612; // @[RAM_ST.scala 32:46]
  assign _GEN_614 = 9'h81 == RADDR ? 9'h81 : _GEN_613; // @[RAM_ST.scala 32:46]
  assign _GEN_615 = 9'h82 == RADDR ? 9'h82 : _GEN_614; // @[RAM_ST.scala 32:46]
  assign _GEN_616 = 9'h83 == RADDR ? 9'h83 : _GEN_615; // @[RAM_ST.scala 32:46]
  assign _GEN_617 = 9'h84 == RADDR ? 9'h84 : _GEN_616; // @[RAM_ST.scala 32:46]
  assign _GEN_618 = 9'h85 == RADDR ? 9'h85 : _GEN_617; // @[RAM_ST.scala 32:46]
  assign _GEN_619 = 9'h86 == RADDR ? 9'h86 : _GEN_618; // @[RAM_ST.scala 32:46]
  assign _GEN_620 = 9'h87 == RADDR ? 9'h87 : _GEN_619; // @[RAM_ST.scala 32:46]
  assign _GEN_621 = 9'h88 == RADDR ? 9'h88 : _GEN_620; // @[RAM_ST.scala 32:46]
  assign _GEN_622 = 9'h89 == RADDR ? 9'h89 : _GEN_621; // @[RAM_ST.scala 32:46]
  assign _GEN_623 = 9'h8a == RADDR ? 9'h8a : _GEN_622; // @[RAM_ST.scala 32:46]
  assign _GEN_624 = 9'h8b == RADDR ? 9'h8b : _GEN_623; // @[RAM_ST.scala 32:46]
  assign _GEN_625 = 9'h8c == RADDR ? 9'h8c : _GEN_624; // @[RAM_ST.scala 32:46]
  assign _GEN_626 = 9'h8d == RADDR ? 9'h8d : _GEN_625; // @[RAM_ST.scala 32:46]
  assign _GEN_627 = 9'h8e == RADDR ? 9'h8e : _GEN_626; // @[RAM_ST.scala 32:46]
  assign _GEN_628 = 9'h8f == RADDR ? 9'h8f : _GEN_627; // @[RAM_ST.scala 32:46]
  assign _GEN_629 = 9'h90 == RADDR ? 9'h90 : _GEN_628; // @[RAM_ST.scala 32:46]
  assign _GEN_630 = 9'h91 == RADDR ? 9'h91 : _GEN_629; // @[RAM_ST.scala 32:46]
  assign _GEN_631 = 9'h92 == RADDR ? 9'h92 : _GEN_630; // @[RAM_ST.scala 32:46]
  assign _GEN_632 = 9'h93 == RADDR ? 9'h93 : _GEN_631; // @[RAM_ST.scala 32:46]
  assign _GEN_633 = 9'h94 == RADDR ? 9'h94 : _GEN_632; // @[RAM_ST.scala 32:46]
  assign _GEN_634 = 9'h95 == RADDR ? 9'h95 : _GEN_633; // @[RAM_ST.scala 32:46]
  assign _GEN_635 = 9'h96 == RADDR ? 9'h96 : _GEN_634; // @[RAM_ST.scala 32:46]
  assign _GEN_636 = 9'h97 == RADDR ? 9'h97 : _GEN_635; // @[RAM_ST.scala 32:46]
  assign _GEN_637 = 9'h98 == RADDR ? 9'h98 : _GEN_636; // @[RAM_ST.scala 32:46]
  assign _GEN_638 = 9'h99 == RADDR ? 9'h99 : _GEN_637; // @[RAM_ST.scala 32:46]
  assign _GEN_639 = 9'h9a == RADDR ? 9'h9a : _GEN_638; // @[RAM_ST.scala 32:46]
  assign _GEN_640 = 9'h9b == RADDR ? 9'h9b : _GEN_639; // @[RAM_ST.scala 32:46]
  assign _GEN_641 = 9'h9c == RADDR ? 9'h9c : _GEN_640; // @[RAM_ST.scala 32:46]
  assign _GEN_642 = 9'h9d == RADDR ? 9'h9d : _GEN_641; // @[RAM_ST.scala 32:46]
  assign _GEN_643 = 9'h9e == RADDR ? 9'h9e : _GEN_642; // @[RAM_ST.scala 32:46]
  assign _GEN_644 = 9'h9f == RADDR ? 9'h9f : _GEN_643; // @[RAM_ST.scala 32:46]
  assign _GEN_645 = 9'ha0 == RADDR ? 9'ha0 : _GEN_644; // @[RAM_ST.scala 32:46]
  assign _GEN_646 = 9'ha1 == RADDR ? 9'ha1 : _GEN_645; // @[RAM_ST.scala 32:46]
  assign _GEN_647 = 9'ha2 == RADDR ? 9'ha2 : _GEN_646; // @[RAM_ST.scala 32:46]
  assign _GEN_648 = 9'ha3 == RADDR ? 9'ha3 : _GEN_647; // @[RAM_ST.scala 32:46]
  assign _GEN_649 = 9'ha4 == RADDR ? 9'ha4 : _GEN_648; // @[RAM_ST.scala 32:46]
  assign _GEN_650 = 9'ha5 == RADDR ? 9'ha5 : _GEN_649; // @[RAM_ST.scala 32:46]
  assign _GEN_651 = 9'ha6 == RADDR ? 9'ha6 : _GEN_650; // @[RAM_ST.scala 32:46]
  assign _GEN_652 = 9'ha7 == RADDR ? 9'ha7 : _GEN_651; // @[RAM_ST.scala 32:46]
  assign _GEN_653 = 9'ha8 == RADDR ? 9'ha8 : _GEN_652; // @[RAM_ST.scala 32:46]
  assign _GEN_654 = 9'ha9 == RADDR ? 9'ha9 : _GEN_653; // @[RAM_ST.scala 32:46]
  assign _GEN_655 = 9'haa == RADDR ? 9'haa : _GEN_654; // @[RAM_ST.scala 32:46]
  assign _GEN_656 = 9'hab == RADDR ? 9'hab : _GEN_655; // @[RAM_ST.scala 32:46]
  assign _GEN_657 = 9'hac == RADDR ? 9'hac : _GEN_656; // @[RAM_ST.scala 32:46]
  assign _GEN_658 = 9'had == RADDR ? 9'had : _GEN_657; // @[RAM_ST.scala 32:46]
  assign _GEN_659 = 9'hae == RADDR ? 9'hae : _GEN_658; // @[RAM_ST.scala 32:46]
  assign _GEN_660 = 9'haf == RADDR ? 9'haf : _GEN_659; // @[RAM_ST.scala 32:46]
  assign _GEN_661 = 9'hb0 == RADDR ? 9'hb0 : _GEN_660; // @[RAM_ST.scala 32:46]
  assign _GEN_662 = 9'hb1 == RADDR ? 9'hb1 : _GEN_661; // @[RAM_ST.scala 32:46]
  assign _GEN_663 = 9'hb2 == RADDR ? 9'hb2 : _GEN_662; // @[RAM_ST.scala 32:46]
  assign _GEN_664 = 9'hb3 == RADDR ? 9'hb3 : _GEN_663; // @[RAM_ST.scala 32:46]
  assign _GEN_665 = 9'hb4 == RADDR ? 9'hb4 : _GEN_664; // @[RAM_ST.scala 32:46]
  assign _GEN_666 = 9'hb5 == RADDR ? 9'hb5 : _GEN_665; // @[RAM_ST.scala 32:46]
  assign _GEN_667 = 9'hb6 == RADDR ? 9'hb6 : _GEN_666; // @[RAM_ST.scala 32:46]
  assign _GEN_668 = 9'hb7 == RADDR ? 9'hb7 : _GEN_667; // @[RAM_ST.scala 32:46]
  assign _GEN_669 = 9'hb8 == RADDR ? 9'hb8 : _GEN_668; // @[RAM_ST.scala 32:46]
  assign _GEN_670 = 9'hb9 == RADDR ? 9'hb9 : _GEN_669; // @[RAM_ST.scala 32:46]
  assign _GEN_671 = 9'hba == RADDR ? 9'hba : _GEN_670; // @[RAM_ST.scala 32:46]
  assign _GEN_672 = 9'hbb == RADDR ? 9'hbb : _GEN_671; // @[RAM_ST.scala 32:46]
  assign _GEN_673 = 9'hbc == RADDR ? 9'hbc : _GEN_672; // @[RAM_ST.scala 32:46]
  assign _GEN_674 = 9'hbd == RADDR ? 9'hbd : _GEN_673; // @[RAM_ST.scala 32:46]
  assign _GEN_675 = 9'hbe == RADDR ? 9'hbe : _GEN_674; // @[RAM_ST.scala 32:46]
  assign _GEN_676 = 9'hbf == RADDR ? 9'hbf : _GEN_675; // @[RAM_ST.scala 32:46]
  assign _GEN_677 = 9'hc0 == RADDR ? 9'hc0 : _GEN_676; // @[RAM_ST.scala 32:46]
  assign _GEN_678 = 9'hc1 == RADDR ? 9'hc1 : _GEN_677; // @[RAM_ST.scala 32:46]
  assign _GEN_679 = 9'hc2 == RADDR ? 9'hc2 : _GEN_678; // @[RAM_ST.scala 32:46]
  assign _GEN_680 = 9'hc3 == RADDR ? 9'hc3 : _GEN_679; // @[RAM_ST.scala 32:46]
  assign _GEN_681 = 9'hc4 == RADDR ? 9'hc4 : _GEN_680; // @[RAM_ST.scala 32:46]
  assign _GEN_682 = 9'hc5 == RADDR ? 9'hc5 : _GEN_681; // @[RAM_ST.scala 32:46]
  assign _GEN_683 = 9'hc6 == RADDR ? 9'hc6 : _GEN_682; // @[RAM_ST.scala 32:46]
  assign _GEN_684 = 9'hc7 == RADDR ? 9'hc7 : _GEN_683; // @[RAM_ST.scala 32:46]
  assign _GEN_685 = 9'hc8 == RADDR ? 9'hc8 : _GEN_684; // @[RAM_ST.scala 32:46]
  assign _GEN_686 = 9'hc9 == RADDR ? 9'hc9 : _GEN_685; // @[RAM_ST.scala 32:46]
  assign _GEN_687 = 9'hca == RADDR ? 9'hca : _GEN_686; // @[RAM_ST.scala 32:46]
  assign _GEN_688 = 9'hcb == RADDR ? 9'hcb : _GEN_687; // @[RAM_ST.scala 32:46]
  assign _GEN_689 = 9'hcc == RADDR ? 9'hcc : _GEN_688; // @[RAM_ST.scala 32:46]
  assign _GEN_690 = 9'hcd == RADDR ? 9'hcd : _GEN_689; // @[RAM_ST.scala 32:46]
  assign _GEN_691 = 9'hce == RADDR ? 9'hce : _GEN_690; // @[RAM_ST.scala 32:46]
  assign _GEN_692 = 9'hcf == RADDR ? 9'hcf : _GEN_691; // @[RAM_ST.scala 32:46]
  assign _GEN_693 = 9'hd0 == RADDR ? 9'hd0 : _GEN_692; // @[RAM_ST.scala 32:46]
  assign _GEN_694 = 9'hd1 == RADDR ? 9'hd1 : _GEN_693; // @[RAM_ST.scala 32:46]
  assign _GEN_695 = 9'hd2 == RADDR ? 9'hd2 : _GEN_694; // @[RAM_ST.scala 32:46]
  assign _GEN_696 = 9'hd3 == RADDR ? 9'hd3 : _GEN_695; // @[RAM_ST.scala 32:46]
  assign _GEN_697 = 9'hd4 == RADDR ? 9'hd4 : _GEN_696; // @[RAM_ST.scala 32:46]
  assign _GEN_698 = 9'hd5 == RADDR ? 9'hd5 : _GEN_697; // @[RAM_ST.scala 32:46]
  assign _GEN_699 = 9'hd6 == RADDR ? 9'hd6 : _GEN_698; // @[RAM_ST.scala 32:46]
  assign _GEN_700 = 9'hd7 == RADDR ? 9'hd7 : _GEN_699; // @[RAM_ST.scala 32:46]
  assign _GEN_701 = 9'hd8 == RADDR ? 9'hd8 : _GEN_700; // @[RAM_ST.scala 32:46]
  assign _GEN_702 = 9'hd9 == RADDR ? 9'hd9 : _GEN_701; // @[RAM_ST.scala 32:46]
  assign _GEN_703 = 9'hda == RADDR ? 9'hda : _GEN_702; // @[RAM_ST.scala 32:46]
  assign _GEN_704 = 9'hdb == RADDR ? 9'hdb : _GEN_703; // @[RAM_ST.scala 32:46]
  assign _GEN_705 = 9'hdc == RADDR ? 9'hdc : _GEN_704; // @[RAM_ST.scala 32:46]
  assign _GEN_706 = 9'hdd == RADDR ? 9'hdd : _GEN_705; // @[RAM_ST.scala 32:46]
  assign _GEN_707 = 9'hde == RADDR ? 9'hde : _GEN_706; // @[RAM_ST.scala 32:46]
  assign _GEN_708 = 9'hdf == RADDR ? 9'hdf : _GEN_707; // @[RAM_ST.scala 32:46]
  assign _GEN_709 = 9'he0 == RADDR ? 9'he0 : _GEN_708; // @[RAM_ST.scala 32:46]
  assign _GEN_710 = 9'he1 == RADDR ? 9'he1 : _GEN_709; // @[RAM_ST.scala 32:46]
  assign _GEN_711 = 9'he2 == RADDR ? 9'he2 : _GEN_710; // @[RAM_ST.scala 32:46]
  assign _GEN_712 = 9'he3 == RADDR ? 9'he3 : _GEN_711; // @[RAM_ST.scala 32:46]
  assign _GEN_713 = 9'he4 == RADDR ? 9'he4 : _GEN_712; // @[RAM_ST.scala 32:46]
  assign _GEN_714 = 9'he5 == RADDR ? 9'he5 : _GEN_713; // @[RAM_ST.scala 32:46]
  assign _GEN_715 = 9'he6 == RADDR ? 9'he6 : _GEN_714; // @[RAM_ST.scala 32:46]
  assign _GEN_716 = 9'he7 == RADDR ? 9'he7 : _GEN_715; // @[RAM_ST.scala 32:46]
  assign _GEN_717 = 9'he8 == RADDR ? 9'he8 : _GEN_716; // @[RAM_ST.scala 32:46]
  assign _GEN_718 = 9'he9 == RADDR ? 9'he9 : _GEN_717; // @[RAM_ST.scala 32:46]
  assign _GEN_719 = 9'hea == RADDR ? 9'hea : _GEN_718; // @[RAM_ST.scala 32:46]
  assign _GEN_720 = 9'heb == RADDR ? 9'heb : _GEN_719; // @[RAM_ST.scala 32:46]
  assign _GEN_721 = 9'hec == RADDR ? 9'hec : _GEN_720; // @[RAM_ST.scala 32:46]
  assign _GEN_722 = 9'hed == RADDR ? 9'hed : _GEN_721; // @[RAM_ST.scala 32:46]
  assign _GEN_723 = 9'hee == RADDR ? 9'hee : _GEN_722; // @[RAM_ST.scala 32:46]
  assign _GEN_724 = 9'hef == RADDR ? 9'hef : _GEN_723; // @[RAM_ST.scala 32:46]
  assign _GEN_725 = 9'hf0 == RADDR ? 9'hf0 : _GEN_724; // @[RAM_ST.scala 32:46]
  assign _GEN_726 = 9'hf1 == RADDR ? 9'hf1 : _GEN_725; // @[RAM_ST.scala 32:46]
  assign _GEN_727 = 9'hf2 == RADDR ? 9'hf2 : _GEN_726; // @[RAM_ST.scala 32:46]
  assign _GEN_728 = 9'hf3 == RADDR ? 9'hf3 : _GEN_727; // @[RAM_ST.scala 32:46]
  assign _GEN_729 = 9'hf4 == RADDR ? 9'hf4 : _GEN_728; // @[RAM_ST.scala 32:46]
  assign _GEN_730 = 9'hf5 == RADDR ? 9'hf5 : _GEN_729; // @[RAM_ST.scala 32:46]
  assign _GEN_731 = 9'hf6 == RADDR ? 9'hf6 : _GEN_730; // @[RAM_ST.scala 32:46]
  assign _GEN_732 = 9'hf7 == RADDR ? 9'hf7 : _GEN_731; // @[RAM_ST.scala 32:46]
  assign _GEN_733 = 9'hf8 == RADDR ? 9'hf8 : _GEN_732; // @[RAM_ST.scala 32:46]
  assign _GEN_734 = 9'hf9 == RADDR ? 9'hf9 : _GEN_733; // @[RAM_ST.scala 32:46]
  assign _GEN_735 = 9'hfa == RADDR ? 9'hfa : _GEN_734; // @[RAM_ST.scala 32:46]
  assign _GEN_736 = 9'hfb == RADDR ? 9'hfb : _GEN_735; // @[RAM_ST.scala 32:46]
  assign _GEN_737 = 9'hfc == RADDR ? 9'hfc : _GEN_736; // @[RAM_ST.scala 32:46]
  assign _GEN_738 = 9'hfd == RADDR ? 9'hfd : _GEN_737; // @[RAM_ST.scala 32:46]
  assign _GEN_739 = 9'hfe == RADDR ? 9'hfe : _GEN_738; // @[RAM_ST.scala 32:46]
  assign _GEN_740 = 9'hff == RADDR ? 9'hff : _GEN_739; // @[RAM_ST.scala 32:46]
  assign _GEN_741 = 9'h100 == RADDR ? 9'h100 : _GEN_740; // @[RAM_ST.scala 32:46]
  assign _GEN_742 = 9'h101 == RADDR ? 9'h101 : _GEN_741; // @[RAM_ST.scala 32:46]
  assign _GEN_743 = 9'h102 == RADDR ? 9'h102 : _GEN_742; // @[RAM_ST.scala 32:46]
  assign _GEN_744 = 9'h103 == RADDR ? 9'h103 : _GEN_743; // @[RAM_ST.scala 32:46]
  assign _GEN_745 = 9'h104 == RADDR ? 9'h104 : _GEN_744; // @[RAM_ST.scala 32:46]
  assign _GEN_746 = 9'h105 == RADDR ? 9'h105 : _GEN_745; // @[RAM_ST.scala 32:46]
  assign _GEN_747 = 9'h106 == RADDR ? 9'h106 : _GEN_746; // @[RAM_ST.scala 32:46]
  assign _GEN_748 = 9'h107 == RADDR ? 9'h107 : _GEN_747; // @[RAM_ST.scala 32:46]
  assign _GEN_749 = 9'h108 == RADDR ? 9'h108 : _GEN_748; // @[RAM_ST.scala 32:46]
  assign _GEN_750 = 9'h109 == RADDR ? 9'h109 : _GEN_749; // @[RAM_ST.scala 32:46]
  assign _GEN_751 = 9'h10a == RADDR ? 9'h10a : _GEN_750; // @[RAM_ST.scala 32:46]
  assign _GEN_752 = 9'h10b == RADDR ? 9'h10b : _GEN_751; // @[RAM_ST.scala 32:46]
  assign _GEN_753 = 9'h10c == RADDR ? 9'h10c : _GEN_752; // @[RAM_ST.scala 32:46]
  assign _GEN_754 = 9'h10d == RADDR ? 9'h10d : _GEN_753; // @[RAM_ST.scala 32:46]
  assign _GEN_755 = 9'h10e == RADDR ? 9'h10e : _GEN_754; // @[RAM_ST.scala 32:46]
  assign _GEN_756 = 9'h10f == RADDR ? 9'h10f : _GEN_755; // @[RAM_ST.scala 32:46]
  assign _GEN_757 = 9'h110 == RADDR ? 9'h110 : _GEN_756; // @[RAM_ST.scala 32:46]
  assign _GEN_758 = 9'h111 == RADDR ? 9'h111 : _GEN_757; // @[RAM_ST.scala 32:46]
  assign _GEN_759 = 9'h112 == RADDR ? 9'h112 : _GEN_758; // @[RAM_ST.scala 32:46]
  assign _GEN_760 = 9'h113 == RADDR ? 9'h113 : _GEN_759; // @[RAM_ST.scala 32:46]
  assign _GEN_761 = 9'h114 == RADDR ? 9'h114 : _GEN_760; // @[RAM_ST.scala 32:46]
  assign _GEN_762 = 9'h115 == RADDR ? 9'h115 : _GEN_761; // @[RAM_ST.scala 32:46]
  assign _GEN_763 = 9'h116 == RADDR ? 9'h116 : _GEN_762; // @[RAM_ST.scala 32:46]
  assign _GEN_764 = 9'h117 == RADDR ? 9'h117 : _GEN_763; // @[RAM_ST.scala 32:46]
  assign _GEN_765 = 9'h118 == RADDR ? 9'h118 : _GEN_764; // @[RAM_ST.scala 32:46]
  assign _GEN_766 = 9'h119 == RADDR ? 9'h119 : _GEN_765; // @[RAM_ST.scala 32:46]
  assign _GEN_767 = 9'h11a == RADDR ? 9'h11a : _GEN_766; // @[RAM_ST.scala 32:46]
  assign _GEN_768 = 9'h11b == RADDR ? 9'h11b : _GEN_767; // @[RAM_ST.scala 32:46]
  assign _GEN_769 = 9'h11c == RADDR ? 9'h11c : _GEN_768; // @[RAM_ST.scala 32:46]
  assign _GEN_770 = 9'h11d == RADDR ? 9'h11d : _GEN_769; // @[RAM_ST.scala 32:46]
  assign _GEN_771 = 9'h11e == RADDR ? 9'h11e : _GEN_770; // @[RAM_ST.scala 32:46]
  assign _GEN_772 = 9'h11f == RADDR ? 9'h11f : _GEN_771; // @[RAM_ST.scala 32:46]
  assign _GEN_773 = 9'h120 == RADDR ? 9'h120 : _GEN_772; // @[RAM_ST.scala 32:46]
  assign _GEN_774 = 9'h121 == RADDR ? 9'h121 : _GEN_773; // @[RAM_ST.scala 32:46]
  assign _GEN_775 = 9'h122 == RADDR ? 9'h122 : _GEN_774; // @[RAM_ST.scala 32:46]
  assign _GEN_776 = 9'h123 == RADDR ? 9'h123 : _GEN_775; // @[RAM_ST.scala 32:46]
  assign _GEN_777 = 9'h124 == RADDR ? 9'h124 : _GEN_776; // @[RAM_ST.scala 32:46]
  assign _GEN_778 = 9'h125 == RADDR ? 9'h125 : _GEN_777; // @[RAM_ST.scala 32:46]
  assign _GEN_779 = 9'h126 == RADDR ? 9'h126 : _GEN_778; // @[RAM_ST.scala 32:46]
  assign _GEN_780 = 9'h127 == RADDR ? 9'h127 : _GEN_779; // @[RAM_ST.scala 32:46]
  assign _GEN_781 = 9'h128 == RADDR ? 9'h128 : _GEN_780; // @[RAM_ST.scala 32:46]
  assign _GEN_782 = 9'h129 == RADDR ? 9'h129 : _GEN_781; // @[RAM_ST.scala 32:46]
  assign _GEN_783 = 9'h12a == RADDR ? 9'h12a : _GEN_782; // @[RAM_ST.scala 32:46]
  assign _GEN_784 = 9'h12b == RADDR ? 9'h12b : _GEN_783; // @[RAM_ST.scala 32:46]
  assign _GEN_785 = 9'h12c == RADDR ? 9'h12c : _GEN_784; // @[RAM_ST.scala 32:46]
  assign _GEN_786 = 9'h12d == RADDR ? 9'h12d : _GEN_785; // @[RAM_ST.scala 32:46]
  assign _GEN_787 = 9'h12e == RADDR ? 9'h12e : _GEN_786; // @[RAM_ST.scala 32:46]
  assign _GEN_788 = 9'h12f == RADDR ? 9'h12f : _GEN_787; // @[RAM_ST.scala 32:46]
  assign _GEN_789 = 9'h130 == RADDR ? 9'h130 : _GEN_788; // @[RAM_ST.scala 32:46]
  assign _GEN_790 = 9'h131 == RADDR ? 9'h131 : _GEN_789; // @[RAM_ST.scala 32:46]
  assign _GEN_791 = 9'h132 == RADDR ? 9'h132 : _GEN_790; // @[RAM_ST.scala 32:46]
  assign _GEN_792 = 9'h133 == RADDR ? 9'h133 : _GEN_791; // @[RAM_ST.scala 32:46]
  assign _GEN_793 = 9'h134 == RADDR ? 9'h134 : _GEN_792; // @[RAM_ST.scala 32:46]
  assign _GEN_794 = 9'h135 == RADDR ? 9'h135 : _GEN_793; // @[RAM_ST.scala 32:46]
  assign _GEN_795 = 9'h136 == RADDR ? 9'h136 : _GEN_794; // @[RAM_ST.scala 32:46]
  assign _GEN_796 = 9'h137 == RADDR ? 9'h137 : _GEN_795; // @[RAM_ST.scala 32:46]
  assign _GEN_797 = 9'h138 == RADDR ? 9'h138 : _GEN_796; // @[RAM_ST.scala 32:46]
  assign _GEN_798 = 9'h139 == RADDR ? 9'h139 : _GEN_797; // @[RAM_ST.scala 32:46]
  assign _GEN_799 = 9'h13a == RADDR ? 9'h13a : _GEN_798; // @[RAM_ST.scala 32:46]
  assign _GEN_800 = 9'h13b == RADDR ? 9'h13b : _GEN_799; // @[RAM_ST.scala 32:46]
  assign _GEN_801 = 9'h13c == RADDR ? 9'h13c : _GEN_800; // @[RAM_ST.scala 32:46]
  assign _GEN_802 = 9'h13d == RADDR ? 9'h13d : _GEN_801; // @[RAM_ST.scala 32:46]
  assign _GEN_803 = 9'h13e == RADDR ? 9'h13e : _GEN_802; // @[RAM_ST.scala 32:46]
  assign _GEN_804 = 9'h13f == RADDR ? 9'h13f : _GEN_803; // @[RAM_ST.scala 32:46]
  assign _GEN_805 = 9'h140 == RADDR ? 9'h140 : _GEN_804; // @[RAM_ST.scala 32:46]
  assign _GEN_806 = 9'h141 == RADDR ? 9'h141 : _GEN_805; // @[RAM_ST.scala 32:46]
  assign _GEN_807 = 9'h142 == RADDR ? 9'h142 : _GEN_806; // @[RAM_ST.scala 32:46]
  assign _GEN_808 = 9'h143 == RADDR ? 9'h143 : _GEN_807; // @[RAM_ST.scala 32:46]
  assign _GEN_809 = 9'h144 == RADDR ? 9'h144 : _GEN_808; // @[RAM_ST.scala 32:46]
  assign _GEN_810 = 9'h145 == RADDR ? 9'h145 : _GEN_809; // @[RAM_ST.scala 32:46]
  assign _GEN_811 = 9'h146 == RADDR ? 9'h146 : _GEN_810; // @[RAM_ST.scala 32:46]
  assign _GEN_812 = 9'h147 == RADDR ? 9'h147 : _GEN_811; // @[RAM_ST.scala 32:46]
  assign _GEN_813 = 9'h148 == RADDR ? 9'h148 : _GEN_812; // @[RAM_ST.scala 32:46]
  assign _GEN_814 = 9'h149 == RADDR ? 9'h149 : _GEN_813; // @[RAM_ST.scala 32:46]
  assign _GEN_815 = 9'h14a == RADDR ? 9'h14a : _GEN_814; // @[RAM_ST.scala 32:46]
  assign _GEN_816 = 9'h14b == RADDR ? 9'h14b : _GEN_815; // @[RAM_ST.scala 32:46]
  assign _GEN_817 = 9'h14c == RADDR ? 9'h14c : _GEN_816; // @[RAM_ST.scala 32:46]
  assign _GEN_818 = 9'h14d == RADDR ? 9'h14d : _GEN_817; // @[RAM_ST.scala 32:46]
  assign _GEN_819 = 9'h14e == RADDR ? 9'h14e : _GEN_818; // @[RAM_ST.scala 32:46]
  assign _GEN_820 = 9'h14f == RADDR ? 9'h14f : _GEN_819; // @[RAM_ST.scala 32:46]
  assign _GEN_821 = 9'h150 == RADDR ? 9'h150 : _GEN_820; // @[RAM_ST.scala 32:46]
  assign _GEN_822 = 9'h151 == RADDR ? 9'h151 : _GEN_821; // @[RAM_ST.scala 32:46]
  assign _GEN_823 = 9'h152 == RADDR ? 9'h152 : _GEN_822; // @[RAM_ST.scala 32:46]
  assign _GEN_824 = 9'h153 == RADDR ? 9'h153 : _GEN_823; // @[RAM_ST.scala 32:46]
  assign _GEN_825 = 9'h154 == RADDR ? 9'h154 : _GEN_824; // @[RAM_ST.scala 32:46]
  assign _GEN_826 = 9'h155 == RADDR ? 9'h155 : _GEN_825; // @[RAM_ST.scala 32:46]
  assign _GEN_827 = 9'h156 == RADDR ? 9'h156 : _GEN_826; // @[RAM_ST.scala 32:46]
  assign _GEN_828 = 9'h157 == RADDR ? 9'h157 : _GEN_827; // @[RAM_ST.scala 32:46]
  assign _GEN_829 = 9'h158 == RADDR ? 9'h158 : _GEN_828; // @[RAM_ST.scala 32:46]
  assign _GEN_830 = 9'h159 == RADDR ? 9'h159 : _GEN_829; // @[RAM_ST.scala 32:46]
  assign _GEN_831 = 9'h15a == RADDR ? 9'h15a : _GEN_830; // @[RAM_ST.scala 32:46]
  assign _GEN_832 = 9'h15b == RADDR ? 9'h15b : _GEN_831; // @[RAM_ST.scala 32:46]
  assign _GEN_833 = 9'h15c == RADDR ? 9'h15c : _GEN_832; // @[RAM_ST.scala 32:46]
  assign _GEN_834 = 9'h15d == RADDR ? 9'h15d : _GEN_833; // @[RAM_ST.scala 32:46]
  assign _GEN_835 = 9'h15e == RADDR ? 9'h15e : _GEN_834; // @[RAM_ST.scala 32:46]
  assign _GEN_836 = 9'h15f == RADDR ? 9'h15f : _GEN_835; // @[RAM_ST.scala 32:46]
  assign _GEN_837 = 9'h160 == RADDR ? 9'h160 : _GEN_836; // @[RAM_ST.scala 32:46]
  assign _GEN_838 = 9'h161 == RADDR ? 9'h161 : _GEN_837; // @[RAM_ST.scala 32:46]
  assign _GEN_839 = 9'h162 == RADDR ? 9'h162 : _GEN_838; // @[RAM_ST.scala 32:46]
  assign _GEN_840 = 9'h163 == RADDR ? 9'h163 : _GEN_839; // @[RAM_ST.scala 32:46]
  assign _GEN_841 = 9'h164 == RADDR ? 9'h164 : _GEN_840; // @[RAM_ST.scala 32:46]
  assign _GEN_842 = 9'h165 == RADDR ? 9'h165 : _GEN_841; // @[RAM_ST.scala 32:46]
  assign _GEN_843 = 9'h166 == RADDR ? 9'h166 : _GEN_842; // @[RAM_ST.scala 32:46]
  assign _GEN_844 = 9'h167 == RADDR ? 9'h167 : _GEN_843; // @[RAM_ST.scala 32:46]
  assign _GEN_845 = 9'h168 == RADDR ? 9'h168 : _GEN_844; // @[RAM_ST.scala 32:46]
  assign _GEN_846 = 9'h169 == RADDR ? 9'h169 : _GEN_845; // @[RAM_ST.scala 32:46]
  assign _GEN_847 = 9'h16a == RADDR ? 9'h16a : _GEN_846; // @[RAM_ST.scala 32:46]
  assign _GEN_848 = 9'h16b == RADDR ? 9'h16b : _GEN_847; // @[RAM_ST.scala 32:46]
  assign _GEN_849 = 9'h16c == RADDR ? 9'h16c : _GEN_848; // @[RAM_ST.scala 32:46]
  assign _GEN_850 = 9'h16d == RADDR ? 9'h16d : _GEN_849; // @[RAM_ST.scala 32:46]
  assign _GEN_851 = 9'h16e == RADDR ? 9'h16e : _GEN_850; // @[RAM_ST.scala 32:46]
  assign _GEN_852 = 9'h16f == RADDR ? 9'h16f : _GEN_851; // @[RAM_ST.scala 32:46]
  assign _GEN_853 = 9'h170 == RADDR ? 9'h170 : _GEN_852; // @[RAM_ST.scala 32:46]
  assign _GEN_854 = 9'h171 == RADDR ? 9'h171 : _GEN_853; // @[RAM_ST.scala 32:46]
  assign _GEN_855 = 9'h172 == RADDR ? 9'h172 : _GEN_854; // @[RAM_ST.scala 32:46]
  assign _GEN_856 = 9'h173 == RADDR ? 9'h173 : _GEN_855; // @[RAM_ST.scala 32:46]
  assign _GEN_857 = 9'h174 == RADDR ? 9'h174 : _GEN_856; // @[RAM_ST.scala 32:46]
  assign _GEN_858 = 9'h175 == RADDR ? 9'h175 : _GEN_857; // @[RAM_ST.scala 32:46]
  assign _GEN_859 = 9'h176 == RADDR ? 9'h176 : _GEN_858; // @[RAM_ST.scala 32:46]
  assign _GEN_860 = 9'h177 == RADDR ? 9'h177 : _GEN_859; // @[RAM_ST.scala 32:46]
  assign _GEN_861 = 9'h178 == RADDR ? 9'h178 : _GEN_860; // @[RAM_ST.scala 32:46]
  assign _GEN_862 = 9'h179 == RADDR ? 9'h179 : _GEN_861; // @[RAM_ST.scala 32:46]
  assign _GEN_863 = 9'h17a == RADDR ? 9'h17a : _GEN_862; // @[RAM_ST.scala 32:46]
  assign _GEN_864 = 9'h17b == RADDR ? 9'h17b : _GEN_863; // @[RAM_ST.scala 32:46]
  assign _GEN_865 = 9'h17c == RADDR ? 9'h17c : _GEN_864; // @[RAM_ST.scala 32:46]
  assign _GEN_866 = 9'h17d == RADDR ? 9'h17d : _GEN_865; // @[RAM_ST.scala 32:46]
  assign _GEN_867 = 9'h17e == RADDR ? 9'h17e : _GEN_866; // @[RAM_ST.scala 32:46]
  assign _GEN_868 = 9'h17f == RADDR ? 9'h17f : _GEN_867; // @[RAM_ST.scala 32:46]
  assign _GEN_869 = 9'h180 == RADDR ? 9'h180 : _GEN_868; // @[RAM_ST.scala 32:46]
  assign _GEN_870 = 9'h181 == RADDR ? 9'h181 : _GEN_869; // @[RAM_ST.scala 32:46]
  assign _GEN_871 = 9'h182 == RADDR ? 9'h182 : _GEN_870; // @[RAM_ST.scala 32:46]
  assign _GEN_872 = 9'h183 == RADDR ? 9'h183 : _GEN_871; // @[RAM_ST.scala 32:46]
  assign _GEN_873 = 9'h184 == RADDR ? 9'h184 : _GEN_872; // @[RAM_ST.scala 32:46]
  assign _GEN_874 = 9'h185 == RADDR ? 9'h185 : _GEN_873; // @[RAM_ST.scala 32:46]
  assign _GEN_875 = 9'h186 == RADDR ? 9'h186 : _GEN_874; // @[RAM_ST.scala 32:46]
  assign _GEN_876 = 9'h187 == RADDR ? 9'h187 : _GEN_875; // @[RAM_ST.scala 32:46]
  assign _GEN_877 = 9'h188 == RADDR ? 9'h188 : _GEN_876; // @[RAM_ST.scala 32:46]
  assign _GEN_878 = 9'h189 == RADDR ? 9'h189 : _GEN_877; // @[RAM_ST.scala 32:46]
  assign _GEN_879 = 9'h18a == RADDR ? 9'h18a : _GEN_878; // @[RAM_ST.scala 32:46]
  assign _GEN_880 = 9'h18b == RADDR ? 9'h18b : _GEN_879; // @[RAM_ST.scala 32:46]
  assign _GEN_881 = 9'h18c == RADDR ? 9'h18c : _GEN_880; // @[RAM_ST.scala 32:46]
  assign _GEN_882 = 9'h18d == RADDR ? 9'h18d : _GEN_881; // @[RAM_ST.scala 32:46]
  assign _GEN_883 = 9'h18e == RADDR ? 9'h18e : _GEN_882; // @[RAM_ST.scala 32:46]
  assign _GEN_884 = 9'h18f == RADDR ? 9'h18f : _GEN_883; // @[RAM_ST.scala 32:46]
  assign _GEN_885 = 9'h190 == RADDR ? 9'h190 : _GEN_884; // @[RAM_ST.scala 32:46]
  assign _GEN_886 = 9'h191 == RADDR ? 9'h191 : _GEN_885; // @[RAM_ST.scala 32:46]
  assign _GEN_887 = 9'h192 == RADDR ? 9'h192 : _GEN_886; // @[RAM_ST.scala 32:46]
  assign _GEN_888 = 9'h193 == RADDR ? 9'h193 : _GEN_887; // @[RAM_ST.scala 32:46]
  assign _GEN_889 = 9'h194 == RADDR ? 9'h194 : _GEN_888; // @[RAM_ST.scala 32:46]
  assign _GEN_890 = 9'h195 == RADDR ? 9'h195 : _GEN_889; // @[RAM_ST.scala 32:46]
  assign _GEN_891 = 9'h196 == RADDR ? 9'h196 : _GEN_890; // @[RAM_ST.scala 32:46]
  assign _GEN_892 = 9'h197 == RADDR ? 9'h197 : _GEN_891; // @[RAM_ST.scala 32:46]
  assign _GEN_893 = 9'h198 == RADDR ? 9'h198 : _GEN_892; // @[RAM_ST.scala 32:46]
  assign _GEN_894 = 9'h199 == RADDR ? 9'h199 : _GEN_893; // @[RAM_ST.scala 32:46]
  assign _GEN_895 = 9'h19a == RADDR ? 9'h19a : _GEN_894; // @[RAM_ST.scala 32:46]
  assign _GEN_896 = 9'h19b == RADDR ? 9'h19b : _GEN_895; // @[RAM_ST.scala 32:46]
  assign _GEN_897 = 9'h19c == RADDR ? 9'h19c : _GEN_896; // @[RAM_ST.scala 32:46]
  assign _GEN_898 = 9'h19d == RADDR ? 9'h19d : _GEN_897; // @[RAM_ST.scala 32:46]
  assign _GEN_899 = 9'h19e == RADDR ? 9'h19e : _GEN_898; // @[RAM_ST.scala 32:46]
  assign _GEN_900 = 9'h19f == RADDR ? 9'h19f : _GEN_899; // @[RAM_ST.scala 32:46]
  assign _GEN_901 = 9'h1a0 == RADDR ? 9'h1a0 : _GEN_900; // @[RAM_ST.scala 32:46]
  assign _GEN_902 = 9'h1a1 == RADDR ? 9'h1a1 : _GEN_901; // @[RAM_ST.scala 32:46]
  assign _GEN_903 = 9'h1a2 == RADDR ? 9'h1a2 : _GEN_902; // @[RAM_ST.scala 32:46]
  assign _GEN_904 = 9'h1a3 == RADDR ? 9'h1a3 : _GEN_903; // @[RAM_ST.scala 32:46]
  assign _GEN_905 = 9'h1a4 == RADDR ? 9'h1a4 : _GEN_904; // @[RAM_ST.scala 32:46]
  assign _GEN_906 = 9'h1a5 == RADDR ? 9'h1a5 : _GEN_905; // @[RAM_ST.scala 32:46]
  assign _GEN_907 = 9'h1a6 == RADDR ? 9'h1a6 : _GEN_906; // @[RAM_ST.scala 32:46]
  assign _GEN_908 = 9'h1a7 == RADDR ? 9'h1a7 : _GEN_907; // @[RAM_ST.scala 32:46]
  assign _GEN_909 = 9'h1a8 == RADDR ? 9'h1a8 : _GEN_908; // @[RAM_ST.scala 32:46]
  assign _GEN_910 = 9'h1a9 == RADDR ? 9'h1a9 : _GEN_909; // @[RAM_ST.scala 32:46]
  assign _GEN_911 = 9'h1aa == RADDR ? 9'h1aa : _GEN_910; // @[RAM_ST.scala 32:46]
  assign _GEN_912 = 9'h1ab == RADDR ? 9'h1ab : _GEN_911; // @[RAM_ST.scala 32:46]
  assign _GEN_913 = 9'h1ac == RADDR ? 9'h1ac : _GEN_912; // @[RAM_ST.scala 32:46]
  assign _GEN_914 = 9'h1ad == RADDR ? 9'h1ad : _GEN_913; // @[RAM_ST.scala 32:46]
  assign _GEN_915 = 9'h1ae == RADDR ? 9'h1ae : _GEN_914; // @[RAM_ST.scala 32:46]
  assign _GEN_916 = 9'h1af == RADDR ? 9'h1af : _GEN_915; // @[RAM_ST.scala 32:46]
  assign _GEN_917 = 9'h1b0 == RADDR ? 9'h1b0 : _GEN_916; // @[RAM_ST.scala 32:46]
  assign _GEN_918 = 9'h1b1 == RADDR ? 9'h1b1 : _GEN_917; // @[RAM_ST.scala 32:46]
  assign _GEN_919 = 9'h1b2 == RADDR ? 9'h1b2 : _GEN_918; // @[RAM_ST.scala 32:46]
  assign _GEN_920 = 9'h1b3 == RADDR ? 9'h1b3 : _GEN_919; // @[RAM_ST.scala 32:46]
  assign _GEN_921 = 9'h1b4 == RADDR ? 9'h1b4 : _GEN_920; // @[RAM_ST.scala 32:46]
  assign _GEN_922 = 9'h1b5 == RADDR ? 9'h1b5 : _GEN_921; // @[RAM_ST.scala 32:46]
  assign _GEN_923 = 9'h1b6 == RADDR ? 9'h1b6 : _GEN_922; // @[RAM_ST.scala 32:46]
  assign _GEN_924 = 9'h1b7 == RADDR ? 9'h1b7 : _GEN_923; // @[RAM_ST.scala 32:46]
  assign _GEN_925 = 9'h1b8 == RADDR ? 9'h1b8 : _GEN_924; // @[RAM_ST.scala 32:46]
  assign _GEN_926 = 9'h1b9 == RADDR ? 9'h1b9 : _GEN_925; // @[RAM_ST.scala 32:46]
  assign _GEN_927 = 9'h1ba == RADDR ? 9'h1ba : _GEN_926; // @[RAM_ST.scala 32:46]
  assign _GEN_928 = 9'h1bb == RADDR ? 9'h1bb : _GEN_927; // @[RAM_ST.scala 32:46]
  assign _GEN_929 = 9'h1bc == RADDR ? 9'h1bc : _GEN_928; // @[RAM_ST.scala 32:46]
  assign _GEN_930 = 9'h1bd == RADDR ? 9'h1bd : _GEN_929; // @[RAM_ST.scala 32:46]
  assign _GEN_931 = 9'h1be == RADDR ? 9'h1be : _GEN_930; // @[RAM_ST.scala 32:46]
  assign _GEN_932 = 9'h1bf == RADDR ? 9'h1bf : _GEN_931; // @[RAM_ST.scala 32:46]
  assign _GEN_933 = 9'h1c0 == RADDR ? 9'h1c0 : _GEN_932; // @[RAM_ST.scala 32:46]
  assign _GEN_934 = 9'h1c1 == RADDR ? 9'h1c1 : _GEN_933; // @[RAM_ST.scala 32:46]
  assign _GEN_935 = 9'h1c2 == RADDR ? 9'h1c2 : _GEN_934; // @[RAM_ST.scala 32:46]
  assign _GEN_936 = 9'h1c3 == RADDR ? 9'h1c3 : _GEN_935; // @[RAM_ST.scala 32:46]
  assign _GEN_937 = 9'h1c4 == RADDR ? 9'h1c4 : _GEN_936; // @[RAM_ST.scala 32:46]
  assign _GEN_938 = 9'h1c5 == RADDR ? 9'h1c5 : _GEN_937; // @[RAM_ST.scala 32:46]
  assign _GEN_939 = 9'h1c6 == RADDR ? 9'h1c6 : _GEN_938; // @[RAM_ST.scala 32:46]
  assign _GEN_940 = 9'h1c7 == RADDR ? 9'h1c7 : _GEN_939; // @[RAM_ST.scala 32:46]
  assign _GEN_941 = 9'h1c8 == RADDR ? 9'h1c8 : _GEN_940; // @[RAM_ST.scala 32:46]
  assign _GEN_942 = 9'h1c9 == RADDR ? 9'h1c9 : _GEN_941; // @[RAM_ST.scala 32:46]
  assign _GEN_943 = 9'h1ca == RADDR ? 9'h1ca : _GEN_942; // @[RAM_ST.scala 32:46]
  assign _GEN_944 = 9'h1cb == RADDR ? 9'h1cb : _GEN_943; // @[RAM_ST.scala 32:46]
  assign _GEN_945 = 9'h1cc == RADDR ? 9'h1cc : _GEN_944; // @[RAM_ST.scala 32:46]
  assign _GEN_946 = 9'h1cd == RADDR ? 9'h1cd : _GEN_945; // @[RAM_ST.scala 32:46]
  assign _GEN_947 = 9'h1ce == RADDR ? 9'h1ce : _GEN_946; // @[RAM_ST.scala 32:46]
  assign _GEN_948 = 9'h1cf == RADDR ? 9'h1cf : _GEN_947; // @[RAM_ST.scala 32:46]
  assign _GEN_949 = 9'h1d0 == RADDR ? 9'h1d0 : _GEN_948; // @[RAM_ST.scala 32:46]
  assign _GEN_950 = 9'h1d1 == RADDR ? 9'h1d1 : _GEN_949; // @[RAM_ST.scala 32:46]
  assign _GEN_951 = 9'h1d2 == RADDR ? 9'h1d2 : _GEN_950; // @[RAM_ST.scala 32:46]
  assign _GEN_952 = 9'h1d3 == RADDR ? 9'h1d3 : _GEN_951; // @[RAM_ST.scala 32:46]
  assign _GEN_953 = 9'h1d4 == RADDR ? 9'h1d4 : _GEN_952; // @[RAM_ST.scala 32:46]
  assign _GEN_954 = 9'h1d5 == RADDR ? 9'h1d5 : _GEN_953; // @[RAM_ST.scala 32:46]
  assign _GEN_955 = 9'h1d6 == RADDR ? 9'h1d6 : _GEN_954; // @[RAM_ST.scala 32:46]
  assign _GEN_956 = 9'h1d7 == RADDR ? 9'h1d7 : _GEN_955; // @[RAM_ST.scala 32:46]
  assign _GEN_957 = 9'h1d8 == RADDR ? 9'h1d8 : _GEN_956; // @[RAM_ST.scala 32:46]
  assign _GEN_958 = 9'h1d9 == RADDR ? 9'h1d9 : _GEN_957; // @[RAM_ST.scala 32:46]
  assign _GEN_959 = 9'h1da == RADDR ? 9'h1da : _GEN_958; // @[RAM_ST.scala 32:46]
  assign _GEN_960 = 9'h1db == RADDR ? 9'h1db : _GEN_959; // @[RAM_ST.scala 32:46]
  assign _GEN_961 = 9'h1dc == RADDR ? 9'h1dc : _GEN_960; // @[RAM_ST.scala 32:46]
  assign _GEN_962 = 9'h1dd == RADDR ? 9'h1dd : _GEN_961; // @[RAM_ST.scala 32:46]
  assign _GEN_963 = 9'h1de == RADDR ? 9'h1de : _GEN_962; // @[RAM_ST.scala 32:46]
  assign _GEN_964 = 9'h1df == RADDR ? 9'h1df : _GEN_963; // @[RAM_ST.scala 32:46]
  assign _T_6 = {{1'd0}, _GEN_964}; // @[RAM_ST.scala 32:46]
  assign _T_13 = ram__T_11_data;
  assign RDATA_0 = _T_13[15:0]; // @[RAM_ST.scala 32:9]
  assign RDATA_1 = _T_13[31:16]; // @[RAM_ST.scala 32:9]
  assign RDATA_2 = _T_13[47:32]; // @[RAM_ST.scala 32:9]
  assign RDATA_3 = _T_13[63:48]; // @[RAM_ST.scala 32:9]
  assign write_elem_counter_CE = WE; // @[RAM_ST.scala 23:25]
  assign read_elem_counter_CE = RE; // @[RAM_ST.scala 24:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 480; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram__T_11_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ram__T_11_addr_pipe_0 = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_5_en & ram__T_5_mask) begin
      ram[ram__T_5_addr] <= ram__T_5_data; // @[RAM_ST.scala 29:24]
    end
    ram__T_11_en_pipe_0 <= read_elem_counter_valid;
    if (read_elem_counter_valid) begin
      ram__T_11_addr_pipe_0 <= _T_6[8:0];
    end
  end
endmodule
module ShiftT(
  input         clock,
  input         reset,
  input         valid_up,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  input  [15:0] I_3,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3
);
  wire  RAM_ST_clock; // @[ShiftT.scala 39:29]
  wire  RAM_ST_RE; // @[ShiftT.scala 39:29]
  wire [8:0] RAM_ST_RADDR; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_RDATA_0; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_RDATA_1; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_RDATA_2; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_RDATA_3; // @[ShiftT.scala 39:29]
  wire  RAM_ST_WE; // @[ShiftT.scala 39:29]
  wire [8:0] RAM_ST_WADDR; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_WDATA_0; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_WDATA_1; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_WDATA_2; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_WDATA_3; // @[ShiftT.scala 39:29]
  wire  NestedCounters_CE; // @[ShiftT.scala 41:31]
  wire  NestedCounters_valid; // @[ShiftT.scala 41:31]
  reg [8:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[Counter.scala 37:24]
  wire [8:0] _T_3; // @[Counter.scala 38:22]
  RAM_ST RAM_ST ( // @[ShiftT.scala 39:29]
    .clock(RAM_ST_clock),
    .RE(RAM_ST_RE),
    .RADDR(RAM_ST_RADDR),
    .RDATA_0(RAM_ST_RDATA_0),
    .RDATA_1(RAM_ST_RDATA_1),
    .RDATA_2(RAM_ST_RDATA_2),
    .RDATA_3(RAM_ST_RDATA_3),
    .WE(RAM_ST_WE),
    .WADDR(RAM_ST_WADDR),
    .WDATA_0(RAM_ST_WDATA_0),
    .WDATA_1(RAM_ST_WDATA_1),
    .WDATA_2(RAM_ST_WDATA_2),
    .WDATA_3(RAM_ST_WDATA_3)
  );
  NestedCounters_1 NestedCounters ( // @[ShiftT.scala 41:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign _T_1 = value == 9'h1df; // @[Counter.scala 37:24]
  assign _T_3 = value + 9'h1; // @[Counter.scala 38:22]
  assign O_0 = RAM_ST_RDATA_0; // @[ShiftT.scala 51:7]
  assign O_1 = RAM_ST_RDATA_1; // @[ShiftT.scala 51:7]
  assign O_2 = RAM_ST_RDATA_2; // @[ShiftT.scala 51:7]
  assign O_3 = RAM_ST_RDATA_3; // @[ShiftT.scala 51:7]
  assign RAM_ST_clock = clock;
  assign RAM_ST_RE = valid_up; // @[ShiftT.scala 49:20]
  assign RAM_ST_RADDR = _T_1 ? 9'h0 : _T_3; // @[ShiftT.scala 46:76 ShiftT.scala 47:38]
  assign RAM_ST_WE = valid_up; // @[ShiftT.scala 48:20]
  assign RAM_ST_WADDR = value; // @[ShiftT.scala 45:23]
  assign RAM_ST_WDATA_0 = I_0; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_1 = I_1; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_2 = I_2; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_3 = I_3; // @[ShiftT.scala 50:23]
  assign NestedCounters_CE = valid_up; // @[ShiftT.scala 42:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 9'h0;
    end else if (valid_up) begin
      if (_T_1) begin
        value <= 9'h0;
      end else begin
        value <= _T_3;
      end
    end
  end
endmodule
module ShiftTS(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  input  [15:0] I_3,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:26]
  wire  ShiftT_reset; // @[ShiftTS.scala 32:26]
  wire  ShiftT_valid_up; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_I_0; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_I_1; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_I_2; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_I_3; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_O_0; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_O_1; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_O_2; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_O_3; // @[ShiftTS.scala 32:26]
  ShiftT ShiftT ( // @[ShiftTS.scala 32:26]
    .clock(ShiftT_clock),
    .reset(ShiftT_reset),
    .valid_up(ShiftT_valid_up),
    .I_0(ShiftT_I_0),
    .I_1(ShiftT_I_1),
    .I_2(ShiftT_I_2),
    .I_3(ShiftT_I_3),
    .O_0(ShiftT_O_0),
    .O_1(ShiftT_O_1),
    .O_2(ShiftT_O_2),
    .O_3(ShiftT_O_3)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 58:14]
  assign O_0 = ShiftT_O_0; // @[ShiftTS.scala 51:36]
  assign O_1 = ShiftT_O_1; // @[ShiftTS.scala 51:36]
  assign O_2 = ShiftT_O_2; // @[ShiftTS.scala 51:36]
  assign O_3 = ShiftT_O_3; // @[ShiftTS.scala 51:36]
  assign ShiftT_clock = clock;
  assign ShiftT_reset = reset;
  assign ShiftT_valid_up = valid_up; // @[ShiftTS.scala 53:29]
  assign ShiftT_I_0 = I_0; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_1 = I_1; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_2 = I_2; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_3 = I_3; // @[ShiftTS.scala 50:25]
endmodule
module ShiftT_2(
  input         clock,
  input  [15:0] I_0,
  output [15:0] O_0
);
  reg [15:0] _T_0; // @[ShiftT.scala 24:82]
  reg [31:0] _RAND_0;
  assign O_0 = _T_0; // @[ShiftT.scala 24:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= I_0;
  end
endmodule
module ShiftTS_2(
  input         clock,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  input  [15:0] I_3,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_I_0; // @[ShiftTS.scala 32:26]
  wire [15:0] ShiftT_O_0; // @[ShiftTS.scala 32:26]
  ShiftT_2 ShiftT ( // @[ShiftTS.scala 32:26]
    .clock(ShiftT_clock),
    .I_0(ShiftT_I_0),
    .O_0(ShiftT_O_0)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 58:14]
  assign O_0 = ShiftT_O_0; // @[ShiftTS.scala 51:36]
  assign O_1 = I_0; // @[ShiftTS.scala 40:36]
  assign O_2 = I_1; // @[ShiftTS.scala 40:36]
  assign O_3 = I_2; // @[ShiftTS.scala 40:36]
  assign ShiftT_clock = clock;
  assign ShiftT_I_0 = I_3; // @[ShiftTS.scala 50:25]
endmodule
module SSeqTupleCreator(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0,
  input  [15:0] I1,
  output [15:0] O_0,
  output [15:0] O_1
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0 = I0; // @[Tuple.scala 12:32]
  assign O_1 = I1; // @[Tuple.scala 13:32]
endmodule
module Map2S(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I0_2,
  input  [15:0] I0_3,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  input  [15:0] I1_3,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_3_0,
  output [15:0] O_3_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  SSeqTupleCreator fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  SSeqTupleCreator other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1)
  );
  SSeqTupleCreator other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1)
  );
  SSeqTupleCreator other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0(other_ops_2_I0),
    .I1(other_ops_2_I1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign O_2_0 = other_ops_1_O_0; // @[Map2S.scala 24:12]
  assign O_2_1 = other_ops_1_O_1; // @[Map2S.scala 24:12]
  assign O_3_0 = other_ops_2_O_0; // @[Map2S.scala 24:12]
  assign O_3_1 = other_ops_2_O_1; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0 = I0_3; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
endmodule
module Map2T(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I0_2,
  input  [15:0] I0_3,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  input  [15:0] I1_3,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_3_0,
  output [15:0] O_3_1
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1; // @[Map2T.scala 8:20]
  Map2S op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I0_2(op_I0_2),
    .I0_3(op_I0_3),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign O_1_0 = op_O_1_0; // @[Map2T.scala 17:7]
  assign O_1_1 = op_O_1_1; // @[Map2T.scala 17:7]
  assign O_2_0 = op_O_2_0; // @[Map2T.scala 17:7]
  assign O_2_1 = op_O_2_1; // @[Map2T.scala 17:7]
  assign O_3_0 = op_O_3_0; // @[Map2T.scala 17:7]
  assign O_3_1 = op_O_3_1; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I0_2 = I0_2; // @[Map2T.scala 15:11]
  assign op_I0_3 = I0_3; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I1,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0 = I0_0; // @[Tuple.scala 24:34]
  assign O_1 = I0_1; // @[Tuple.scala 24:34]
  assign O_2 = I1; // @[Tuple.scala 26:32]
endmodule
module Map2S_1(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_3_0,
  input  [15:0] I0_3_1,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  input  [15:0] I1_3,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_3_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  SSeqTupleAppender fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  SSeqTupleAppender other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  SSeqTupleAppender other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I1(other_ops_1_I1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  SSeqTupleAppender other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I1(other_ops_2_I1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1),
    .O_2(other_ops_2_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_0_2 = fst_op_O_2; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign O_1_2 = other_ops_0_O_2; // @[Map2S.scala 24:12]
  assign O_2_0 = other_ops_1_O_0; // @[Map2S.scala 24:12]
  assign O_2_1 = other_ops_1_O_1; // @[Map2S.scala 24:12]
  assign O_2_2 = other_ops_1_O_2; // @[Map2S.scala 24:12]
  assign O_3_0 = other_ops_2_O_0; // @[Map2S.scala 24:12]
  assign O_3_1 = other_ops_2_O_1; // @[Map2S.scala 24:12]
  assign O_3_2 = other_ops_2_O_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
endmodule
module Map2T_1(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_3_0,
  input  [15:0] I0_3_1,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  input  [15:0] I1_3,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_3_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_2; // @[Map2T.scala 8:20]
  Map2S_1 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I0_2_0(op_I0_2_0),
    .I0_2_1(op_I0_2_1),
    .I0_3_0(op_I0_3_0),
    .I0_3_1(op_I0_3_1),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_0_2(op_O_0_2),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_1_2(op_O_1_2),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_2_2(op_O_2_2),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_3_2(op_O_3_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign O_0_2 = op_O_0_2; // @[Map2T.scala 17:7]
  assign O_1_0 = op_O_1_0; // @[Map2T.scala 17:7]
  assign O_1_1 = op_O_1_1; // @[Map2T.scala 17:7]
  assign O_1_2 = op_O_1_2; // @[Map2T.scala 17:7]
  assign O_2_0 = op_O_2_0; // @[Map2T.scala 17:7]
  assign O_2_1 = op_O_2_1; // @[Map2T.scala 17:7]
  assign O_2_2 = op_O_2_2; // @[Map2T.scala 17:7]
  assign O_3_0 = op_O_3_0; // @[Map2T.scala 17:7]
  assign O_3_1 = op_O_3_1; // @[Map2T.scala 17:7]
  assign O_3_2 = op_O_3_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0 = I0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1 = I0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0 = I0_3_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1 = I0_3_1; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
endmodule
module PartitionS(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  input  [15:0] I_3_0,
  input  [15:0] I_3_1,
  input  [15:0] I_3_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0 = I_0_0; // @[Partition.scala 15:39]
  assign O_0_0_1 = I_0_1; // @[Partition.scala 15:39]
  assign O_0_0_2 = I_0_2; // @[Partition.scala 15:39]
  assign O_1_0_0 = I_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1 = I_1_1; // @[Partition.scala 15:39]
  assign O_1_0_2 = I_1_2; // @[Partition.scala 15:39]
  assign O_2_0_0 = I_2_0; // @[Partition.scala 15:39]
  assign O_2_0_1 = I_2_1; // @[Partition.scala 15:39]
  assign O_2_0_2 = I_2_2; // @[Partition.scala 15:39]
  assign O_3_0_0 = I_3_0; // @[Partition.scala 15:39]
  assign O_3_0_1 = I_3_1; // @[Partition.scala 15:39]
  assign O_3_0_2 = I_3_2; // @[Partition.scala 15:39]
endmodule
module MapT(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  input  [15:0] I_3_0,
  input  [15:0] I_3_1,
  input  [15:0] I_3_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_2; // @[MapT.scala 8:20]
  PartitionS op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0(op_I_0_0),
    .I_0_1(op_I_0_1),
    .I_0_2(op_I_0_2),
    .I_1_0(op_I_1_0),
    .I_1_1(op_I_1_1),
    .I_1_2(op_I_1_2),
    .I_2_0(op_I_2_0),
    .I_2_1(op_I_2_1),
    .I_2_2(op_I_2_2),
    .I_3_0(op_I_3_0),
    .I_3_1(op_I_3_1),
    .I_3_2(op_I_3_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0 = I_0_0; // @[MapT.scala 14:10]
  assign op_I_0_1 = I_0_1; // @[MapT.scala 14:10]
  assign op_I_0_2 = I_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0 = I_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1 = I_1_1; // @[MapT.scala 14:10]
  assign op_I_1_2 = I_1_2; // @[MapT.scala 14:10]
  assign op_I_2_0 = I_2_0; // @[MapT.scala 14:10]
  assign op_I_2_1 = I_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2 = I_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0 = I_3_0; // @[MapT.scala 14:10]
  assign op_I_3_1 = I_3_1; // @[MapT.scala 14:10]
  assign op_I_3_2 = I_3_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0 = I_0; // @[Tuple.scala 41:5]
  assign O_1 = I_1; // @[Tuple.scala 41:5]
  assign O_2 = I_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0(op_inst_I_0),
    .I_1(op_inst_I_1),
    .I_2(op_inst_I_2),
    .O_0(op_inst_O_0),
    .O_1(op_inst_O_1),
    .O_2(op_inst_O_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0 = op_inst_O_0; // @[Remove1S.scala 14:5]
  assign O_1 = op_inst_O_1; // @[Remove1S.scala 14:5]
  assign O_2 = op_inst_O_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0 = I_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1 = I_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2 = I_0_2; // @[Remove1S.scala 13:13]
endmodule
module MapS(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_3_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  Remove1S fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  Remove1S other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  Remove1S other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  Remove1S other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1),
    .O_2(other_ops_2_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign O_3_0 = other_ops_2_O_0; // @[MapS.scala 21:12]
  assign O_3_1 = other_ops_2_O_1; // @[MapS.scala 21:12]
  assign O_3_2 = other_ops_2_O_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
endmodule
module MapT_1(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_3_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_2; // @[MapT.scala 8:20]
  MapS op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_0_2(op_O_0_2),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_1_2(op_O_1_2),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_2_2(op_O_2_2),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_3_2(op_O_3_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0 = op_O_0_0; // @[MapT.scala 15:7]
  assign O_0_1 = op_O_0_1; // @[MapT.scala 15:7]
  assign O_0_2 = op_O_0_2; // @[MapT.scala 15:7]
  assign O_1_0 = op_O_1_0; // @[MapT.scala 15:7]
  assign O_1_1 = op_O_1_1; // @[MapT.scala 15:7]
  assign O_1_2 = op_O_1_2; // @[MapT.scala 15:7]
  assign O_2_0 = op_O_2_0; // @[MapT.scala 15:7]
  assign O_2_1 = op_O_2_1; // @[MapT.scala 15:7]
  assign O_2_2 = op_O_2_2; // @[MapT.scala 15:7]
  assign O_3_0 = op_O_3_0; // @[MapT.scala 15:7]
  assign O_3_1 = op_O_3_1; // @[MapT.scala 15:7]
  assign O_3_2 = op_O_3_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleCreator_2(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I0_2,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0_0 = I0_0; // @[Tuple.scala 12:32]
  assign O_0_1 = I0_1; // @[Tuple.scala 12:32]
  assign O_0_2 = I0_2; // @[Tuple.scala 12:32]
  assign O_1_0 = I1_0; // @[Tuple.scala 13:32]
  assign O_1_1 = I1_1; // @[Tuple.scala 13:32]
  assign O_1_2 = I1_2; // @[Tuple.scala 13:32]
endmodule
module Map2S_4(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_0_2,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_1_2,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_2_2,
  input  [15:0] I0_3_0,
  input  [15:0] I0_3_1,
  input  [15:0] I0_3_2,
  input  [15:0] I1_0_0,
  input  [15:0] I1_0_1,
  input  [15:0] I1_0_2,
  input  [15:0] I1_1_0,
  input  [15:0] I1_1_1,
  input  [15:0] I1_1_2,
  input  [15:0] I1_2_0,
  input  [15:0] I1_2_1,
  input  [15:0] I1_2_2,
  input  [15:0] I1_3_0,
  input  [15:0] I1_3_1,
  input  [15:0] I1_3_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  SSeqTupleCreator_2 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I0_2(other_ops_2_I0_2),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .I1_2(other_ops_2_I1_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = I1_2_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_2 = I0_3_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_2 = I1_3_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_4(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_0_2,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_1_2,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_2_2,
  input  [15:0] I0_3_0,
  input  [15:0] I0_3_1,
  input  [15:0] I0_3_2,
  input  [15:0] I1_0_0,
  input  [15:0] I1_0_1,
  input  [15:0] I1_0_2,
  input  [15:0] I1_1_0,
  input  [15:0] I1_1_1,
  input  [15:0] I1_1_2,
  input  [15:0] I1_2_0,
  input  [15:0] I1_2_1,
  input  [15:0] I1_2_2,
  input  [15:0] I1_3_0,
  input  [15:0] I1_3_1,
  input  [15:0] I1_3_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_2; // @[Map2T.scala 8:20]
  Map2S_4 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_0_2(op_I0_0_2),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I0_1_2(op_I0_1_2),
    .I0_2_0(op_I0_2_0),
    .I0_2_1(op_I0_2_1),
    .I0_2_2(op_I0_2_2),
    .I0_3_0(op_I0_3_0),
    .I0_3_1(op_I0_3_1),
    .I0_3_2(op_I0_3_2),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_0_2(op_I1_0_2),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_1_2(op_I1_1_2),
    .I1_2_0(op_I1_2_0),
    .I1_2_1(op_I1_2_1),
    .I1_2_2(op_I1_2_2),
    .I1_3_0(op_I1_3_0),
    .I1_3_1(op_I1_3_1),
    .I1_3_2(op_I1_3_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_2 = op_O_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_1_2 = op_O_0_1_2; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_2 = op_O_1_0_2; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_1_1_2 = op_O_1_1_2; // @[Map2T.scala 17:7]
  assign O_2_0_0 = op_O_2_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_1 = op_O_2_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_2 = op_O_2_0_2; // @[Map2T.scala 17:7]
  assign O_2_1_0 = op_O_2_1_0; // @[Map2T.scala 17:7]
  assign O_2_1_1 = op_O_2_1_1; // @[Map2T.scala 17:7]
  assign O_2_1_2 = op_O_2_1_2; // @[Map2T.scala 17:7]
  assign O_3_0_0 = op_O_3_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_1 = op_O_3_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_2 = op_O_3_0_2; // @[Map2T.scala 17:7]
  assign O_3_1_0 = op_O_3_1_0; // @[Map2T.scala 17:7]
  assign O_3_1_1 = op_O_3_1_1; // @[Map2T.scala 17:7]
  assign O_3_1_2 = op_O_3_1_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_2 = I0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_2 = I0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0 = I0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1 = I0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_2_2 = I0_2_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0 = I0_3_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1 = I0_3_1; // @[Map2T.scala 15:11]
  assign op_I0_3_2 = I0_3_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_2 = I1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_1_2 = I1_1_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0 = I1_2_0; // @[Map2T.scala 16:11]
  assign op_I1_2_1 = I1_2_1; // @[Map2T.scala 16:11]
  assign op_I1_2_2 = I1_2_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0 = I1_3_0; // @[Map2T.scala 16:11]
  assign op_I1_3_1 = I1_3_1; // @[Map2T.scala 16:11]
  assign op_I1_3_2 = I1_3_2; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender_3(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_0_2,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_1_2,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0_0 = I0_0_0; // @[Tuple.scala 24:34]
  assign O_0_1 = I0_0_1; // @[Tuple.scala 24:34]
  assign O_0_2 = I0_0_2; // @[Tuple.scala 24:34]
  assign O_1_0 = I0_1_0; // @[Tuple.scala 24:34]
  assign O_1_1 = I0_1_1; // @[Tuple.scala 24:34]
  assign O_1_2 = I0_1_2; // @[Tuple.scala 24:34]
  assign O_2_0 = I1_0; // @[Tuple.scala 26:32]
  assign O_2_1 = I1_1; // @[Tuple.scala 26:32]
  assign O_2_2 = I1_2; // @[Tuple.scala 26:32]
endmodule
module Map2S_7(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0_0,
  input  [15:0] I0_0_0_1,
  input  [15:0] I0_0_0_2,
  input  [15:0] I0_0_1_0,
  input  [15:0] I0_0_1_1,
  input  [15:0] I0_0_1_2,
  input  [15:0] I0_1_0_0,
  input  [15:0] I0_1_0_1,
  input  [15:0] I0_1_0_2,
  input  [15:0] I0_1_1_0,
  input  [15:0] I0_1_1_1,
  input  [15:0] I0_1_1_2,
  input  [15:0] I0_2_0_0,
  input  [15:0] I0_2_0_1,
  input  [15:0] I0_2_0_2,
  input  [15:0] I0_2_1_0,
  input  [15:0] I0_2_1_1,
  input  [15:0] I0_2_1_2,
  input  [15:0] I0_3_0_0,
  input  [15:0] I0_3_0_1,
  input  [15:0] I0_3_0_2,
  input  [15:0] I0_3_1_0,
  input  [15:0] I0_3_1_1,
  input  [15:0] I0_3_1_2,
  input  [15:0] I1_0_0,
  input  [15:0] I1_0_1,
  input  [15:0] I1_0_2,
  input  [15:0] I1_1_0,
  input  [15:0] I1_1_1,
  input  [15:0] I1_1_2,
  input  [15:0] I1_2_0,
  input  [15:0] I1_2_1,
  input  [15:0] I1_2_2,
  input  [15:0] I1_3_0,
  input  [15:0] I1_3_1,
  input  [15:0] I1_3_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_0_2_0,
  output [15:0] O_0_2_1,
  output [15:0] O_0_2_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_1_2_0,
  output [15:0] O_1_2_1,
  output [15:0] O_1_2_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_2_2_0,
  output [15:0] O_2_2_1,
  output [15:0] O_2_2_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_3_2_0,
  output [15:0] O_3_2_1,
  output [15:0] O_3_2_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_2_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  SSeqTupleAppender_3 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I0_1_0(fst_op_I0_1_0),
    .I0_1_1(fst_op_I0_1_1),
    .I0_1_2(fst_op_I0_1_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0(other_ops_0_I0_0_0),
    .I0_0_1(other_ops_0_I0_0_1),
    .I0_0_2(other_ops_0_I0_0_2),
    .I0_1_0(other_ops_0_I0_1_0),
    .I0_1_1(other_ops_0_I0_1_1),
    .I0_1_2(other_ops_0_I0_1_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0(other_ops_1_I0_0_0),
    .I0_0_1(other_ops_1_I0_0_1),
    .I0_0_2(other_ops_1_I0_0_2),
    .I0_1_0(other_ops_1_I0_1_0),
    .I0_1_1(other_ops_1_I0_1_1),
    .I0_1_2(other_ops_1_I0_1_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0(other_ops_2_I0_0_0),
    .I0_0_1(other_ops_2_I0_0_1),
    .I0_0_2(other_ops_2_I0_0_2),
    .I0_1_0(other_ops_2_I0_1_0),
    .I0_1_1(other_ops_2_I0_1_1),
    .I0_1_2(other_ops_2_I0_1_2),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .I1_2(other_ops_2_I1_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[Map2S.scala 19:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[Map2S.scala 19:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[Map2S.scala 24:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[Map2S.scala 24:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[Map2S.scala 24:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[Map2S.scala 24:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[Map2S.scala 24:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[Map2S.scala 24:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[Map2S.scala 24:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[Map2S.scala 24:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_0 = I0_0_1_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_1 = I0_0_1_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_2 = I0_0_1_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0 = I0_1_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1 = I0_1_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_2 = I0_1_0_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_0 = I0_1_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_1 = I0_1_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_2 = I0_1_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0 = I0_2_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1 = I0_2_0_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_2 = I0_2_0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_0 = I0_2_1_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_1 = I0_2_1_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_2 = I0_2_1_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = I1_2_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0 = I0_3_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1 = I0_3_0_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_2 = I0_3_0_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_0 = I0_3_1_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_1 = I0_3_1_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_2 = I0_3_1_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_2 = I1_3_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_7(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0_0,
  input  [15:0] I0_0_0_1,
  input  [15:0] I0_0_0_2,
  input  [15:0] I0_0_1_0,
  input  [15:0] I0_0_1_1,
  input  [15:0] I0_0_1_2,
  input  [15:0] I0_1_0_0,
  input  [15:0] I0_1_0_1,
  input  [15:0] I0_1_0_2,
  input  [15:0] I0_1_1_0,
  input  [15:0] I0_1_1_1,
  input  [15:0] I0_1_1_2,
  input  [15:0] I0_2_0_0,
  input  [15:0] I0_2_0_1,
  input  [15:0] I0_2_0_2,
  input  [15:0] I0_2_1_0,
  input  [15:0] I0_2_1_1,
  input  [15:0] I0_2_1_2,
  input  [15:0] I0_3_0_0,
  input  [15:0] I0_3_0_1,
  input  [15:0] I0_3_0_2,
  input  [15:0] I0_3_1_0,
  input  [15:0] I0_3_1_1,
  input  [15:0] I0_3_1_2,
  input  [15:0] I1_0_0,
  input  [15:0] I1_0_1,
  input  [15:0] I1_0_2,
  input  [15:0] I1_1_0,
  input  [15:0] I1_1_1,
  input  [15:0] I1_1_2,
  input  [15:0] I1_2_0,
  input  [15:0] I1_2_1,
  input  [15:0] I1_2_2,
  input  [15:0] I1_3_0,
  input  [15:0] I1_3_1,
  input  [15:0] I1_3_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_0_2_0,
  output [15:0] O_0_2_1,
  output [15:0] O_0_2_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_1_2_0,
  output [15:0] O_1_2_1,
  output [15:0] O_1_2_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_2_2_0,
  output [15:0] O_2_2_1,
  output [15:0] O_2_2_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_3_2_0,
  output [15:0] O_3_2_1,
  output [15:0] O_3_2_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_2_2; // @[Map2T.scala 8:20]
  Map2S_7 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0(op_I0_0_0_0),
    .I0_0_0_1(op_I0_0_0_1),
    .I0_0_0_2(op_I0_0_0_2),
    .I0_0_1_0(op_I0_0_1_0),
    .I0_0_1_1(op_I0_0_1_1),
    .I0_0_1_2(op_I0_0_1_2),
    .I0_1_0_0(op_I0_1_0_0),
    .I0_1_0_1(op_I0_1_0_1),
    .I0_1_0_2(op_I0_1_0_2),
    .I0_1_1_0(op_I0_1_1_0),
    .I0_1_1_1(op_I0_1_1_1),
    .I0_1_1_2(op_I0_1_1_2),
    .I0_2_0_0(op_I0_2_0_0),
    .I0_2_0_1(op_I0_2_0_1),
    .I0_2_0_2(op_I0_2_0_2),
    .I0_2_1_0(op_I0_2_1_0),
    .I0_2_1_1(op_I0_2_1_1),
    .I0_2_1_2(op_I0_2_1_2),
    .I0_3_0_0(op_I0_3_0_0),
    .I0_3_0_1(op_I0_3_0_1),
    .I0_3_0_2(op_I0_3_0_2),
    .I0_3_1_0(op_I0_3_1_0),
    .I0_3_1_1(op_I0_3_1_1),
    .I0_3_1_2(op_I0_3_1_2),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_0_2(op_I1_0_2),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_1_2(op_I1_1_2),
    .I1_2_0(op_I1_2_0),
    .I1_2_1(op_I1_2_1),
    .I1_2_2(op_I1_2_2),
    .I1_3_0(op_I1_3_0),
    .I1_3_1(op_I1_3_1),
    .I1_3_2(op_I1_3_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_2_2_0(op_O_2_2_0),
    .O_2_2_1(op_O_2_2_1),
    .O_2_2_2(op_O_2_2_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_3_2_0(op_O_3_2_0),
    .O_3_2_1(op_O_3_2_1),
    .O_3_2_2(op_O_3_2_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_2 = op_O_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_1_2 = op_O_0_1_2; // @[Map2T.scala 17:7]
  assign O_0_2_0 = op_O_0_2_0; // @[Map2T.scala 17:7]
  assign O_0_2_1 = op_O_0_2_1; // @[Map2T.scala 17:7]
  assign O_0_2_2 = op_O_0_2_2; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_2 = op_O_1_0_2; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_1_1_2 = op_O_1_1_2; // @[Map2T.scala 17:7]
  assign O_1_2_0 = op_O_1_2_0; // @[Map2T.scala 17:7]
  assign O_1_2_1 = op_O_1_2_1; // @[Map2T.scala 17:7]
  assign O_1_2_2 = op_O_1_2_2; // @[Map2T.scala 17:7]
  assign O_2_0_0 = op_O_2_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_1 = op_O_2_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_2 = op_O_2_0_2; // @[Map2T.scala 17:7]
  assign O_2_1_0 = op_O_2_1_0; // @[Map2T.scala 17:7]
  assign O_2_1_1 = op_O_2_1_1; // @[Map2T.scala 17:7]
  assign O_2_1_2 = op_O_2_1_2; // @[Map2T.scala 17:7]
  assign O_2_2_0 = op_O_2_2_0; // @[Map2T.scala 17:7]
  assign O_2_2_1 = op_O_2_2_1; // @[Map2T.scala 17:7]
  assign O_2_2_2 = op_O_2_2_2; // @[Map2T.scala 17:7]
  assign O_3_0_0 = op_O_3_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_1 = op_O_3_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_2 = op_O_3_0_2; // @[Map2T.scala 17:7]
  assign O_3_1_0 = op_O_3_1_0; // @[Map2T.scala 17:7]
  assign O_3_1_1 = op_O_3_1_1; // @[Map2T.scala 17:7]
  assign O_3_1_2 = op_O_3_1_2; // @[Map2T.scala 17:7]
  assign O_3_2_0 = op_O_3_2_0; // @[Map2T.scala 17:7]
  assign O_3_2_1 = op_O_3_2_1; // @[Map2T.scala 17:7]
  assign O_3_2_2 = op_O_3_2_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0 = I0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1 = I0_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_0_2 = I0_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_0_1_0 = I0_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1_1 = I0_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_0_1_2 = I0_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0 = I0_1_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1 = I0_1_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_2 = I0_1_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_1_0 = I0_1_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1_1 = I0_1_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_1_2 = I0_1_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0 = I0_2_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1 = I0_2_0_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_2 = I0_2_0_2; // @[Map2T.scala 15:11]
  assign op_I0_2_1_0 = I0_2_1_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1_1 = I0_2_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_1_2 = I0_2_1_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0 = I0_3_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1 = I0_3_0_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_2 = I0_3_0_2; // @[Map2T.scala 15:11]
  assign op_I0_3_1_0 = I0_3_1_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1_1 = I0_3_1_1; // @[Map2T.scala 15:11]
  assign op_I0_3_1_2 = I0_3_1_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_2 = I1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_1_2 = I1_1_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0 = I1_2_0; // @[Map2T.scala 16:11]
  assign op_I1_2_1 = I1_2_1; // @[Map2T.scala 16:11]
  assign op_I1_2_2 = I1_2_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0 = I1_3_0; // @[Map2T.scala 16:11]
  assign op_I1_3_1 = I1_3_1; // @[Map2T.scala 16:11]
  assign op_I1_3_2 = I1_3_2; // @[Map2T.scala 16:11]
endmodule
module PartitionS_3(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_0_1_2,
  input  [15:0] I_0_2_0,
  input  [15:0] I_0_2_1,
  input  [15:0] I_0_2_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_1_1_2,
  input  [15:0] I_1_2_0,
  input  [15:0] I_1_2_1,
  input  [15:0] I_1_2_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_2_1_2,
  input  [15:0] I_2_2_0,
  input  [15:0] I_2_2_1,
  input  [15:0] I_2_2_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  input  [15:0] I_3_1_2,
  input  [15:0] I_3_2_0,
  input  [15:0] I_3_2_1,
  input  [15:0] I_3_2_2,
  output [15:0] O_0_0_0_0,
  output [15:0] O_0_0_0_1,
  output [15:0] O_0_0_0_2,
  output [15:0] O_0_0_1_0,
  output [15:0] O_0_0_1_1,
  output [15:0] O_0_0_1_2,
  output [15:0] O_0_0_2_0,
  output [15:0] O_0_0_2_1,
  output [15:0] O_0_0_2_2,
  output [15:0] O_1_0_0_0,
  output [15:0] O_1_0_0_1,
  output [15:0] O_1_0_0_2,
  output [15:0] O_1_0_1_0,
  output [15:0] O_1_0_1_1,
  output [15:0] O_1_0_1_2,
  output [15:0] O_1_0_2_0,
  output [15:0] O_1_0_2_1,
  output [15:0] O_1_0_2_2,
  output [15:0] O_2_0_0_0,
  output [15:0] O_2_0_0_1,
  output [15:0] O_2_0_0_2,
  output [15:0] O_2_0_1_0,
  output [15:0] O_2_0_1_1,
  output [15:0] O_2_0_1_2,
  output [15:0] O_2_0_2_0,
  output [15:0] O_2_0_2_1,
  output [15:0] O_2_0_2_2,
  output [15:0] O_3_0_0_0,
  output [15:0] O_3_0_0_1,
  output [15:0] O_3_0_0_2,
  output [15:0] O_3_0_1_0,
  output [15:0] O_3_0_1_1,
  output [15:0] O_3_0_1_2,
  output [15:0] O_3_0_2_0,
  output [15:0] O_3_0_2_1,
  output [15:0] O_3_0_2_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0_0 = I_0_0_0; // @[Partition.scala 15:39]
  assign O_0_0_0_1 = I_0_0_1; // @[Partition.scala 15:39]
  assign O_0_0_0_2 = I_0_0_2; // @[Partition.scala 15:39]
  assign O_0_0_1_0 = I_0_1_0; // @[Partition.scala 15:39]
  assign O_0_0_1_1 = I_0_1_1; // @[Partition.scala 15:39]
  assign O_0_0_1_2 = I_0_1_2; // @[Partition.scala 15:39]
  assign O_0_0_2_0 = I_0_2_0; // @[Partition.scala 15:39]
  assign O_0_0_2_1 = I_0_2_1; // @[Partition.scala 15:39]
  assign O_0_0_2_2 = I_0_2_2; // @[Partition.scala 15:39]
  assign O_1_0_0_0 = I_1_0_0; // @[Partition.scala 15:39]
  assign O_1_0_0_1 = I_1_0_1; // @[Partition.scala 15:39]
  assign O_1_0_0_2 = I_1_0_2; // @[Partition.scala 15:39]
  assign O_1_0_1_0 = I_1_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1_1 = I_1_1_1; // @[Partition.scala 15:39]
  assign O_1_0_1_2 = I_1_1_2; // @[Partition.scala 15:39]
  assign O_1_0_2_0 = I_1_2_0; // @[Partition.scala 15:39]
  assign O_1_0_2_1 = I_1_2_1; // @[Partition.scala 15:39]
  assign O_1_0_2_2 = I_1_2_2; // @[Partition.scala 15:39]
  assign O_2_0_0_0 = I_2_0_0; // @[Partition.scala 15:39]
  assign O_2_0_0_1 = I_2_0_1; // @[Partition.scala 15:39]
  assign O_2_0_0_2 = I_2_0_2; // @[Partition.scala 15:39]
  assign O_2_0_1_0 = I_2_1_0; // @[Partition.scala 15:39]
  assign O_2_0_1_1 = I_2_1_1; // @[Partition.scala 15:39]
  assign O_2_0_1_2 = I_2_1_2; // @[Partition.scala 15:39]
  assign O_2_0_2_0 = I_2_2_0; // @[Partition.scala 15:39]
  assign O_2_0_2_1 = I_2_2_1; // @[Partition.scala 15:39]
  assign O_2_0_2_2 = I_2_2_2; // @[Partition.scala 15:39]
  assign O_3_0_0_0 = I_3_0_0; // @[Partition.scala 15:39]
  assign O_3_0_0_1 = I_3_0_1; // @[Partition.scala 15:39]
  assign O_3_0_0_2 = I_3_0_2; // @[Partition.scala 15:39]
  assign O_3_0_1_0 = I_3_1_0; // @[Partition.scala 15:39]
  assign O_3_0_1_1 = I_3_1_1; // @[Partition.scala 15:39]
  assign O_3_0_1_2 = I_3_1_2; // @[Partition.scala 15:39]
  assign O_3_0_2_0 = I_3_2_0; // @[Partition.scala 15:39]
  assign O_3_0_2_1 = I_3_2_1; // @[Partition.scala 15:39]
  assign O_3_0_2_2 = I_3_2_2; // @[Partition.scala 15:39]
endmodule
module MapT_6(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_0_1_2,
  input  [15:0] I_0_2_0,
  input  [15:0] I_0_2_1,
  input  [15:0] I_0_2_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_1_1_2,
  input  [15:0] I_1_2_0,
  input  [15:0] I_1_2_1,
  input  [15:0] I_1_2_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_2_1_2,
  input  [15:0] I_2_2_0,
  input  [15:0] I_2_2_1,
  input  [15:0] I_2_2_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  input  [15:0] I_3_1_2,
  input  [15:0] I_3_2_0,
  input  [15:0] I_3_2_1,
  input  [15:0] I_3_2_2,
  output [15:0] O_0_0_0_0,
  output [15:0] O_0_0_0_1,
  output [15:0] O_0_0_0_2,
  output [15:0] O_0_0_1_0,
  output [15:0] O_0_0_1_1,
  output [15:0] O_0_0_1_2,
  output [15:0] O_0_0_2_0,
  output [15:0] O_0_0_2_1,
  output [15:0] O_0_0_2_2,
  output [15:0] O_1_0_0_0,
  output [15:0] O_1_0_0_1,
  output [15:0] O_1_0_0_2,
  output [15:0] O_1_0_1_0,
  output [15:0] O_1_0_1_1,
  output [15:0] O_1_0_1_2,
  output [15:0] O_1_0_2_0,
  output [15:0] O_1_0_2_1,
  output [15:0] O_1_0_2_2,
  output [15:0] O_2_0_0_0,
  output [15:0] O_2_0_0_1,
  output [15:0] O_2_0_0_2,
  output [15:0] O_2_0_1_0,
  output [15:0] O_2_0_1_1,
  output [15:0] O_2_0_1_2,
  output [15:0] O_2_0_2_0,
  output [15:0] O_2_0_2_1,
  output [15:0] O_2_0_2_2,
  output [15:0] O_3_0_0_0,
  output [15:0] O_3_0_0_1,
  output [15:0] O_3_0_0_2,
  output [15:0] O_3_0_1_0,
  output [15:0] O_3_0_1_1,
  output [15:0] O_3_0_1_2,
  output [15:0] O_3_0_2_0,
  output [15:0] O_3_0_2_1,
  output [15:0] O_3_0_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_2_2; // @[MapT.scala 8:20]
  PartitionS_3 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_0_0_0_2(op_O_0_0_0_2),
    .O_0_0_1_0(op_O_0_0_1_0),
    .O_0_0_1_1(op_O_0_0_1_1),
    .O_0_0_1_2(op_O_0_0_1_2),
    .O_0_0_2_0(op_O_0_0_2_0),
    .O_0_0_2_1(op_O_0_0_2_1),
    .O_0_0_2_2(op_O_0_0_2_2),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_1_0_0_2(op_O_1_0_0_2),
    .O_1_0_1_0(op_O_1_0_1_0),
    .O_1_0_1_1(op_O_1_0_1_1),
    .O_1_0_1_2(op_O_1_0_1_2),
    .O_1_0_2_0(op_O_1_0_2_0),
    .O_1_0_2_1(op_O_1_0_2_1),
    .O_1_0_2_2(op_O_1_0_2_2),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_2_0_0_2(op_O_2_0_0_2),
    .O_2_0_1_0(op_O_2_0_1_0),
    .O_2_0_1_1(op_O_2_0_1_1),
    .O_2_0_1_2(op_O_2_0_1_2),
    .O_2_0_2_0(op_O_2_0_2_0),
    .O_2_0_2_1(op_O_2_0_2_1),
    .O_2_0_2_2(op_O_2_0_2_2),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_3_0_0_2(op_O_3_0_0_2),
    .O_3_0_1_0(op_O_3_0_1_0),
    .O_3_0_1_1(op_O_3_0_1_1),
    .O_3_0_1_2(op_O_3_0_1_2),
    .O_3_0_2_0(op_O_3_0_2_0),
    .O_3_0_2_1(op_O_3_0_2_1),
    .O_3_0_2_2(op_O_3_0_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_0_2 = op_O_0_0_0_2; // @[MapT.scala 15:7]
  assign O_0_0_1_0 = op_O_0_0_1_0; // @[MapT.scala 15:7]
  assign O_0_0_1_1 = op_O_0_0_1_1; // @[MapT.scala 15:7]
  assign O_0_0_1_2 = op_O_0_0_1_2; // @[MapT.scala 15:7]
  assign O_0_0_2_0 = op_O_0_0_2_0; // @[MapT.scala 15:7]
  assign O_0_0_2_1 = op_O_0_0_2_1; // @[MapT.scala 15:7]
  assign O_0_0_2_2 = op_O_0_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[MapT.scala 15:7]
  assign O_1_0_0_2 = op_O_1_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_1_0 = op_O_1_0_1_0; // @[MapT.scala 15:7]
  assign O_1_0_1_1 = op_O_1_0_1_1; // @[MapT.scala 15:7]
  assign O_1_0_1_2 = op_O_1_0_1_2; // @[MapT.scala 15:7]
  assign O_1_0_2_0 = op_O_1_0_2_0; // @[MapT.scala 15:7]
  assign O_1_0_2_1 = op_O_1_0_2_1; // @[MapT.scala 15:7]
  assign O_1_0_2_2 = op_O_1_0_2_2; // @[MapT.scala 15:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[MapT.scala 15:7]
  assign O_2_0_0_2 = op_O_2_0_0_2; // @[MapT.scala 15:7]
  assign O_2_0_1_0 = op_O_2_0_1_0; // @[MapT.scala 15:7]
  assign O_2_0_1_1 = op_O_2_0_1_1; // @[MapT.scala 15:7]
  assign O_2_0_1_2 = op_O_2_0_1_2; // @[MapT.scala 15:7]
  assign O_2_0_2_0 = op_O_2_0_2_0; // @[MapT.scala 15:7]
  assign O_2_0_2_1 = op_O_2_0_2_1; // @[MapT.scala 15:7]
  assign O_2_0_2_2 = op_O_2_0_2_2; // @[MapT.scala 15:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[MapT.scala 15:7]
  assign O_3_0_0_2 = op_O_3_0_0_2; // @[MapT.scala 15:7]
  assign O_3_0_1_0 = op_O_3_0_1_0; // @[MapT.scala 15:7]
  assign O_3_0_1_1 = op_O_3_0_1_1; // @[MapT.scala 15:7]
  assign O_3_0_1_2 = op_O_3_0_1_2; // @[MapT.scala 15:7]
  assign O_3_0_2_0 = op_O_3_0_2_0; // @[MapT.scala 15:7]
  assign O_3_0_2_1 = op_O_3_0_2_1; // @[MapT.scala 15:7]
  assign O_3_0_2_2 = op_O_3_0_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq_3(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0_0 = I_0_0; // @[Tuple.scala 41:5]
  assign O_0_1 = I_0_1; // @[Tuple.scala 41:5]
  assign O_0_2 = I_0_2; // @[Tuple.scala 41:5]
  assign O_1_0 = I_1_0; // @[Tuple.scala 41:5]
  assign O_1_1 = I_1_1; // @[Tuple.scala 41:5]
  assign O_1_2 = I_1_2; // @[Tuple.scala 41:5]
  assign O_2_0 = I_2_0; // @[Tuple.scala 41:5]
  assign O_2_1 = I_2_1; // @[Tuple.scala 41:5]
  assign O_2_2 = I_2_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S_3(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_0_1_2,
  input  [15:0] I_0_2_0,
  input  [15:0] I_0_2_1,
  input  [15:0] I_0_2_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_0_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_0_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_0_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_1_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_1_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_1_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_2_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_2_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_2_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_0_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_0_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_0_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_1_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_1_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_1_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_2_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_2_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_2_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_3 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0_0(op_inst_I_0_0),
    .I_0_1(op_inst_I_0_1),
    .I_0_2(op_inst_I_0_2),
    .I_1_0(op_inst_I_1_0),
    .I_1_1(op_inst_I_1_1),
    .I_1_2(op_inst_I_1_2),
    .I_2_0(op_inst_I_2_0),
    .I_2_1(op_inst_I_2_1),
    .I_2_2(op_inst_I_2_2),
    .O_0_0(op_inst_O_0_0),
    .O_0_1(op_inst_O_0_1),
    .O_0_2(op_inst_O_0_2),
    .O_1_0(op_inst_O_1_0),
    .O_1_1(op_inst_O_1_1),
    .O_1_2(op_inst_O_1_2),
    .O_2_0(op_inst_O_2_0),
    .O_2_1(op_inst_O_2_1),
    .O_2_2(op_inst_O_2_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0_0 = op_inst_O_0_0; // @[Remove1S.scala 14:5]
  assign O_0_1 = op_inst_O_0_1; // @[Remove1S.scala 14:5]
  assign O_0_2 = op_inst_O_0_2; // @[Remove1S.scala 14:5]
  assign O_1_0 = op_inst_O_1_0; // @[Remove1S.scala 14:5]
  assign O_1_1 = op_inst_O_1_1; // @[Remove1S.scala 14:5]
  assign O_1_2 = op_inst_O_1_2; // @[Remove1S.scala 14:5]
  assign O_2_0 = op_inst_O_2_0; // @[Remove1S.scala 14:5]
  assign O_2_1 = op_inst_O_2_1; // @[Remove1S.scala 14:5]
  assign O_2_2 = op_inst_O_2_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0_0 = I_0_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_1 = I_0_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_2 = I_0_0_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_0 = I_0_1_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_1 = I_0_1_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_2 = I_0_1_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_0 = I_0_2_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_1 = I_0_2_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_2 = I_0_2_2; // @[Remove1S.scala 13:13]
endmodule
module MapS_3(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0_0,
  input  [15:0] I_0_0_0_1,
  input  [15:0] I_0_0_0_2,
  input  [15:0] I_0_0_1_0,
  input  [15:0] I_0_0_1_1,
  input  [15:0] I_0_0_1_2,
  input  [15:0] I_0_0_2_0,
  input  [15:0] I_0_0_2_1,
  input  [15:0] I_0_0_2_2,
  input  [15:0] I_1_0_0_0,
  input  [15:0] I_1_0_0_1,
  input  [15:0] I_1_0_0_2,
  input  [15:0] I_1_0_1_0,
  input  [15:0] I_1_0_1_1,
  input  [15:0] I_1_0_1_2,
  input  [15:0] I_1_0_2_0,
  input  [15:0] I_1_0_2_1,
  input  [15:0] I_1_0_2_2,
  input  [15:0] I_2_0_0_0,
  input  [15:0] I_2_0_0_1,
  input  [15:0] I_2_0_0_2,
  input  [15:0] I_2_0_1_0,
  input  [15:0] I_2_0_1_1,
  input  [15:0] I_2_0_1_2,
  input  [15:0] I_2_0_2_0,
  input  [15:0] I_2_0_2_1,
  input  [15:0] I_2_0_2_2,
  input  [15:0] I_3_0_0_0,
  input  [15:0] I_3_0_0_1,
  input  [15:0] I_3_0_0_2,
  input  [15:0] I_3_0_1_0,
  input  [15:0] I_3_0_1_1,
  input  [15:0] I_3_0_1_2,
  input  [15:0] I_3_0_2_0,
  input  [15:0] I_3_0_2_1,
  input  [15:0] I_3_0_2_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_0_2_0,
  output [15:0] O_0_2_1,
  output [15:0] O_0_2_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_1_2_0,
  output [15:0] O_1_2_1,
  output [15:0] O_1_2_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_2_2_0,
  output [15:0] O_2_2_1,
  output [15:0] O_2_2_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_3_2_0,
  output [15:0] O_3_2_1,
  output [15:0] O_3_2_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_2_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_2_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_2_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_2_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_2_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_2_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_2_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  Remove1S_3 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0_0(fst_op_I_0_0_0),
    .I_0_0_1(fst_op_I_0_0_1),
    .I_0_0_2(fst_op_I_0_0_2),
    .I_0_1_0(fst_op_I_0_1_0),
    .I_0_1_1(fst_op_I_0_1_1),
    .I_0_1_2(fst_op_I_0_1_2),
    .I_0_2_0(fst_op_I_0_2_0),
    .I_0_2_1(fst_op_I_0_2_1),
    .I_0_2_2(fst_op_I_0_2_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  Remove1S_3 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0_0(other_ops_0_I_0_0_0),
    .I_0_0_1(other_ops_0_I_0_0_1),
    .I_0_0_2(other_ops_0_I_0_0_2),
    .I_0_1_0(other_ops_0_I_0_1_0),
    .I_0_1_1(other_ops_0_I_0_1_1),
    .I_0_1_2(other_ops_0_I_0_1_2),
    .I_0_2_0(other_ops_0_I_0_2_0),
    .I_0_2_1(other_ops_0_I_0_2_1),
    .I_0_2_2(other_ops_0_I_0_2_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  Remove1S_3 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0_0(other_ops_1_I_0_0_0),
    .I_0_0_1(other_ops_1_I_0_0_1),
    .I_0_0_2(other_ops_1_I_0_0_2),
    .I_0_1_0(other_ops_1_I_0_1_0),
    .I_0_1_1(other_ops_1_I_0_1_1),
    .I_0_1_2(other_ops_1_I_0_1_2),
    .I_0_2_0(other_ops_1_I_0_2_0),
    .I_0_2_1(other_ops_1_I_0_2_1),
    .I_0_2_2(other_ops_1_I_0_2_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  Remove1S_3 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0_0(other_ops_2_I_0_0_0),
    .I_0_0_1(other_ops_2_I_0_0_1),
    .I_0_0_2(other_ops_2_I_0_0_2),
    .I_0_1_0(other_ops_2_I_0_1_0),
    .I_0_1_1(other_ops_2_I_0_1_1),
    .I_0_1_2(other_ops_2_I_0_1_2),
    .I_0_2_0(other_ops_2_I_0_2_0),
    .I_0_2_1(other_ops_2_I_0_2_1),
    .I_0_2_2(other_ops_2_I_0_2_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[MapS.scala 17:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[MapS.scala 17:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[MapS.scala 17:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[MapS.scala 17:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[MapS.scala 17:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[MapS.scala 17:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[MapS.scala 17:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[MapS.scala 21:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[MapS.scala 21:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[MapS.scala 21:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[MapS.scala 21:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[MapS.scala 21:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[MapS.scala 21:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[MapS.scala 21:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[MapS.scala 21:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[MapS.scala 21:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[MapS.scala 21:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[MapS.scala 21:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[MapS.scala 21:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[MapS.scala 21:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[MapS.scala 21:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[MapS.scala 21:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[MapS.scala 21:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[MapS.scala 21:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[MapS.scala 21:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[MapS.scala 21:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[MapS.scala 21:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[MapS.scala 21:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0_0 = I_0_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_1 = I_0_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_2 = I_0_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_0 = I_0_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_1 = I_0_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_2 = I_0_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_0 = I_0_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_1 = I_0_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_2 = I_0_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0_0 = I_1_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_1 = I_1_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_2 = I_1_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_0 = I_1_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_1 = I_1_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_2 = I_1_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_0 = I_1_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_1 = I_1_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_2 = I_1_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0_0 = I_2_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_1 = I_2_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_2 = I_2_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_0 = I_2_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_1 = I_2_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_2 = I_2_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_0 = I_2_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_1 = I_2_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_2 = I_2_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0_0 = I_3_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_1 = I_3_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_2 = I_3_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_0 = I_3_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_1 = I_3_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_2 = I_3_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_0 = I_3_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_1 = I_3_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_2 = I_3_0_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_7(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0_0,
  input  [15:0] I_0_0_0_1,
  input  [15:0] I_0_0_0_2,
  input  [15:0] I_0_0_1_0,
  input  [15:0] I_0_0_1_1,
  input  [15:0] I_0_0_1_2,
  input  [15:0] I_0_0_2_0,
  input  [15:0] I_0_0_2_1,
  input  [15:0] I_0_0_2_2,
  input  [15:0] I_1_0_0_0,
  input  [15:0] I_1_0_0_1,
  input  [15:0] I_1_0_0_2,
  input  [15:0] I_1_0_1_0,
  input  [15:0] I_1_0_1_1,
  input  [15:0] I_1_0_1_2,
  input  [15:0] I_1_0_2_0,
  input  [15:0] I_1_0_2_1,
  input  [15:0] I_1_0_2_2,
  input  [15:0] I_2_0_0_0,
  input  [15:0] I_2_0_0_1,
  input  [15:0] I_2_0_0_2,
  input  [15:0] I_2_0_1_0,
  input  [15:0] I_2_0_1_1,
  input  [15:0] I_2_0_1_2,
  input  [15:0] I_2_0_2_0,
  input  [15:0] I_2_0_2_1,
  input  [15:0] I_2_0_2_2,
  input  [15:0] I_3_0_0_0,
  input  [15:0] I_3_0_0_1,
  input  [15:0] I_3_0_0_2,
  input  [15:0] I_3_0_1_0,
  input  [15:0] I_3_0_1_1,
  input  [15:0] I_3_0_1_2,
  input  [15:0] I_3_0_2_0,
  input  [15:0] I_3_0_2_1,
  input  [15:0] I_3_0_2_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_0_2_0,
  output [15:0] O_0_2_1,
  output [15:0] O_0_2_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_1_2_0,
  output [15:0] O_1_2_1,
  output [15:0] O_1_2_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_2_2_0,
  output [15:0] O_2_2_1,
  output [15:0] O_2_2_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_3_2_0,
  output [15:0] O_3_2_1,
  output [15:0] O_3_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_2_2; // @[MapT.scala 8:20]
  MapS_3 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0_0(op_I_0_0_0_0),
    .I_0_0_0_1(op_I_0_0_0_1),
    .I_0_0_0_2(op_I_0_0_0_2),
    .I_0_0_1_0(op_I_0_0_1_0),
    .I_0_0_1_1(op_I_0_0_1_1),
    .I_0_0_1_2(op_I_0_0_1_2),
    .I_0_0_2_0(op_I_0_0_2_0),
    .I_0_0_2_1(op_I_0_0_2_1),
    .I_0_0_2_2(op_I_0_0_2_2),
    .I_1_0_0_0(op_I_1_0_0_0),
    .I_1_0_0_1(op_I_1_0_0_1),
    .I_1_0_0_2(op_I_1_0_0_2),
    .I_1_0_1_0(op_I_1_0_1_0),
    .I_1_0_1_1(op_I_1_0_1_1),
    .I_1_0_1_2(op_I_1_0_1_2),
    .I_1_0_2_0(op_I_1_0_2_0),
    .I_1_0_2_1(op_I_1_0_2_1),
    .I_1_0_2_2(op_I_1_0_2_2),
    .I_2_0_0_0(op_I_2_0_0_0),
    .I_2_0_0_1(op_I_2_0_0_1),
    .I_2_0_0_2(op_I_2_0_0_2),
    .I_2_0_1_0(op_I_2_0_1_0),
    .I_2_0_1_1(op_I_2_0_1_1),
    .I_2_0_1_2(op_I_2_0_1_2),
    .I_2_0_2_0(op_I_2_0_2_0),
    .I_2_0_2_1(op_I_2_0_2_1),
    .I_2_0_2_2(op_I_2_0_2_2),
    .I_3_0_0_0(op_I_3_0_0_0),
    .I_3_0_0_1(op_I_3_0_0_1),
    .I_3_0_0_2(op_I_3_0_0_2),
    .I_3_0_1_0(op_I_3_0_1_0),
    .I_3_0_1_1(op_I_3_0_1_1),
    .I_3_0_1_2(op_I_3_0_1_2),
    .I_3_0_2_0(op_I_3_0_2_0),
    .I_3_0_2_1(op_I_3_0_2_1),
    .I_3_0_2_2(op_I_3_0_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_2_2_0(op_O_2_2_0),
    .O_2_2_1(op_O_2_2_1),
    .O_2_2_2(op_O_2_2_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_3_2_0(op_O_3_2_0),
    .O_3_2_1(op_O_3_2_1),
    .O_3_2_2(op_O_3_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_0_1_0 = op_O_0_1_0; // @[MapT.scala 15:7]
  assign O_0_1_1 = op_O_0_1_1; // @[MapT.scala 15:7]
  assign O_0_1_2 = op_O_0_1_2; // @[MapT.scala 15:7]
  assign O_0_2_0 = op_O_0_2_0; // @[MapT.scala 15:7]
  assign O_0_2_1 = op_O_0_2_1; // @[MapT.scala 15:7]
  assign O_0_2_2 = op_O_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_1_1_0 = op_O_1_1_0; // @[MapT.scala 15:7]
  assign O_1_1_1 = op_O_1_1_1; // @[MapT.scala 15:7]
  assign O_1_1_2 = op_O_1_1_2; // @[MapT.scala 15:7]
  assign O_1_2_0 = op_O_1_2_0; // @[MapT.scala 15:7]
  assign O_1_2_1 = op_O_1_2_1; // @[MapT.scala 15:7]
  assign O_1_2_2 = op_O_1_2_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_2_1_0 = op_O_2_1_0; // @[MapT.scala 15:7]
  assign O_2_1_1 = op_O_2_1_1; // @[MapT.scala 15:7]
  assign O_2_1_2 = op_O_2_1_2; // @[MapT.scala 15:7]
  assign O_2_2_0 = op_O_2_2_0; // @[MapT.scala 15:7]
  assign O_2_2_1 = op_O_2_2_1; // @[MapT.scala 15:7]
  assign O_2_2_2 = op_O_2_2_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign O_3_1_0 = op_O_3_1_0; // @[MapT.scala 15:7]
  assign O_3_1_1 = op_O_3_1_1; // @[MapT.scala 15:7]
  assign O_3_1_2 = op_O_3_1_2; // @[MapT.scala 15:7]
  assign O_3_2_0 = op_O_3_2_0; // @[MapT.scala 15:7]
  assign O_3_2_1 = op_O_3_2_1; // @[MapT.scala 15:7]
  assign O_3_2_2 = op_O_3_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0_0 = I_0_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_0_1 = I_0_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_0_2 = I_0_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_0_1_0 = I_0_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1_1 = I_0_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_0_1_2 = I_0_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_0_2_0 = I_0_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_0_2_1 = I_0_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2_2 = I_0_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0_0 = I_1_0_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_0_1 = I_1_0_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0_2 = I_1_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_1_0 = I_1_0_1_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1_1 = I_1_0_1_1; // @[MapT.scala 14:10]
  assign op_I_1_0_1_2 = I_1_0_1_2; // @[MapT.scala 14:10]
  assign op_I_1_0_2_0 = I_1_0_2_0; // @[MapT.scala 14:10]
  assign op_I_1_0_2_1 = I_1_0_2_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2_2 = I_1_0_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0_0 = I_2_0_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_0_1 = I_2_0_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0_2 = I_2_0_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_1_0 = I_2_0_1_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1_1 = I_2_0_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0_1_2 = I_2_0_1_2; // @[MapT.scala 14:10]
  assign op_I_2_0_2_0 = I_2_0_2_0; // @[MapT.scala 14:10]
  assign op_I_2_0_2_1 = I_2_0_2_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2_2 = I_2_0_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0_0 = I_3_0_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_0_1 = I_3_0_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0_2 = I_3_0_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_1_0 = I_3_0_1_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1_1 = I_3_0_1_1; // @[MapT.scala 14:10]
  assign op_I_3_0_1_2 = I_3_0_1_2; // @[MapT.scala 14:10]
  assign op_I_3_0_2_0 = I_3_0_2_0; // @[MapT.scala 14:10]
  assign op_I_3_0_2_1 = I_3_0_2_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2_2 = I_3_0_2_2; // @[MapT.scala 14:10]
endmodule
module InitialDelayCounter(
  input   clock,
  input   reset,
  output  valid_down
);
  reg  value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire  _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 1'h1; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 1'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 1'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module AtomTuple(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0,
  input  [15:0] I1,
  output [15:0] O_t0b,
  output [15:0] O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Map2S_8(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I0_2,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  output [15:0] O_0_t0b,
  output [15:0] O_0_t1b,
  output [15:0] O_1_t0b,
  output [15:0] O_1_t1b,
  output [15:0] O_2_t0b,
  output [15:0] O_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  AtomTuple other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  AtomTuple other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_t0b(other_ops_1_O_t0b),
    .O_t1b(other_ops_1_O_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign O_2_t0b = other_ops_1_O_t0b; // @[Map2S.scala 24:12]
  assign O_2_t1b = other_ops_1_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
endmodule
module Map2S_9(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_0_2,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_1_2,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_2_2,
  output [15:0] O_0_0_t0b,
  output [15:0] O_0_0_t1b,
  output [15:0] O_0_1_t0b,
  output [15:0] O_0_1_t1b,
  output [15:0] O_0_2_t0b,
  output [15:0] O_0_2_t1b,
  output [15:0] O_1_0_t0b,
  output [15:0] O_1_0_t1b,
  output [15:0] O_1_1_t0b,
  output [15:0] O_1_1_t1b,
  output [15:0] O_1_2_t0b,
  output [15:0] O_1_2_t1b,
  output [15:0] O_2_0_t0b,
  output [15:0] O_2_0_t1b,
  output [15:0] O_2_1_t0b,
  output [15:0] O_2_1_t1b,
  output [15:0] O_2_2_t0b,
  output [15:0] O_2_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_t0b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_t1b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2_t0b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_t1b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_t1b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_t1b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_t1b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  Map2S_8 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b),
    .O_1_t0b(fst_op_O_1_t0b),
    .O_1_t1b(fst_op_O_1_t1b),
    .O_2_t0b(fst_op_O_2_t0b),
    .O_2_t1b(fst_op_O_2_t1b)
  );
  Map2S_8 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_t0b(other_ops_0_O_0_t0b),
    .O_0_t1b(other_ops_0_O_0_t1b),
    .O_1_t0b(other_ops_0_O_1_t0b),
    .O_1_t1b(other_ops_0_O_1_t1b),
    .O_2_t0b(other_ops_0_O_2_t0b),
    .O_2_t1b(other_ops_0_O_2_t1b)
  );
  Map2S_8 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_t0b(other_ops_1_O_0_t0b),
    .O_0_t1b(other_ops_1_O_0_t1b),
    .O_1_t0b(other_ops_1_O_1_t0b),
    .O_1_t1b(other_ops_1_O_1_t1b),
    .O_2_t0b(other_ops_1_O_2_t0b),
    .O_2_t1b(other_ops_1_O_2_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign O_0_1_t0b = fst_op_O_1_t0b; // @[Map2S.scala 19:8]
  assign O_0_1_t1b = fst_op_O_1_t1b; // @[Map2S.scala 19:8]
  assign O_0_2_t0b = fst_op_O_2_t0b; // @[Map2S.scala 19:8]
  assign O_0_2_t1b = fst_op_O_2_t1b; // @[Map2S.scala 19:8]
  assign O_1_0_t0b = other_ops_0_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_1_0_t1b = other_ops_0_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_1_1_t0b = other_ops_0_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_1_1_t1b = other_ops_0_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_1_2_t0b = other_ops_0_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_1_2_t1b = other_ops_0_O_2_t1b; // @[Map2S.scala 24:12]
  assign O_2_0_t0b = other_ops_1_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_2_0_t1b = other_ops_1_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_2_1_t0b = other_ops_1_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_2_1_t1b = other_ops_1_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_2_2_t0b = other_ops_1_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_2_2_t1b = other_ops_1_O_2_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = 16'h1; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = 16'h2; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = 16'h1; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = 16'h2; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = 16'h4; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = 16'h2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = 16'h1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = 16'h2; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = 16'h1; // @[Map2S.scala 23:43]
endmodule
module Mul(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_t0b,
  input  [15:0] I_t1b,
  output [15:0] O
);
  wire [15:0] BlackBoxMulUInt16_I0; // @[Arithmetic.scala 180:27]
  wire [15:0] BlackBoxMulUInt16_I1; // @[Arithmetic.scala 180:27]
  wire [31:0] BlackBoxMulUInt16_O; // @[Arithmetic.scala 180:27]
  wire  BlackBoxMulUInt16_clock; // @[Arithmetic.scala 180:27]
  reg  _T_1; // @[Arithmetic.scala 217:42]
  reg [31:0] _RAND_0;
  reg  _T_2; // @[Arithmetic.scala 217:34]
  reg [31:0] _RAND_1;
  reg  _T_3; // @[Arithmetic.scala 217:26]
  reg [31:0] _RAND_2;
  BlackBoxMulUInt16 BlackBoxMulUInt16 ( // @[Arithmetic.scala 180:27]
    .I0(BlackBoxMulUInt16_I0),
    .I1(BlackBoxMulUInt16_I1),
    .O(BlackBoxMulUInt16_O),
    .clock(BlackBoxMulUInt16_clock)
  );
  assign valid_down = _T_3; // @[Arithmetic.scala 217:16]
  assign O = BlackBoxMulUInt16_O[15:0]; // @[Arithmetic.scala 183:7]
  assign BlackBoxMulUInt16_I0 = I_t0b; // @[Arithmetic.scala 181:21]
  assign BlackBoxMulUInt16_I1 = I_t1b; // @[Arithmetic.scala 182:21]
  assign BlackBoxMulUInt16_clock = clock; // @[Arithmetic.scala 184:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_3 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
    if (reset) begin
      _T_2 <= 1'h0;
    end else begin
      _T_2 <= _T_1;
    end
    if (reset) begin
      _T_3 <= 1'h0;
    end else begin
      _T_3 <= _T_2;
    end
  end
endmodule
module MapS_4(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_t0b,
  input  [15:0] I_0_t1b,
  input  [15:0] I_1_t0b,
  input  [15:0] I_1_t1b,
  input  [15:0] I_2_t0b,
  input  [15:0] I_2_t1b,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  Mul fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  Mul other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t0b(other_ops_0_I_t0b),
    .I_t1b(other_ops_0_I_t1b),
    .O(other_ops_0_O)
  );
  Mul other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_t0b(other_ops_1_I_t0b),
    .I_t1b(other_ops_1_I_t1b),
    .O(other_ops_1_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t0b = I_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_t1b = I_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_t0b = I_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_t1b = I_2_t1b; // @[MapS.scala 20:41]
endmodule
module MapS_5(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_t0b,
  input  [15:0] I_0_0_t1b,
  input  [15:0] I_0_1_t0b,
  input  [15:0] I_0_1_t1b,
  input  [15:0] I_0_2_t0b,
  input  [15:0] I_0_2_t1b,
  input  [15:0] I_1_0_t0b,
  input  [15:0] I_1_0_t1b,
  input  [15:0] I_1_1_t0b,
  input  [15:0] I_1_1_t1b,
  input  [15:0] I_1_2_t0b,
  input  [15:0] I_1_2_t1b,
  input  [15:0] I_2_0_t0b,
  input  [15:0] I_2_0_t1b,
  input  [15:0] I_2_1_t0b,
  input  [15:0] I_2_1_t1b,
  input  [15:0] I_2_2_t0b,
  input  [15:0] I_2_2_t1b,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_t0b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2_t0b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  MapS_4 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .I_1_t0b(fst_op_I_1_t0b),
    .I_1_t1b(fst_op_I_1_t1b),
    .I_2_t0b(fst_op_I_2_t0b),
    .I_2_t1b(fst_op_I_2_t1b),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  MapS_4 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_t0b(other_ops_0_I_0_t0b),
    .I_0_t1b(other_ops_0_I_0_t1b),
    .I_1_t0b(other_ops_0_I_1_t0b),
    .I_1_t1b(other_ops_0_I_1_t1b),
    .I_2_t0b(other_ops_0_I_2_t0b),
    .I_2_t1b(other_ops_0_I_2_t1b),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  MapS_4 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_t0b(other_ops_1_I_0_t0b),
    .I_0_t1b(other_ops_1_I_0_t1b),
    .I_1_t0b(other_ops_1_I_1_t0b),
    .I_1_t1b(other_ops_1_I_1_t1b),
    .I_2_t0b(other_ops_1_I_2_t0b),
    .I_2_t1b(other_ops_1_I_2_t1b),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t0b = I_0_1_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t1b = I_0_1_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t0b = I_0_2_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t1b = I_0_2_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_t0b = I_1_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_t1b = I_1_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t0b = I_1_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t1b = I_1_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t0b = I_1_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t1b = I_1_2_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_t0b = I_2_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_t1b = I_2_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t0b = I_2_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t1b = I_2_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t0b = I_2_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t1b = I_2_2_t1b; // @[MapS.scala 20:41]
endmodule
module AddNoValid(
  input  [15:0] I_t0b,
  input  [15:0] I_t1b,
  output [15:0] O
);
  assign O = I_t0b + I_t1b; // @[Arithmetic.scala 122:7]
endmodule
module ReduceS(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  output [15:0] O_0
);
  wire [15:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_1_O; // @[ReduceS.scala 20:43]
  reg [15:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [15:0] _T_1; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [15:0] _T_2; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [15:0] _T_3; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_5;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  AddNoValid AddNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_1_I_t0b),
    .I_t1b(AddNoValid_1_I_t1b),
    .O(AddNoValid_1_O)
  );
  assign valid_down = _T_5; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = _T_3; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = AddNoValid_1_O; // @[ReduceS.scala 36:18]
  assign AddNoValid_1_I_t0b = _T_2; // @[ReduceS.scala 43:18]
  assign AddNoValid_1_I_t1b = _T_1; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    _T_1 <= I_0;
    _T_2 <= I_1;
    _T_3 <= I_2;
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= valid_up;
    end
    _T_5 <= _T_4;
  end
endmodule
module MapS_6(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  output [15:0] O_0_0,
  output [15:0] O_1_0,
  output [15:0] O_2_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  ReduceS fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .O_0(fst_op_O_0)
  );
  ReduceS other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0(other_ops_0_I_0),
    .I_1(other_ops_0_I_1),
    .I_2(other_ops_0_I_2),
    .O_0(other_ops_0_O_0)
  );
  ReduceS other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0(other_ops_1_I_0),
    .I_1(other_ops_1_I_1),
    .I_2(other_ops_1_I_2),
    .O_0(other_ops_1_O_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0 = I_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1 = I_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2 = I_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0 = I_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1 = I_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2 = I_2_2; // @[MapS.scala 20:41]
endmodule
module MapSNoValid(
  input  [15:0] I_0_t0b,
  input  [15:0] I_0_t1b,
  output [15:0] O_0
);
  wire [15:0] fst_op_I_t0b; // @[MapS.scala 28:22]
  wire [15:0] fst_op_I_t1b; // @[MapS.scala 28:22]
  wire [15:0] fst_op_O; // @[MapS.scala 28:22]
  AddNoValid fst_op ( // @[MapS.scala 28:22]
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign O_0 = fst_op_O; // @[MapS.scala 35:8]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 34:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 34:12]
endmodule
module ReduceS_1(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_1_0,
  input  [15:0] I_2_0,
  output [15:0] O_0_0
);
  wire [15:0] MapSNoValid_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_O_0; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_1_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_1_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_1_O_0; // @[ReduceS.scala 20:43]
  reg [15:0] _T_0; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [15:0] _T_1_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [15:0] _T_2_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [15:0] _T_3_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_5;
  MapSNoValid MapSNoValid ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_I_0_t0b),
    .I_0_t1b(MapSNoValid_I_0_t1b),
    .O_0(MapSNoValid_O_0)
  );
  MapSNoValid MapSNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_1_I_0_t0b),
    .I_0_t1b(MapSNoValid_1_I_0_t1b),
    .O_0(MapSNoValid_1_O_0)
  );
  assign valid_down = _T_5; // @[ReduceS.scala 47:14]
  assign O_0_0 = _T_0; // @[ReduceS.scala 27:14]
  assign MapSNoValid_I_0_t0b = _T_2_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_I_0_t1b = MapSNoValid_1_O_0; // @[ReduceS.scala 36:18]
  assign MapSNoValid_1_I_0_t0b = _T_1_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_1_I_0_t1b = _T_3_0; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1_0 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2_0 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3_0 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= MapSNoValid_O_0;
    _T_1_0 <= I_0_0;
    _T_2_0 <= I_1_0;
    _T_3_0 <= I_2_0;
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= valid_up;
    end
    _T_5 <= _T_4;
  end
endmodule
module InitialDelayCounter_1(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [3:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [3:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 4'h8; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 4'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 4'h8; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 4'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module AtomTuple_1(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0,
  input  [7:0]  I1,
  output [15:0] O_t0b,
  output [7:0]  O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Map2S_10(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [7:0]  I1_0,
  output [15:0] O_0_t0b,
  output [7:0]  O_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  AtomTuple_1 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_11(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [7:0]  I1_0_0,
  output [15:0] O_0_0_t0b,
  output [7:0]  O_0_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  Map2S_10 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I1_0(fst_op_I1_0),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
endmodule
module Div(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_t0b,
  input  [7:0]  I_t1b,
  output [15:0] O
);
  wire [15:0] BlackBoxMulUInt16_I0; // @[Arithmetic.scala 349:27]
  wire [15:0] BlackBoxMulUInt16_I1; // @[Arithmetic.scala 349:27]
  wire [31:0] BlackBoxMulUInt16_O; // @[Arithmetic.scala 349:27]
  wire  BlackBoxMulUInt16_clock; // @[Arithmetic.scala 349:27]
  wire [8:0] _T_1; // @[Cat.scala 29:58]
  reg  _T_3; // @[Arithmetic.scala 370:42]
  reg [31:0] _RAND_0;
  reg  _T_4; // @[Arithmetic.scala 370:34]
  reg [31:0] _RAND_1;
  reg  _T_5; // @[Arithmetic.scala 370:26]
  reg [31:0] _RAND_2;
  BlackBoxMulUInt16 BlackBoxMulUInt16 ( // @[Arithmetic.scala 349:27]
    .I0(BlackBoxMulUInt16_I0),
    .I1(BlackBoxMulUInt16_I1),
    .O(BlackBoxMulUInt16_O),
    .clock(BlackBoxMulUInt16_clock)
  );
  assign _T_1 = {1'h0,I_t1b}; // @[Cat.scala 29:58]
  assign valid_down = _T_5; // @[Arithmetic.scala 370:16]
  assign O = BlackBoxMulUInt16_O[22:7]; // @[Arithmetic.scala 352:7]
  assign BlackBoxMulUInt16_I0 = I_t0b; // @[Arithmetic.scala 350:21]
  assign BlackBoxMulUInt16_I1 = {{7'd0}, _T_1}; // @[Arithmetic.scala 351:21]
  assign BlackBoxMulUInt16_clock = clock; // @[Arithmetic.scala 353:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_3 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_4 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_5 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_3 <= 1'h0;
    end else begin
      _T_3 <= valid_up;
    end
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= _T_3;
    end
    if (reset) begin
      _T_5 <= 1'h0;
    end else begin
      _T_5 <= _T_4;
    end
  end
endmodule
module MapS_7(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_t0b,
  input  [7:0]  I_0_t1b,
  output [15:0] O_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O; // @[MapS.scala 9:22]
  Div fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
endmodule
module MapS_8(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_t0b,
  input  [7:0]  I_0_0_t1b,
  output [15:0] O_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0; // @[MapS.scala 9:22]
  MapS_7 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
endmodule
module Module_0(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  output [15:0] O_0_0
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n110_valid_up; // @[Top.scala 18:22]
  wire  n110_valid_down; // @[Top.scala 18:22]
  wire [15:0] n110_I0_0_0; // @[Top.scala 18:22]
  wire [15:0] n110_I0_0_1; // @[Top.scala 18:22]
  wire [15:0] n110_I0_0_2; // @[Top.scala 18:22]
  wire [15:0] n110_I0_1_0; // @[Top.scala 18:22]
  wire [15:0] n110_I0_1_1; // @[Top.scala 18:22]
  wire [15:0] n110_I0_1_2; // @[Top.scala 18:22]
  wire [15:0] n110_I0_2_0; // @[Top.scala 18:22]
  wire [15:0] n110_I0_2_1; // @[Top.scala 18:22]
  wire [15:0] n110_I0_2_2; // @[Top.scala 18:22]
  wire [15:0] n110_O_0_0_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_0_0_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_0_1_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_0_1_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_0_2_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_0_2_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_1_0_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_1_0_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_1_1_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_1_1_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_1_2_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_1_2_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_2_0_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_2_0_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_2_1_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_2_1_t1b; // @[Top.scala 18:22]
  wire [15:0] n110_O_2_2_t0b; // @[Top.scala 18:22]
  wire [15:0] n110_O_2_2_t1b; // @[Top.scala 18:22]
  wire  n121_clock; // @[Top.scala 22:22]
  wire  n121_reset; // @[Top.scala 22:22]
  wire  n121_valid_up; // @[Top.scala 22:22]
  wire  n121_valid_down; // @[Top.scala 22:22]
  wire [15:0] n121_I_0_0_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_0_0_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_0_1_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_0_1_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_0_2_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_0_2_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_1_0_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_1_0_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_1_1_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_1_1_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_1_2_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_1_2_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_2_0_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_2_0_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_2_1_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_2_1_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_I_2_2_t0b; // @[Top.scala 22:22]
  wire [15:0] n121_I_2_2_t1b; // @[Top.scala 22:22]
  wire [15:0] n121_O_0_0; // @[Top.scala 22:22]
  wire [15:0] n121_O_0_1; // @[Top.scala 22:22]
  wire [15:0] n121_O_0_2; // @[Top.scala 22:22]
  wire [15:0] n121_O_1_0; // @[Top.scala 22:22]
  wire [15:0] n121_O_1_1; // @[Top.scala 22:22]
  wire [15:0] n121_O_1_2; // @[Top.scala 22:22]
  wire [15:0] n121_O_2_0; // @[Top.scala 22:22]
  wire [15:0] n121_O_2_1; // @[Top.scala 22:22]
  wire [15:0] n121_O_2_2; // @[Top.scala 22:22]
  wire  n126_clock; // @[Top.scala 25:22]
  wire  n126_reset; // @[Top.scala 25:22]
  wire  n126_valid_up; // @[Top.scala 25:22]
  wire  n126_valid_down; // @[Top.scala 25:22]
  wire [15:0] n126_I_0_0; // @[Top.scala 25:22]
  wire [15:0] n126_I_0_1; // @[Top.scala 25:22]
  wire [15:0] n126_I_0_2; // @[Top.scala 25:22]
  wire [15:0] n126_I_1_0; // @[Top.scala 25:22]
  wire [15:0] n126_I_1_1; // @[Top.scala 25:22]
  wire [15:0] n126_I_1_2; // @[Top.scala 25:22]
  wire [15:0] n126_I_2_0; // @[Top.scala 25:22]
  wire [15:0] n126_I_2_1; // @[Top.scala 25:22]
  wire [15:0] n126_I_2_2; // @[Top.scala 25:22]
  wire [15:0] n126_O_0_0; // @[Top.scala 25:22]
  wire [15:0] n126_O_1_0; // @[Top.scala 25:22]
  wire [15:0] n126_O_2_0; // @[Top.scala 25:22]
  wire  n131_clock; // @[Top.scala 28:22]
  wire  n131_reset; // @[Top.scala 28:22]
  wire  n131_valid_up; // @[Top.scala 28:22]
  wire  n131_valid_down; // @[Top.scala 28:22]
  wire [15:0] n131_I_0_0; // @[Top.scala 28:22]
  wire [15:0] n131_I_1_0; // @[Top.scala 28:22]
  wire [15:0] n131_I_2_0; // @[Top.scala 28:22]
  wire [15:0] n131_O_0_0; // @[Top.scala 28:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n134_valid_up; // @[Top.scala 32:22]
  wire  n134_valid_down; // @[Top.scala 32:22]
  wire [15:0] n134_I0_0_0; // @[Top.scala 32:22]
  wire [7:0] n134_I1_0_0; // @[Top.scala 32:22]
  wire [15:0] n134_O_0_0_t0b; // @[Top.scala 32:22]
  wire [7:0] n134_O_0_0_t1b; // @[Top.scala 32:22]
  wire  n145_clock; // @[Top.scala 36:22]
  wire  n145_reset; // @[Top.scala 36:22]
  wire  n145_valid_up; // @[Top.scala 36:22]
  wire  n145_valid_down; // @[Top.scala 36:22]
  wire [15:0] n145_I_0_0_t0b; // @[Top.scala 36:22]
  wire [7:0] n145_I_0_0_t1b; // @[Top.scala 36:22]
  wire [15:0] n145_O_0_0; // @[Top.scala 36:22]
  InitialDelayCounter InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  Map2S_9 n110 ( // @[Top.scala 18:22]
    .valid_up(n110_valid_up),
    .valid_down(n110_valid_down),
    .I0_0_0(n110_I0_0_0),
    .I0_0_1(n110_I0_0_1),
    .I0_0_2(n110_I0_0_2),
    .I0_1_0(n110_I0_1_0),
    .I0_1_1(n110_I0_1_1),
    .I0_1_2(n110_I0_1_2),
    .I0_2_0(n110_I0_2_0),
    .I0_2_1(n110_I0_2_1),
    .I0_2_2(n110_I0_2_2),
    .O_0_0_t0b(n110_O_0_0_t0b),
    .O_0_0_t1b(n110_O_0_0_t1b),
    .O_0_1_t0b(n110_O_0_1_t0b),
    .O_0_1_t1b(n110_O_0_1_t1b),
    .O_0_2_t0b(n110_O_0_2_t0b),
    .O_0_2_t1b(n110_O_0_2_t1b),
    .O_1_0_t0b(n110_O_1_0_t0b),
    .O_1_0_t1b(n110_O_1_0_t1b),
    .O_1_1_t0b(n110_O_1_1_t0b),
    .O_1_1_t1b(n110_O_1_1_t1b),
    .O_1_2_t0b(n110_O_1_2_t0b),
    .O_1_2_t1b(n110_O_1_2_t1b),
    .O_2_0_t0b(n110_O_2_0_t0b),
    .O_2_0_t1b(n110_O_2_0_t1b),
    .O_2_1_t0b(n110_O_2_1_t0b),
    .O_2_1_t1b(n110_O_2_1_t1b),
    .O_2_2_t0b(n110_O_2_2_t0b),
    .O_2_2_t1b(n110_O_2_2_t1b)
  );
  MapS_5 n121 ( // @[Top.scala 22:22]
    .clock(n121_clock),
    .reset(n121_reset),
    .valid_up(n121_valid_up),
    .valid_down(n121_valid_down),
    .I_0_0_t0b(n121_I_0_0_t0b),
    .I_0_0_t1b(n121_I_0_0_t1b),
    .I_0_1_t0b(n121_I_0_1_t0b),
    .I_0_1_t1b(n121_I_0_1_t1b),
    .I_0_2_t0b(n121_I_0_2_t0b),
    .I_0_2_t1b(n121_I_0_2_t1b),
    .I_1_0_t0b(n121_I_1_0_t0b),
    .I_1_0_t1b(n121_I_1_0_t1b),
    .I_1_1_t0b(n121_I_1_1_t0b),
    .I_1_1_t1b(n121_I_1_1_t1b),
    .I_1_2_t0b(n121_I_1_2_t0b),
    .I_1_2_t1b(n121_I_1_2_t1b),
    .I_2_0_t0b(n121_I_2_0_t0b),
    .I_2_0_t1b(n121_I_2_0_t1b),
    .I_2_1_t0b(n121_I_2_1_t0b),
    .I_2_1_t1b(n121_I_2_1_t1b),
    .I_2_2_t0b(n121_I_2_2_t0b),
    .I_2_2_t1b(n121_I_2_2_t1b),
    .O_0_0(n121_O_0_0),
    .O_0_1(n121_O_0_1),
    .O_0_2(n121_O_0_2),
    .O_1_0(n121_O_1_0),
    .O_1_1(n121_O_1_1),
    .O_1_2(n121_O_1_2),
    .O_2_0(n121_O_2_0),
    .O_2_1(n121_O_2_1),
    .O_2_2(n121_O_2_2)
  );
  MapS_6 n126 ( // @[Top.scala 25:22]
    .clock(n126_clock),
    .reset(n126_reset),
    .valid_up(n126_valid_up),
    .valid_down(n126_valid_down),
    .I_0_0(n126_I_0_0),
    .I_0_1(n126_I_0_1),
    .I_0_2(n126_I_0_2),
    .I_1_0(n126_I_1_0),
    .I_1_1(n126_I_1_1),
    .I_1_2(n126_I_1_2),
    .I_2_0(n126_I_2_0),
    .I_2_1(n126_I_2_1),
    .I_2_2(n126_I_2_2),
    .O_0_0(n126_O_0_0),
    .O_1_0(n126_O_1_0),
    .O_2_0(n126_O_2_0)
  );
  ReduceS_1 n131 ( // @[Top.scala 28:22]
    .clock(n131_clock),
    .reset(n131_reset),
    .valid_up(n131_valid_up),
    .valid_down(n131_valid_down),
    .I_0_0(n131_I_0_0),
    .I_1_0(n131_I_1_0),
    .I_2_0(n131_I_2_0),
    .O_0_0(n131_O_0_0)
  );
  InitialDelayCounter_1 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  Map2S_11 n134 ( // @[Top.scala 32:22]
    .valid_up(n134_valid_up),
    .valid_down(n134_valid_down),
    .I0_0_0(n134_I0_0_0),
    .I1_0_0(n134_I1_0_0),
    .O_0_0_t0b(n134_O_0_0_t0b),
    .O_0_0_t1b(n134_O_0_0_t1b)
  );
  MapS_8 n145 ( // @[Top.scala 36:22]
    .clock(n145_clock),
    .reset(n145_reset),
    .valid_up(n145_valid_up),
    .valid_down(n145_valid_down),
    .I_0_0_t0b(n145_I_0_0_t0b),
    .I_0_0_t1b(n145_I_0_0_t1b),
    .O_0_0(n145_O_0_0)
  );
  assign valid_down = n145_valid_down; // @[Top.scala 40:16]
  assign O_0_0 = n145_O_0_0; // @[Top.scala 39:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n110_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 21:19]
  assign n110_I0_0_0 = I_0_0; // @[Top.scala 19:13]
  assign n110_I0_0_1 = I_0_1; // @[Top.scala 19:13]
  assign n110_I0_0_2 = I_0_2; // @[Top.scala 19:13]
  assign n110_I0_1_0 = I_1_0; // @[Top.scala 19:13]
  assign n110_I0_1_1 = I_1_1; // @[Top.scala 19:13]
  assign n110_I0_1_2 = I_1_2; // @[Top.scala 19:13]
  assign n110_I0_2_0 = I_2_0; // @[Top.scala 19:13]
  assign n110_I0_2_1 = I_2_1; // @[Top.scala 19:13]
  assign n110_I0_2_2 = I_2_2; // @[Top.scala 19:13]
  assign n121_clock = clock;
  assign n121_reset = reset;
  assign n121_valid_up = n110_valid_down; // @[Top.scala 24:19]
  assign n121_I_0_0_t0b = n110_O_0_0_t0b; // @[Top.scala 23:12]
  assign n121_I_0_0_t1b = n110_O_0_0_t1b; // @[Top.scala 23:12]
  assign n121_I_0_1_t0b = n110_O_0_1_t0b; // @[Top.scala 23:12]
  assign n121_I_0_1_t1b = n110_O_0_1_t1b; // @[Top.scala 23:12]
  assign n121_I_0_2_t0b = n110_O_0_2_t0b; // @[Top.scala 23:12]
  assign n121_I_0_2_t1b = n110_O_0_2_t1b; // @[Top.scala 23:12]
  assign n121_I_1_0_t0b = n110_O_1_0_t0b; // @[Top.scala 23:12]
  assign n121_I_1_0_t1b = n110_O_1_0_t1b; // @[Top.scala 23:12]
  assign n121_I_1_1_t0b = n110_O_1_1_t0b; // @[Top.scala 23:12]
  assign n121_I_1_1_t1b = n110_O_1_1_t1b; // @[Top.scala 23:12]
  assign n121_I_1_2_t0b = n110_O_1_2_t0b; // @[Top.scala 23:12]
  assign n121_I_1_2_t1b = n110_O_1_2_t1b; // @[Top.scala 23:12]
  assign n121_I_2_0_t0b = n110_O_2_0_t0b; // @[Top.scala 23:12]
  assign n121_I_2_0_t1b = n110_O_2_0_t1b; // @[Top.scala 23:12]
  assign n121_I_2_1_t0b = n110_O_2_1_t0b; // @[Top.scala 23:12]
  assign n121_I_2_1_t1b = n110_O_2_1_t1b; // @[Top.scala 23:12]
  assign n121_I_2_2_t0b = n110_O_2_2_t0b; // @[Top.scala 23:12]
  assign n121_I_2_2_t1b = n110_O_2_2_t1b; // @[Top.scala 23:12]
  assign n126_clock = clock;
  assign n126_reset = reset;
  assign n126_valid_up = n121_valid_down; // @[Top.scala 27:19]
  assign n126_I_0_0 = n121_O_0_0; // @[Top.scala 26:12]
  assign n126_I_0_1 = n121_O_0_1; // @[Top.scala 26:12]
  assign n126_I_0_2 = n121_O_0_2; // @[Top.scala 26:12]
  assign n126_I_1_0 = n121_O_1_0; // @[Top.scala 26:12]
  assign n126_I_1_1 = n121_O_1_1; // @[Top.scala 26:12]
  assign n126_I_1_2 = n121_O_1_2; // @[Top.scala 26:12]
  assign n126_I_2_0 = n121_O_2_0; // @[Top.scala 26:12]
  assign n126_I_2_1 = n121_O_2_1; // @[Top.scala 26:12]
  assign n126_I_2_2 = n121_O_2_2; // @[Top.scala 26:12]
  assign n131_clock = clock;
  assign n131_reset = reset;
  assign n131_valid_up = n126_valid_down; // @[Top.scala 30:19]
  assign n131_I_0_0 = n126_O_0_0; // @[Top.scala 29:12]
  assign n131_I_1_0 = n126_O_1_0; // @[Top.scala 29:12]
  assign n131_I_2_0 = n126_O_2_0; // @[Top.scala 29:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n134_valid_up = n131_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 35:19]
  assign n134_I0_0_0 = n131_O_0_0; // @[Top.scala 33:13]
  assign n134_I1_0_0 = 8'sh8; // @[Top.scala 34:13]
  assign n145_clock = clock;
  assign n145_reset = reset;
  assign n145_valid_up = n134_valid_down; // @[Top.scala 38:19]
  assign n145_I_0_0_t0b = n134_O_0_0_t0b; // @[Top.scala 37:12]
  assign n145_I_0_0_t1b = n134_O_0_0_t1b; // @[Top.scala 37:12]
endmodule
module MapS_9(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_0_1_2,
  input  [15:0] I_0_2_0,
  input  [15:0] I_0_2_1,
  input  [15:0] I_0_2_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_1_1_2,
  input  [15:0] I_1_2_0,
  input  [15:0] I_1_2_1,
  input  [15:0] I_1_2_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_2_1_2,
  input  [15:0] I_2_2_0,
  input  [15:0] I_2_2_1,
  input  [15:0] I_2_2_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  input  [15:0] I_3_1_2,
  input  [15:0] I_3_2_0,
  input  [15:0] I_3_2_1,
  input  [15:0] I_3_2_2,
  output [15:0] O_0_0_0,
  output [15:0] O_1_0_0,
  output [15:0] O_2_0_0,
  output [15:0] O_3_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_2_clock; // @[MapS.scala 10:86]
  wire  other_ops_2_reset; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  Module_0 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .I_1_0(fst_op_I_1_0),
    .I_1_1(fst_op_I_1_1),
    .I_1_2(fst_op_I_1_2),
    .I_2_0(fst_op_I_2_0),
    .I_2_1(fst_op_I_2_1),
    .I_2_2(fst_op_I_2_2),
    .O_0_0(fst_op_O_0_0)
  );
  Module_0 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .I_1_0(other_ops_0_I_1_0),
    .I_1_1(other_ops_0_I_1_1),
    .I_1_2(other_ops_0_I_1_2),
    .I_2_0(other_ops_0_I_2_0),
    .I_2_1(other_ops_0_I_2_1),
    .I_2_2(other_ops_0_I_2_2),
    .O_0_0(other_ops_0_O_0_0)
  );
  Module_0 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .I_1_0(other_ops_1_I_1_0),
    .I_1_1(other_ops_1_I_1_1),
    .I_1_2(other_ops_1_I_1_2),
    .I_2_0(other_ops_1_I_2_0),
    .I_2_1(other_ops_1_I_2_1),
    .I_2_2(other_ops_1_I_2_2),
    .O_0_0(other_ops_1_O_0_0)
  );
  Module_0 other_ops_2 ( // @[MapS.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .I_1_0(other_ops_2_I_1_0),
    .I_1_1(other_ops_2_I_1_1),
    .I_1_2(other_ops_2_I_1_2),
    .I_2_0(other_ops_2_I_2_0),
    .I_2_1(other_ops_2_I_2_1),
    .I_2_2(other_ops_2_I_2_2),
    .O_0_0(other_ops_2_O_0_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_1_0 = I_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_1_1 = I_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_1_2 = I_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_2_0 = I_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_2_1 = I_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_2_2 = I_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_0 = I_1_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_1 = I_1_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_2 = I_1_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_0 = I_1_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_1 = I_1_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_2 = I_1_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_0 = I_2_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_1 = I_2_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_2 = I_2_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_0 = I_2_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_1 = I_2_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_2 = I_2_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_2_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_0 = I_3_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_1 = I_3_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_2 = I_3_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_0 = I_3_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_1 = I_3_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_2 = I_3_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_8(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_0_1_2,
  input  [15:0] I_0_2_0,
  input  [15:0] I_0_2_1,
  input  [15:0] I_0_2_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_1_1_2,
  input  [15:0] I_1_2_0,
  input  [15:0] I_1_2_1,
  input  [15:0] I_1_2_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_2_1_2,
  input  [15:0] I_2_2_0,
  input  [15:0] I_2_2_1,
  input  [15:0] I_2_2_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  input  [15:0] I_3_1_2,
  input  [15:0] I_3_2_0,
  input  [15:0] I_3_2_1,
  input  [15:0] I_3_2_2,
  output [15:0] O_0_0_0,
  output [15:0] O_1_0_0,
  output [15:0] O_2_0_0,
  output [15:0] O_3_0_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[MapT.scala 8:20]
  MapS_9 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_1_0_0(op_O_1_0_0),
    .O_2_0_0(op_O_2_0_0),
    .O_3_0_0(op_O_3_0_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
endmodule
module Passthrough(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_1_0_0,
  input  [15:0] I_2_0_0,
  input  [15:0] I_3_0_0,
  output [15:0] O_0_0,
  output [15:0] O_1_0,
  output [15:0] O_2_0,
  output [15:0] O_3_0
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0 = I_0_0_0; // @[Passthrough.scala 17:68]
  assign O_1_0 = I_1_0_0; // @[Passthrough.scala 17:68]
  assign O_2_0 = I_2_0_0; // @[Passthrough.scala 17:68]
  assign O_3_0 = I_3_0_0; // @[Passthrough.scala 17:68]
endmodule
module Passthrough_1(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_1_0,
  input  [15:0] I_2_0,
  input  [15:0] I_3_0,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0 = I_0_0; // @[Passthrough.scala 17:68]
  assign O_1 = I_1_0; // @[Passthrough.scala 17:68]
  assign O_2 = I_2_0; // @[Passthrough.scala 17:68]
  assign O_3 = I_3_0; // @[Passthrough.scala 17:68]
endmodule
module PartitionS_4(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_3_0,
  input  [15:0] I_3_1,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0 = I_0_0; // @[Partition.scala 15:39]
  assign O_0_0_1 = I_0_1; // @[Partition.scala 15:39]
  assign O_1_0_0 = I_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1 = I_1_1; // @[Partition.scala 15:39]
  assign O_2_0_0 = I_2_0; // @[Partition.scala 15:39]
  assign O_2_0_1 = I_2_1; // @[Partition.scala 15:39]
  assign O_3_0_0 = I_3_0; // @[Partition.scala 15:39]
  assign O_3_0_1 = I_3_1; // @[Partition.scala 15:39]
endmodule
module MapT_9(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_3_0,
  input  [15:0] I_3_1,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1; // @[MapT.scala 8:20]
  PartitionS_4 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0(op_I_0_0),
    .I_0_1(op_I_0_1),
    .I_1_0(op_I_1_0),
    .I_1_1(op_I_1_1),
    .I_2_0(op_I_2_0),
    .I_2_1(op_I_2_1),
    .I_3_0(op_I_3_0),
    .I_3_1(op_I_3_1),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0 = I_0_0; // @[MapT.scala 14:10]
  assign op_I_0_1 = I_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0 = I_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1 = I_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0 = I_2_0; // @[MapT.scala 14:10]
  assign op_I_2_1 = I_2_1; // @[MapT.scala 14:10]
  assign op_I_3_0 = I_3_0; // @[MapT.scala 14:10]
  assign op_I_3_1 = I_3_1; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq_4(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  output [15:0] O_0,
  output [15:0] O_1
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0 = I_0; // @[Tuple.scala 41:5]
  assign O_1 = I_1; // @[Tuple.scala 41:5]
endmodule
module Remove1S_4(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  output [15:0] O_0,
  output [15:0] O_1
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_1; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_4 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0(op_inst_I_0),
    .I_1(op_inst_I_1),
    .O_0(op_inst_O_0),
    .O_1(op_inst_O_1)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0 = op_inst_O_0; // @[Remove1S.scala 14:5]
  assign O_1 = op_inst_O_1; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0 = I_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1 = I_0_1; // @[Remove1S.scala 13:13]
endmodule
module MapS_10(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_3_0,
  output [15:0] O_3_1
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_1; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  Remove1S_4 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  Remove1S_4 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1)
  );
  Remove1S_4 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1)
  );
  Remove1S_4 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_3_0 = other_ops_2_O_0; // @[MapS.scala 21:12]
  assign O_3_1 = other_ops_2_O_1; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
endmodule
module MapT_10(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_3_0,
  output [15:0] O_3_1
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_1; // @[MapT.scala 8:20]
  MapS_10 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0 = op_O_0_0; // @[MapT.scala 15:7]
  assign O_0_1 = op_O_0_1; // @[MapT.scala 15:7]
  assign O_1_0 = op_O_1_0; // @[MapT.scala 15:7]
  assign O_1_1 = op_O_1_1; // @[MapT.scala 15:7]
  assign O_2_0 = op_O_2_0; // @[MapT.scala 15:7]
  assign O_2_1 = op_O_2_1; // @[MapT.scala 15:7]
  assign O_3_0 = op_O_3_0; // @[MapT.scala 15:7]
  assign O_3_1 = op_O_3_1; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
endmodule
module SSeqTupleCreator_6(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_1_0,
  output [15:0] O_1_1
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0_0 = I0_0; // @[Tuple.scala 12:32]
  assign O_0_1 = I0_1; // @[Tuple.scala 12:32]
  assign O_1_0 = I1_0; // @[Tuple.scala 13:32]
  assign O_1_1 = I1_1; // @[Tuple.scala 13:32]
endmodule
module Map2S_14(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_3_0,
  input  [15:0] I0_3_1,
  input  [15:0] I1_0_0,
  input  [15:0] I1_0_1,
  input  [15:0] I1_1_0,
  input  [15:0] I1_1_1,
  input  [15:0] I1_2_0,
  input  [15:0] I1_2_1,
  input  [15:0] I1_3_0,
  input  [15:0] I1_3_1,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  SSeqTupleCreator_6 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
endmodule
module Map2T_10(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_3_0,
  input  [15:0] I0_3_1,
  input  [15:0] I1_0_0,
  input  [15:0] I1_0_1,
  input  [15:0] I1_1_0,
  input  [15:0] I1_1_1,
  input  [15:0] I1_2_0,
  input  [15:0] I1_2_1,
  input  [15:0] I1_3_0,
  input  [15:0] I1_3_1,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_1; // @[Map2T.scala 8:20]
  Map2S_14 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I0_2_0(op_I0_2_0),
    .I0_2_1(op_I0_2_1),
    .I0_3_0(op_I0_3_0),
    .I0_3_1(op_I0_3_1),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_2_0(op_I1_2_0),
    .I1_2_1(op_I1_2_1),
    .I1_3_0(op_I1_3_0),
    .I1_3_1(op_I1_3_1),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_2_0_0 = op_O_2_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_1 = op_O_2_0_1; // @[Map2T.scala 17:7]
  assign O_2_1_0 = op_O_2_1_0; // @[Map2T.scala 17:7]
  assign O_2_1_1 = op_O_2_1_1; // @[Map2T.scala 17:7]
  assign O_3_0_0 = op_O_3_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_1 = op_O_3_0_1; // @[Map2T.scala 17:7]
  assign O_3_1_0 = op_O_3_1_0; // @[Map2T.scala 17:7]
  assign O_3_1_1 = op_O_3_1_1; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0 = I0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1 = I0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0 = I0_3_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1 = I0_3_1; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_2_0 = I1_2_0; // @[Map2T.scala 16:11]
  assign op_I1_2_1 = I1_2_1; // @[Map2T.scala 16:11]
  assign op_I1_3_0 = I1_3_0; // @[Map2T.scala 16:11]
  assign op_I1_3_1 = I1_3_1; // @[Map2T.scala 16:11]
endmodule
module PartitionS_6(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  output [15:0] O_0_0_0_0,
  output [15:0] O_0_0_0_1,
  output [15:0] O_0_0_1_0,
  output [15:0] O_0_0_1_1,
  output [15:0] O_1_0_0_0,
  output [15:0] O_1_0_0_1,
  output [15:0] O_1_0_1_0,
  output [15:0] O_1_0_1_1,
  output [15:0] O_2_0_0_0,
  output [15:0] O_2_0_0_1,
  output [15:0] O_2_0_1_0,
  output [15:0] O_2_0_1_1,
  output [15:0] O_3_0_0_0,
  output [15:0] O_3_0_0_1,
  output [15:0] O_3_0_1_0,
  output [15:0] O_3_0_1_1
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0_0 = I_0_0_0; // @[Partition.scala 15:39]
  assign O_0_0_0_1 = I_0_0_1; // @[Partition.scala 15:39]
  assign O_0_0_1_0 = I_0_1_0; // @[Partition.scala 15:39]
  assign O_0_0_1_1 = I_0_1_1; // @[Partition.scala 15:39]
  assign O_1_0_0_0 = I_1_0_0; // @[Partition.scala 15:39]
  assign O_1_0_0_1 = I_1_0_1; // @[Partition.scala 15:39]
  assign O_1_0_1_0 = I_1_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1_1 = I_1_1_1; // @[Partition.scala 15:39]
  assign O_2_0_0_0 = I_2_0_0; // @[Partition.scala 15:39]
  assign O_2_0_0_1 = I_2_0_1; // @[Partition.scala 15:39]
  assign O_2_0_1_0 = I_2_1_0; // @[Partition.scala 15:39]
  assign O_2_0_1_1 = I_2_1_1; // @[Partition.scala 15:39]
  assign O_3_0_0_0 = I_3_0_0; // @[Partition.scala 15:39]
  assign O_3_0_0_1 = I_3_0_1; // @[Partition.scala 15:39]
  assign O_3_0_1_0 = I_3_1_0; // @[Partition.scala 15:39]
  assign O_3_0_1_1 = I_3_1_1; // @[Partition.scala 15:39]
endmodule
module MapT_13(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  output [15:0] O_0_0_0_0,
  output [15:0] O_0_0_0_1,
  output [15:0] O_0_0_1_0,
  output [15:0] O_0_0_1_1,
  output [15:0] O_1_0_0_0,
  output [15:0] O_1_0_0_1,
  output [15:0] O_1_0_1_0,
  output [15:0] O_1_0_1_1,
  output [15:0] O_2_0_0_0,
  output [15:0] O_2_0_0_1,
  output [15:0] O_2_0_1_0,
  output [15:0] O_2_0_1_1,
  output [15:0] O_3_0_0_0,
  output [15:0] O_3_0_0_1,
  output [15:0] O_3_0_1_0,
  output [15:0] O_3_0_1_1
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1_1; // @[MapT.scala 8:20]
  PartitionS_6 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_0_0_1_0(op_O_0_0_1_0),
    .O_0_0_1_1(op_O_0_0_1_1),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_1_0_1_0(op_O_1_0_1_0),
    .O_1_0_1_1(op_O_1_0_1_1),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_2_0_1_0(op_O_2_0_1_0),
    .O_2_0_1_1(op_O_2_0_1_1),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_3_0_1_0(op_O_3_0_1_0),
    .O_3_0_1_1(op_O_3_0_1_1)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_1_0 = op_O_0_0_1_0; // @[MapT.scala 15:7]
  assign O_0_0_1_1 = op_O_0_0_1_1; // @[MapT.scala 15:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[MapT.scala 15:7]
  assign O_1_0_1_0 = op_O_1_0_1_0; // @[MapT.scala 15:7]
  assign O_1_0_1_1 = op_O_1_0_1_1; // @[MapT.scala 15:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[MapT.scala 15:7]
  assign O_2_0_1_0 = op_O_2_0_1_0; // @[MapT.scala 15:7]
  assign O_2_0_1_1 = op_O_2_0_1_1; // @[MapT.scala 15:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[MapT.scala 15:7]
  assign O_3_0_1_0 = op_O_3_0_1_0; // @[MapT.scala 15:7]
  assign O_3_0_1_1 = op_O_3_0_1_1; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq_6(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_1_0,
  output [15:0] O_1_1
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0_0 = I_0_0; // @[Tuple.scala 41:5]
  assign O_0_1 = I_0_1; // @[Tuple.scala 41:5]
  assign O_1_0 = I_1_0; // @[Tuple.scala 41:5]
  assign O_1_1 = I_1_1; // @[Tuple.scala 41:5]
endmodule
module Remove1S_6(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_1_0,
  output [15:0] O_1_1
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_0_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_0_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_1_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_1_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_0_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_0_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_1_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_1_1; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_6 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0_0(op_inst_I_0_0),
    .I_0_1(op_inst_I_0_1),
    .I_1_0(op_inst_I_1_0),
    .I_1_1(op_inst_I_1_1),
    .O_0_0(op_inst_O_0_0),
    .O_0_1(op_inst_O_0_1),
    .O_1_0(op_inst_O_1_0),
    .O_1_1(op_inst_O_1_1)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0_0 = op_inst_O_0_0; // @[Remove1S.scala 14:5]
  assign O_0_1 = op_inst_O_0_1; // @[Remove1S.scala 14:5]
  assign O_1_0 = op_inst_O_1_0; // @[Remove1S.scala 14:5]
  assign O_1_1 = op_inst_O_1_1; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0_0 = I_0_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_1 = I_0_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_0 = I_0_1_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_1 = I_0_1_1; // @[Remove1S.scala 13:13]
endmodule
module MapS_12(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0_0,
  input  [15:0] I_0_0_0_1,
  input  [15:0] I_0_0_1_0,
  input  [15:0] I_0_0_1_1,
  input  [15:0] I_1_0_0_0,
  input  [15:0] I_1_0_0_1,
  input  [15:0] I_1_0_1_0,
  input  [15:0] I_1_0_1_1,
  input  [15:0] I_2_0_0_0,
  input  [15:0] I_2_0_0_1,
  input  [15:0] I_2_0_1_0,
  input  [15:0] I_2_0_1_1,
  input  [15:0] I_3_0_0_0,
  input  [15:0] I_3_0_0_1,
  input  [15:0] I_3_0_1_0,
  input  [15:0] I_3_0_1_1,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1_1; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_1_1; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  Remove1S_6 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0_0(fst_op_I_0_0_0),
    .I_0_0_1(fst_op_I_0_0_1),
    .I_0_1_0(fst_op_I_0_1_0),
    .I_0_1_1(fst_op_I_0_1_1),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1)
  );
  Remove1S_6 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0_0(other_ops_0_I_0_0_0),
    .I_0_0_1(other_ops_0_I_0_0_1),
    .I_0_1_0(other_ops_0_I_0_1_0),
    .I_0_1_1(other_ops_0_I_0_1_1),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1)
  );
  Remove1S_6 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0_0(other_ops_1_I_0_0_0),
    .I_0_0_1(other_ops_1_I_0_0_1),
    .I_0_1_0(other_ops_1_I_0_1_0),
    .I_0_1_1(other_ops_1_I_0_1_1),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1)
  );
  Remove1S_6 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0_0(other_ops_2_I_0_0_0),
    .I_0_0_1(other_ops_2_I_0_0_1),
    .I_0_1_0(other_ops_2_I_0_1_0),
    .I_0_1_1(other_ops_2_I_0_1_1),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[MapS.scala 17:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[MapS.scala 17:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[MapS.scala 21:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[MapS.scala 21:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[MapS.scala 21:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[MapS.scala 21:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[MapS.scala 21:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[MapS.scala 21:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0_0 = I_0_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_1 = I_0_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_0 = I_0_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_1 = I_0_0_1_1; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0_0 = I_1_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_1 = I_1_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_0 = I_1_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_1 = I_1_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0_0 = I_2_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_1 = I_2_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_0 = I_2_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_1 = I_2_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0_0 = I_3_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_1 = I_3_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_0 = I_3_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_1 = I_3_0_1_1; // @[MapS.scala 20:41]
endmodule
module MapT_14(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0_0,
  input  [15:0] I_0_0_0_1,
  input  [15:0] I_0_0_1_0,
  input  [15:0] I_0_0_1_1,
  input  [15:0] I_1_0_0_0,
  input  [15:0] I_1_0_0_1,
  input  [15:0] I_1_0_1_0,
  input  [15:0] I_1_0_1_1,
  input  [15:0] I_2_0_0_0,
  input  [15:0] I_2_0_0_1,
  input  [15:0] I_2_0_1_0,
  input  [15:0] I_2_0_1_1,
  input  [15:0] I_3_0_0_0,
  input  [15:0] I_3_0_0_1,
  input  [15:0] I_3_0_1_0,
  input  [15:0] I_3_0_1_1,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_1_1; // @[MapT.scala 8:20]
  MapS_12 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0_0(op_I_0_0_0_0),
    .I_0_0_0_1(op_I_0_0_0_1),
    .I_0_0_1_0(op_I_0_0_1_0),
    .I_0_0_1_1(op_I_0_0_1_1),
    .I_1_0_0_0(op_I_1_0_0_0),
    .I_1_0_0_1(op_I_1_0_0_1),
    .I_1_0_1_0(op_I_1_0_1_0),
    .I_1_0_1_1(op_I_1_0_1_1),
    .I_2_0_0_0(op_I_2_0_0_0),
    .I_2_0_0_1(op_I_2_0_0_1),
    .I_2_0_1_0(op_I_2_0_1_0),
    .I_2_0_1_1(op_I_2_0_1_1),
    .I_3_0_0_0(op_I_3_0_0_0),
    .I_3_0_0_1(op_I_3_0_0_1),
    .I_3_0_1_0(op_I_3_0_1_0),
    .I_3_0_1_1(op_I_3_0_1_1),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_1_0 = op_O_0_1_0; // @[MapT.scala 15:7]
  assign O_0_1_1 = op_O_0_1_1; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_1_0 = op_O_1_1_0; // @[MapT.scala 15:7]
  assign O_1_1_1 = op_O_1_1_1; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_1_0 = op_O_2_1_0; // @[MapT.scala 15:7]
  assign O_2_1_1 = op_O_2_1_1; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_1_0 = op_O_3_1_0; // @[MapT.scala 15:7]
  assign O_3_1_1 = op_O_3_1_1; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0_0 = I_0_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_0_1 = I_0_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_1_0 = I_0_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1_1 = I_0_0_1_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0_0 = I_1_0_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_0_1 = I_1_0_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_1_0 = I_1_0_1_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1_1 = I_1_0_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0_0 = I_2_0_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_0_1 = I_2_0_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_1_0 = I_2_0_1_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1_1 = I_2_0_1_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0_0 = I_3_0_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_0_1 = I_3_0_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_1_0 = I_3_0_1_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1_1 = I_3_0_1_1; // @[MapT.scala 14:10]
endmodule
module InitialDelayCounter_2(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [3:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [3:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 4'hb; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 4'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 4'hb; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 4'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Map2S_15(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  output [15:0] O_0_t0b,
  output [15:0] O_0_t1b,
  output [15:0] O_1_t0b,
  output [15:0] O_1_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  AtomTuple other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
endmodule
module Map2S_16(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  output [15:0] O_0_0_t0b,
  output [15:0] O_0_0_t1b,
  output [15:0] O_0_1_t0b,
  output [15:0] O_0_1_t1b,
  output [15:0] O_1_0_t0b,
  output [15:0] O_1_0_t1b,
  output [15:0] O_1_1_t0b,
  output [15:0] O_1_1_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_t0b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_t1b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_t0b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_t1b; // @[Map2S.scala 10:86]
  Map2S_15 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b),
    .O_1_t0b(fst_op_O_1_t0b),
    .O_1_t1b(fst_op_O_1_t1b)
  );
  Map2S_15 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .O_0_t0b(other_ops_0_O_0_t0b),
    .O_0_t1b(other_ops_0_O_0_t1b),
    .O_1_t0b(other_ops_0_O_1_t0b),
    .O_1_t1b(other_ops_0_O_1_t1b)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign O_0_1_t0b = fst_op_O_1_t0b; // @[Map2S.scala 19:8]
  assign O_0_1_t1b = fst_op_O_1_t1b; // @[Map2S.scala 19:8]
  assign O_1_0_t0b = other_ops_0_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_1_0_t1b = other_ops_0_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_1_1_t0b = other_ops_0_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_1_1_t1b = other_ops_0_O_1_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = 16'h1; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = 16'h4; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = 16'h2; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = 16'h1; // @[Map2S.scala 23:43]
endmodule
module MapS_13(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_t0b,
  input  [15:0] I_0_t1b,
  input  [15:0] I_1_t0b,
  input  [15:0] I_1_t1b,
  output [15:0] O_0,
  output [15:0] O_1
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O; // @[MapS.scala 10:86]
  Mul fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  Mul other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t0b(other_ops_0_I_t0b),
    .I_t1b(other_ops_0_I_t1b),
    .O(other_ops_0_O)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t0b = I_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_t1b = I_1_t1b; // @[MapS.scala 20:41]
endmodule
module MapS_14(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_t0b,
  input  [15:0] I_0_0_t1b,
  input  [15:0] I_0_1_t0b,
  input  [15:0] I_0_1_t1b,
  input  [15:0] I_1_0_t0b,
  input  [15:0] I_1_0_t1b,
  input  [15:0] I_1_1_t0b,
  input  [15:0] I_1_1_t1b,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_1_0,
  output [15:0] O_1_1
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_t0b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_t0b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  MapS_13 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .I_1_t0b(fst_op_I_1_t0b),
    .I_1_t1b(fst_op_I_1_t1b),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  MapS_13 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_t0b(other_ops_0_I_0_t0b),
    .I_0_t1b(other_ops_0_I_0_t1b),
    .I_1_t0b(other_ops_0_I_1_t0b),
    .I_1_t1b(other_ops_0_I_1_t1b),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t0b = I_0_1_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t1b = I_0_1_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_t0b = I_1_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_t1b = I_1_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t0b = I_1_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t1b = I_1_1_t1b; // @[MapS.scala 20:41]
endmodule
module ReduceS_2(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  output [15:0] O_0
);
  wire [15:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  reg [15:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [15:0] _T_1; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [15:0] _T_2; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg  _T_3; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_4;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  assign valid_down = _T_4; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = _T_2; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = _T_1; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    _T_1 <= I_0;
    _T_2 <= I_1;
    if (reset) begin
      _T_3 <= 1'h0;
    end else begin
      _T_3 <= valid_up;
    end
    _T_4 <= _T_3;
  end
endmodule
module MapS_15(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  output [15:0] O_0_0,
  output [15:0] O_1_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  ReduceS_2 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .O_0(fst_op_O_0)
  );
  ReduceS_2 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0(other_ops_0_I_0),
    .I_1(other_ops_0_I_1),
    .O_0(other_ops_0_O_0)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0 = I_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1 = I_1_1; // @[MapS.scala 20:41]
endmodule
module ReduceS_3(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_1_0,
  output [15:0] O_0_0
);
  wire [15:0] MapSNoValid_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_O_0; // @[ReduceS.scala 20:43]
  reg [15:0] _T_0; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [15:0] _T_1_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [15:0] _T_2_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg  _T_3; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_4;
  MapSNoValid MapSNoValid ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_I_0_t0b),
    .I_0_t1b(MapSNoValid_I_0_t1b),
    .O_0(MapSNoValid_O_0)
  );
  assign valid_down = _T_4; // @[ReduceS.scala 47:14]
  assign O_0_0 = _T_0; // @[ReduceS.scala 27:14]
  assign MapSNoValid_I_0_t0b = _T_1_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_I_0_t1b = _T_2_0; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1_0 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2_0 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= MapSNoValid_O_0;
    _T_1_0 <= I_0_0;
    _T_2_0 <= I_1_0;
    if (reset) begin
      _T_3 <= 1'h0;
    end else begin
      _T_3 <= valid_up;
    end
    _T_4 <= _T_3;
  end
endmodule
module InitialDelayCounter_3(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [4:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [4:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 5'h12; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 5'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 5'h12; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 5'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Module_1(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  output [15:0] O_0_0
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n208_valid_up; // @[Top.scala 47:22]
  wire  n208_valid_down; // @[Top.scala 47:22]
  wire [15:0] n208_I0_0_0; // @[Top.scala 47:22]
  wire [15:0] n208_I0_0_1; // @[Top.scala 47:22]
  wire [15:0] n208_I0_1_0; // @[Top.scala 47:22]
  wire [15:0] n208_I0_1_1; // @[Top.scala 47:22]
  wire [15:0] n208_O_0_0_t0b; // @[Top.scala 47:22]
  wire [15:0] n208_O_0_0_t1b; // @[Top.scala 47:22]
  wire [15:0] n208_O_0_1_t0b; // @[Top.scala 47:22]
  wire [15:0] n208_O_0_1_t1b; // @[Top.scala 47:22]
  wire [15:0] n208_O_1_0_t0b; // @[Top.scala 47:22]
  wire [15:0] n208_O_1_0_t1b; // @[Top.scala 47:22]
  wire [15:0] n208_O_1_1_t0b; // @[Top.scala 47:22]
  wire [15:0] n208_O_1_1_t1b; // @[Top.scala 47:22]
  wire  n219_clock; // @[Top.scala 51:22]
  wire  n219_reset; // @[Top.scala 51:22]
  wire  n219_valid_up; // @[Top.scala 51:22]
  wire  n219_valid_down; // @[Top.scala 51:22]
  wire [15:0] n219_I_0_0_t0b; // @[Top.scala 51:22]
  wire [15:0] n219_I_0_0_t1b; // @[Top.scala 51:22]
  wire [15:0] n219_I_0_1_t0b; // @[Top.scala 51:22]
  wire [15:0] n219_I_0_1_t1b; // @[Top.scala 51:22]
  wire [15:0] n219_I_1_0_t0b; // @[Top.scala 51:22]
  wire [15:0] n219_I_1_0_t1b; // @[Top.scala 51:22]
  wire [15:0] n219_I_1_1_t0b; // @[Top.scala 51:22]
  wire [15:0] n219_I_1_1_t1b; // @[Top.scala 51:22]
  wire [15:0] n219_O_0_0; // @[Top.scala 51:22]
  wire [15:0] n219_O_0_1; // @[Top.scala 51:22]
  wire [15:0] n219_O_1_0; // @[Top.scala 51:22]
  wire [15:0] n219_O_1_1; // @[Top.scala 51:22]
  wire  n224_clock; // @[Top.scala 54:22]
  wire  n224_reset; // @[Top.scala 54:22]
  wire  n224_valid_up; // @[Top.scala 54:22]
  wire  n224_valid_down; // @[Top.scala 54:22]
  wire [15:0] n224_I_0_0; // @[Top.scala 54:22]
  wire [15:0] n224_I_0_1; // @[Top.scala 54:22]
  wire [15:0] n224_I_1_0; // @[Top.scala 54:22]
  wire [15:0] n224_I_1_1; // @[Top.scala 54:22]
  wire [15:0] n224_O_0_0; // @[Top.scala 54:22]
  wire [15:0] n224_O_1_0; // @[Top.scala 54:22]
  wire  n229_clock; // @[Top.scala 57:22]
  wire  n229_reset; // @[Top.scala 57:22]
  wire  n229_valid_up; // @[Top.scala 57:22]
  wire  n229_valid_down; // @[Top.scala 57:22]
  wire [15:0] n229_I_0_0; // @[Top.scala 57:22]
  wire [15:0] n229_I_1_0; // @[Top.scala 57:22]
  wire [15:0] n229_O_0_0; // @[Top.scala 57:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n232_valid_up; // @[Top.scala 61:22]
  wire  n232_valid_down; // @[Top.scala 61:22]
  wire [15:0] n232_I0_0_0; // @[Top.scala 61:22]
  wire [7:0] n232_I1_0_0; // @[Top.scala 61:22]
  wire [15:0] n232_O_0_0_t0b; // @[Top.scala 61:22]
  wire [7:0] n232_O_0_0_t1b; // @[Top.scala 61:22]
  wire  n243_clock; // @[Top.scala 65:22]
  wire  n243_reset; // @[Top.scala 65:22]
  wire  n243_valid_up; // @[Top.scala 65:22]
  wire  n243_valid_down; // @[Top.scala 65:22]
  wire [15:0] n243_I_0_0_t0b; // @[Top.scala 65:22]
  wire [7:0] n243_I_0_0_t1b; // @[Top.scala 65:22]
  wire [15:0] n243_O_0_0; // @[Top.scala 65:22]
  InitialDelayCounter_2 InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  Map2S_16 n208 ( // @[Top.scala 47:22]
    .valid_up(n208_valid_up),
    .valid_down(n208_valid_down),
    .I0_0_0(n208_I0_0_0),
    .I0_0_1(n208_I0_0_1),
    .I0_1_0(n208_I0_1_0),
    .I0_1_1(n208_I0_1_1),
    .O_0_0_t0b(n208_O_0_0_t0b),
    .O_0_0_t1b(n208_O_0_0_t1b),
    .O_0_1_t0b(n208_O_0_1_t0b),
    .O_0_1_t1b(n208_O_0_1_t1b),
    .O_1_0_t0b(n208_O_1_0_t0b),
    .O_1_0_t1b(n208_O_1_0_t1b),
    .O_1_1_t0b(n208_O_1_1_t0b),
    .O_1_1_t1b(n208_O_1_1_t1b)
  );
  MapS_14 n219 ( // @[Top.scala 51:22]
    .clock(n219_clock),
    .reset(n219_reset),
    .valid_up(n219_valid_up),
    .valid_down(n219_valid_down),
    .I_0_0_t0b(n219_I_0_0_t0b),
    .I_0_0_t1b(n219_I_0_0_t1b),
    .I_0_1_t0b(n219_I_0_1_t0b),
    .I_0_1_t1b(n219_I_0_1_t1b),
    .I_1_0_t0b(n219_I_1_0_t0b),
    .I_1_0_t1b(n219_I_1_0_t1b),
    .I_1_1_t0b(n219_I_1_1_t0b),
    .I_1_1_t1b(n219_I_1_1_t1b),
    .O_0_0(n219_O_0_0),
    .O_0_1(n219_O_0_1),
    .O_1_0(n219_O_1_0),
    .O_1_1(n219_O_1_1)
  );
  MapS_15 n224 ( // @[Top.scala 54:22]
    .clock(n224_clock),
    .reset(n224_reset),
    .valid_up(n224_valid_up),
    .valid_down(n224_valid_down),
    .I_0_0(n224_I_0_0),
    .I_0_1(n224_I_0_1),
    .I_1_0(n224_I_1_0),
    .I_1_1(n224_I_1_1),
    .O_0_0(n224_O_0_0),
    .O_1_0(n224_O_1_0)
  );
  ReduceS_3 n229 ( // @[Top.scala 57:22]
    .clock(n229_clock),
    .reset(n229_reset),
    .valid_up(n229_valid_up),
    .valid_down(n229_valid_down),
    .I_0_0(n229_I_0_0),
    .I_1_0(n229_I_1_0),
    .O_0_0(n229_O_0_0)
  );
  InitialDelayCounter_3 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  Map2S_11 n232 ( // @[Top.scala 61:22]
    .valid_up(n232_valid_up),
    .valid_down(n232_valid_down),
    .I0_0_0(n232_I0_0_0),
    .I1_0_0(n232_I1_0_0),
    .O_0_0_t0b(n232_O_0_0_t0b),
    .O_0_0_t1b(n232_O_0_0_t1b)
  );
  MapS_8 n243 ( // @[Top.scala 65:22]
    .clock(n243_clock),
    .reset(n243_reset),
    .valid_up(n243_valid_up),
    .valid_down(n243_valid_down),
    .I_0_0_t0b(n243_I_0_0_t0b),
    .I_0_0_t1b(n243_I_0_0_t1b),
    .O_0_0(n243_O_0_0)
  );
  assign valid_down = n243_valid_down; // @[Top.scala 69:16]
  assign O_0_0 = n243_O_0_0; // @[Top.scala 68:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n208_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 50:19]
  assign n208_I0_0_0 = I_0_0; // @[Top.scala 48:13]
  assign n208_I0_0_1 = I_0_1; // @[Top.scala 48:13]
  assign n208_I0_1_0 = I_1_0; // @[Top.scala 48:13]
  assign n208_I0_1_1 = I_1_1; // @[Top.scala 48:13]
  assign n219_clock = clock;
  assign n219_reset = reset;
  assign n219_valid_up = n208_valid_down; // @[Top.scala 53:19]
  assign n219_I_0_0_t0b = n208_O_0_0_t0b; // @[Top.scala 52:12]
  assign n219_I_0_0_t1b = n208_O_0_0_t1b; // @[Top.scala 52:12]
  assign n219_I_0_1_t0b = n208_O_0_1_t0b; // @[Top.scala 52:12]
  assign n219_I_0_1_t1b = n208_O_0_1_t1b; // @[Top.scala 52:12]
  assign n219_I_1_0_t0b = n208_O_1_0_t0b; // @[Top.scala 52:12]
  assign n219_I_1_0_t1b = n208_O_1_0_t1b; // @[Top.scala 52:12]
  assign n219_I_1_1_t0b = n208_O_1_1_t0b; // @[Top.scala 52:12]
  assign n219_I_1_1_t1b = n208_O_1_1_t1b; // @[Top.scala 52:12]
  assign n224_clock = clock;
  assign n224_reset = reset;
  assign n224_valid_up = n219_valid_down; // @[Top.scala 56:19]
  assign n224_I_0_0 = n219_O_0_0; // @[Top.scala 55:12]
  assign n224_I_0_1 = n219_O_0_1; // @[Top.scala 55:12]
  assign n224_I_1_0 = n219_O_1_0; // @[Top.scala 55:12]
  assign n224_I_1_1 = n219_O_1_1; // @[Top.scala 55:12]
  assign n229_clock = clock;
  assign n229_reset = reset;
  assign n229_valid_up = n224_valid_down; // @[Top.scala 59:19]
  assign n229_I_0_0 = n224_O_0_0; // @[Top.scala 58:12]
  assign n229_I_1_0 = n224_O_1_0; // @[Top.scala 58:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n232_valid_up = n229_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 64:19]
  assign n232_I0_0_0 = n229_O_0_0; // @[Top.scala 62:13]
  assign n232_I1_0_0 = 8'sh10; // @[Top.scala 63:13]
  assign n243_clock = clock;
  assign n243_reset = reset;
  assign n243_valid_up = n232_valid_down; // @[Top.scala 67:19]
  assign n243_I_0_0_t0b = n232_O_0_0_t0b; // @[Top.scala 66:12]
  assign n243_I_0_0_t1b = n232_O_0_0_t1b; // @[Top.scala 66:12]
endmodule
module MapS_18(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  output [15:0] O_0_0_0,
  output [15:0] O_1_0_0,
  output [15:0] O_2_0_0,
  output [15:0] O_3_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_2_clock; // @[MapS.scala 10:86]
  wire  other_ops_2_reset; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  Module_1 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_1_0(fst_op_I_1_0),
    .I_1_1(fst_op_I_1_1),
    .O_0_0(fst_op_O_0_0)
  );
  Module_1 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_1_0(other_ops_0_I_1_0),
    .I_1_1(other_ops_0_I_1_1),
    .O_0_0(other_ops_0_O_0_0)
  );
  Module_1 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_1_0(other_ops_1_I_1_0),
    .I_1_1(other_ops_1_I_1_1),
    .O_0_0(other_ops_1_O_0_0)
  );
  Module_1 other_ops_2 ( // @[MapS.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_1_0(other_ops_2_I_1_0),
    .I_1_1(other_ops_2_I_1_1),
    .O_0_0(other_ops_2_O_0_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_1_0 = I_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_1_1 = I_0_1_1; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_0 = I_1_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_1 = I_1_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_0 = I_2_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_1 = I_2_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_2_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_0 = I_3_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_1 = I_3_1_1; // @[MapS.scala 20:41]
endmodule
module MapT_15(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  output [15:0] O_0_0_0,
  output [15:0] O_1_0_0,
  output [15:0] O_2_0_0,
  output [15:0] O_3_0_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[MapT.scala 8:20]
  MapS_18 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .O_0_0_0(op_O_0_0_0),
    .O_1_0_0(op_O_1_0_0),
    .O_2_0_0(op_O_2_0_0),
    .O_3_0_0(op_O_3_0_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
endmodule
module Top(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  input  [15:0] I_3,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3
);
  wire  n1_clock; // @[Top.scala 75:20]
  wire  n1_reset; // @[Top.scala 75:20]
  wire  n1_valid_up; // @[Top.scala 75:20]
  wire  n1_valid_down; // @[Top.scala 75:20]
  wire [15:0] n1_I_0; // @[Top.scala 75:20]
  wire [15:0] n1_I_1; // @[Top.scala 75:20]
  wire [15:0] n1_I_2; // @[Top.scala 75:20]
  wire [15:0] n1_I_3; // @[Top.scala 75:20]
  wire [15:0] n1_O_0; // @[Top.scala 75:20]
  wire [15:0] n1_O_1; // @[Top.scala 75:20]
  wire [15:0] n1_O_2; // @[Top.scala 75:20]
  wire [15:0] n1_O_3; // @[Top.scala 75:20]
  wire  n2_clock; // @[Top.scala 78:20]
  wire  n2_reset; // @[Top.scala 78:20]
  wire  n2_valid_up; // @[Top.scala 78:20]
  wire  n2_valid_down; // @[Top.scala 78:20]
  wire [15:0] n2_I_0; // @[Top.scala 78:20]
  wire [15:0] n2_I_1; // @[Top.scala 78:20]
  wire [15:0] n2_I_2; // @[Top.scala 78:20]
  wire [15:0] n2_I_3; // @[Top.scala 78:20]
  wire [15:0] n2_O_0; // @[Top.scala 78:20]
  wire [15:0] n2_O_1; // @[Top.scala 78:20]
  wire [15:0] n2_O_2; // @[Top.scala 78:20]
  wire [15:0] n2_O_3; // @[Top.scala 78:20]
  wire  n3_clock; // @[Top.scala 81:20]
  wire  n3_reset; // @[Top.scala 81:20]
  wire  n3_valid_up; // @[Top.scala 81:20]
  wire  n3_valid_down; // @[Top.scala 81:20]
  wire [15:0] n3_I_0; // @[Top.scala 81:20]
  wire [15:0] n3_I_1; // @[Top.scala 81:20]
  wire [15:0] n3_I_2; // @[Top.scala 81:20]
  wire [15:0] n3_I_3; // @[Top.scala 81:20]
  wire [15:0] n3_O_0; // @[Top.scala 81:20]
  wire [15:0] n3_O_1; // @[Top.scala 81:20]
  wire [15:0] n3_O_2; // @[Top.scala 81:20]
  wire [15:0] n3_O_3; // @[Top.scala 81:20]
  wire  n4_clock; // @[Top.scala 84:20]
  wire  n4_valid_up; // @[Top.scala 84:20]
  wire  n4_valid_down; // @[Top.scala 84:20]
  wire [15:0] n4_I_0; // @[Top.scala 84:20]
  wire [15:0] n4_I_1; // @[Top.scala 84:20]
  wire [15:0] n4_I_2; // @[Top.scala 84:20]
  wire [15:0] n4_I_3; // @[Top.scala 84:20]
  wire [15:0] n4_O_0; // @[Top.scala 84:20]
  wire [15:0] n4_O_1; // @[Top.scala 84:20]
  wire [15:0] n4_O_2; // @[Top.scala 84:20]
  wire [15:0] n4_O_3; // @[Top.scala 84:20]
  wire  n5_clock; // @[Top.scala 87:20]
  wire  n5_valid_up; // @[Top.scala 87:20]
  wire  n5_valid_down; // @[Top.scala 87:20]
  wire [15:0] n5_I_0; // @[Top.scala 87:20]
  wire [15:0] n5_I_1; // @[Top.scala 87:20]
  wire [15:0] n5_I_2; // @[Top.scala 87:20]
  wire [15:0] n5_I_3; // @[Top.scala 87:20]
  wire [15:0] n5_O_0; // @[Top.scala 87:20]
  wire [15:0] n5_O_1; // @[Top.scala 87:20]
  wire [15:0] n5_O_2; // @[Top.scala 87:20]
  wire [15:0] n5_O_3; // @[Top.scala 87:20]
  wire  n6_valid_up; // @[Top.scala 90:20]
  wire  n6_valid_down; // @[Top.scala 90:20]
  wire [15:0] n6_I0_0; // @[Top.scala 90:20]
  wire [15:0] n6_I0_1; // @[Top.scala 90:20]
  wire [15:0] n6_I0_2; // @[Top.scala 90:20]
  wire [15:0] n6_I0_3; // @[Top.scala 90:20]
  wire [15:0] n6_I1_0; // @[Top.scala 90:20]
  wire [15:0] n6_I1_1; // @[Top.scala 90:20]
  wire [15:0] n6_I1_2; // @[Top.scala 90:20]
  wire [15:0] n6_I1_3; // @[Top.scala 90:20]
  wire [15:0] n6_O_0_0; // @[Top.scala 90:20]
  wire [15:0] n6_O_0_1; // @[Top.scala 90:20]
  wire [15:0] n6_O_1_0; // @[Top.scala 90:20]
  wire [15:0] n6_O_1_1; // @[Top.scala 90:20]
  wire [15:0] n6_O_2_0; // @[Top.scala 90:20]
  wire [15:0] n6_O_2_1; // @[Top.scala 90:20]
  wire [15:0] n6_O_3_0; // @[Top.scala 90:20]
  wire [15:0] n6_O_3_1; // @[Top.scala 90:20]
  wire  n13_valid_up; // @[Top.scala 94:21]
  wire  n13_valid_down; // @[Top.scala 94:21]
  wire [15:0] n13_I0_0_0; // @[Top.scala 94:21]
  wire [15:0] n13_I0_0_1; // @[Top.scala 94:21]
  wire [15:0] n13_I0_1_0; // @[Top.scala 94:21]
  wire [15:0] n13_I0_1_1; // @[Top.scala 94:21]
  wire [15:0] n13_I0_2_0; // @[Top.scala 94:21]
  wire [15:0] n13_I0_2_1; // @[Top.scala 94:21]
  wire [15:0] n13_I0_3_0; // @[Top.scala 94:21]
  wire [15:0] n13_I0_3_1; // @[Top.scala 94:21]
  wire [15:0] n13_I1_0; // @[Top.scala 94:21]
  wire [15:0] n13_I1_1; // @[Top.scala 94:21]
  wire [15:0] n13_I1_2; // @[Top.scala 94:21]
  wire [15:0] n13_I1_3; // @[Top.scala 94:21]
  wire [15:0] n13_O_0_0; // @[Top.scala 94:21]
  wire [15:0] n13_O_0_1; // @[Top.scala 94:21]
  wire [15:0] n13_O_0_2; // @[Top.scala 94:21]
  wire [15:0] n13_O_1_0; // @[Top.scala 94:21]
  wire [15:0] n13_O_1_1; // @[Top.scala 94:21]
  wire [15:0] n13_O_1_2; // @[Top.scala 94:21]
  wire [15:0] n13_O_2_0; // @[Top.scala 94:21]
  wire [15:0] n13_O_2_1; // @[Top.scala 94:21]
  wire [15:0] n13_O_2_2; // @[Top.scala 94:21]
  wire [15:0] n13_O_3_0; // @[Top.scala 94:21]
  wire [15:0] n13_O_3_1; // @[Top.scala 94:21]
  wire [15:0] n13_O_3_2; // @[Top.scala 94:21]
  wire  n22_valid_up; // @[Top.scala 98:21]
  wire  n22_valid_down; // @[Top.scala 98:21]
  wire [15:0] n22_I_0_0; // @[Top.scala 98:21]
  wire [15:0] n22_I_0_1; // @[Top.scala 98:21]
  wire [15:0] n22_I_0_2; // @[Top.scala 98:21]
  wire [15:0] n22_I_1_0; // @[Top.scala 98:21]
  wire [15:0] n22_I_1_1; // @[Top.scala 98:21]
  wire [15:0] n22_I_1_2; // @[Top.scala 98:21]
  wire [15:0] n22_I_2_0; // @[Top.scala 98:21]
  wire [15:0] n22_I_2_1; // @[Top.scala 98:21]
  wire [15:0] n22_I_2_2; // @[Top.scala 98:21]
  wire [15:0] n22_I_3_0; // @[Top.scala 98:21]
  wire [15:0] n22_I_3_1; // @[Top.scala 98:21]
  wire [15:0] n22_I_3_2; // @[Top.scala 98:21]
  wire [15:0] n22_O_0_0_0; // @[Top.scala 98:21]
  wire [15:0] n22_O_0_0_1; // @[Top.scala 98:21]
  wire [15:0] n22_O_0_0_2; // @[Top.scala 98:21]
  wire [15:0] n22_O_1_0_0; // @[Top.scala 98:21]
  wire [15:0] n22_O_1_0_1; // @[Top.scala 98:21]
  wire [15:0] n22_O_1_0_2; // @[Top.scala 98:21]
  wire [15:0] n22_O_2_0_0; // @[Top.scala 98:21]
  wire [15:0] n22_O_2_0_1; // @[Top.scala 98:21]
  wire [15:0] n22_O_2_0_2; // @[Top.scala 98:21]
  wire [15:0] n22_O_3_0_0; // @[Top.scala 98:21]
  wire [15:0] n22_O_3_0_1; // @[Top.scala 98:21]
  wire [15:0] n22_O_3_0_2; // @[Top.scala 98:21]
  wire  n29_valid_up; // @[Top.scala 101:21]
  wire  n29_valid_down; // @[Top.scala 101:21]
  wire [15:0] n29_I_0_0_0; // @[Top.scala 101:21]
  wire [15:0] n29_I_0_0_1; // @[Top.scala 101:21]
  wire [15:0] n29_I_0_0_2; // @[Top.scala 101:21]
  wire [15:0] n29_I_1_0_0; // @[Top.scala 101:21]
  wire [15:0] n29_I_1_0_1; // @[Top.scala 101:21]
  wire [15:0] n29_I_1_0_2; // @[Top.scala 101:21]
  wire [15:0] n29_I_2_0_0; // @[Top.scala 101:21]
  wire [15:0] n29_I_2_0_1; // @[Top.scala 101:21]
  wire [15:0] n29_I_2_0_2; // @[Top.scala 101:21]
  wire [15:0] n29_I_3_0_0; // @[Top.scala 101:21]
  wire [15:0] n29_I_3_0_1; // @[Top.scala 101:21]
  wire [15:0] n29_I_3_0_2; // @[Top.scala 101:21]
  wire [15:0] n29_O_0_0; // @[Top.scala 101:21]
  wire [15:0] n29_O_0_1; // @[Top.scala 101:21]
  wire [15:0] n29_O_0_2; // @[Top.scala 101:21]
  wire [15:0] n29_O_1_0; // @[Top.scala 101:21]
  wire [15:0] n29_O_1_1; // @[Top.scala 101:21]
  wire [15:0] n29_O_1_2; // @[Top.scala 101:21]
  wire [15:0] n29_O_2_0; // @[Top.scala 101:21]
  wire [15:0] n29_O_2_1; // @[Top.scala 101:21]
  wire [15:0] n29_O_2_2; // @[Top.scala 101:21]
  wire [15:0] n29_O_3_0; // @[Top.scala 101:21]
  wire [15:0] n29_O_3_1; // @[Top.scala 101:21]
  wire [15:0] n29_O_3_2; // @[Top.scala 101:21]
  wire  n30_clock; // @[Top.scala 104:21]
  wire  n30_valid_up; // @[Top.scala 104:21]
  wire  n30_valid_down; // @[Top.scala 104:21]
  wire [15:0] n30_I_0; // @[Top.scala 104:21]
  wire [15:0] n30_I_1; // @[Top.scala 104:21]
  wire [15:0] n30_I_2; // @[Top.scala 104:21]
  wire [15:0] n30_I_3; // @[Top.scala 104:21]
  wire [15:0] n30_O_0; // @[Top.scala 104:21]
  wire [15:0] n30_O_1; // @[Top.scala 104:21]
  wire [15:0] n30_O_2; // @[Top.scala 104:21]
  wire [15:0] n30_O_3; // @[Top.scala 104:21]
  wire  n31_clock; // @[Top.scala 107:21]
  wire  n31_valid_up; // @[Top.scala 107:21]
  wire  n31_valid_down; // @[Top.scala 107:21]
  wire [15:0] n31_I_0; // @[Top.scala 107:21]
  wire [15:0] n31_I_1; // @[Top.scala 107:21]
  wire [15:0] n31_I_2; // @[Top.scala 107:21]
  wire [15:0] n31_I_3; // @[Top.scala 107:21]
  wire [15:0] n31_O_0; // @[Top.scala 107:21]
  wire [15:0] n31_O_1; // @[Top.scala 107:21]
  wire [15:0] n31_O_2; // @[Top.scala 107:21]
  wire [15:0] n31_O_3; // @[Top.scala 107:21]
  wire  n32_valid_up; // @[Top.scala 110:21]
  wire  n32_valid_down; // @[Top.scala 110:21]
  wire [15:0] n32_I0_0; // @[Top.scala 110:21]
  wire [15:0] n32_I0_1; // @[Top.scala 110:21]
  wire [15:0] n32_I0_2; // @[Top.scala 110:21]
  wire [15:0] n32_I0_3; // @[Top.scala 110:21]
  wire [15:0] n32_I1_0; // @[Top.scala 110:21]
  wire [15:0] n32_I1_1; // @[Top.scala 110:21]
  wire [15:0] n32_I1_2; // @[Top.scala 110:21]
  wire [15:0] n32_I1_3; // @[Top.scala 110:21]
  wire [15:0] n32_O_0_0; // @[Top.scala 110:21]
  wire [15:0] n32_O_0_1; // @[Top.scala 110:21]
  wire [15:0] n32_O_1_0; // @[Top.scala 110:21]
  wire [15:0] n32_O_1_1; // @[Top.scala 110:21]
  wire [15:0] n32_O_2_0; // @[Top.scala 110:21]
  wire [15:0] n32_O_2_1; // @[Top.scala 110:21]
  wire [15:0] n32_O_3_0; // @[Top.scala 110:21]
  wire [15:0] n32_O_3_1; // @[Top.scala 110:21]
  wire  n39_valid_up; // @[Top.scala 114:21]
  wire  n39_valid_down; // @[Top.scala 114:21]
  wire [15:0] n39_I0_0_0; // @[Top.scala 114:21]
  wire [15:0] n39_I0_0_1; // @[Top.scala 114:21]
  wire [15:0] n39_I0_1_0; // @[Top.scala 114:21]
  wire [15:0] n39_I0_1_1; // @[Top.scala 114:21]
  wire [15:0] n39_I0_2_0; // @[Top.scala 114:21]
  wire [15:0] n39_I0_2_1; // @[Top.scala 114:21]
  wire [15:0] n39_I0_3_0; // @[Top.scala 114:21]
  wire [15:0] n39_I0_3_1; // @[Top.scala 114:21]
  wire [15:0] n39_I1_0; // @[Top.scala 114:21]
  wire [15:0] n39_I1_1; // @[Top.scala 114:21]
  wire [15:0] n39_I1_2; // @[Top.scala 114:21]
  wire [15:0] n39_I1_3; // @[Top.scala 114:21]
  wire [15:0] n39_O_0_0; // @[Top.scala 114:21]
  wire [15:0] n39_O_0_1; // @[Top.scala 114:21]
  wire [15:0] n39_O_0_2; // @[Top.scala 114:21]
  wire [15:0] n39_O_1_0; // @[Top.scala 114:21]
  wire [15:0] n39_O_1_1; // @[Top.scala 114:21]
  wire [15:0] n39_O_1_2; // @[Top.scala 114:21]
  wire [15:0] n39_O_2_0; // @[Top.scala 114:21]
  wire [15:0] n39_O_2_1; // @[Top.scala 114:21]
  wire [15:0] n39_O_2_2; // @[Top.scala 114:21]
  wire [15:0] n39_O_3_0; // @[Top.scala 114:21]
  wire [15:0] n39_O_3_1; // @[Top.scala 114:21]
  wire [15:0] n39_O_3_2; // @[Top.scala 114:21]
  wire  n48_valid_up; // @[Top.scala 118:21]
  wire  n48_valid_down; // @[Top.scala 118:21]
  wire [15:0] n48_I_0_0; // @[Top.scala 118:21]
  wire [15:0] n48_I_0_1; // @[Top.scala 118:21]
  wire [15:0] n48_I_0_2; // @[Top.scala 118:21]
  wire [15:0] n48_I_1_0; // @[Top.scala 118:21]
  wire [15:0] n48_I_1_1; // @[Top.scala 118:21]
  wire [15:0] n48_I_1_2; // @[Top.scala 118:21]
  wire [15:0] n48_I_2_0; // @[Top.scala 118:21]
  wire [15:0] n48_I_2_1; // @[Top.scala 118:21]
  wire [15:0] n48_I_2_2; // @[Top.scala 118:21]
  wire [15:0] n48_I_3_0; // @[Top.scala 118:21]
  wire [15:0] n48_I_3_1; // @[Top.scala 118:21]
  wire [15:0] n48_I_3_2; // @[Top.scala 118:21]
  wire [15:0] n48_O_0_0_0; // @[Top.scala 118:21]
  wire [15:0] n48_O_0_0_1; // @[Top.scala 118:21]
  wire [15:0] n48_O_0_0_2; // @[Top.scala 118:21]
  wire [15:0] n48_O_1_0_0; // @[Top.scala 118:21]
  wire [15:0] n48_O_1_0_1; // @[Top.scala 118:21]
  wire [15:0] n48_O_1_0_2; // @[Top.scala 118:21]
  wire [15:0] n48_O_2_0_0; // @[Top.scala 118:21]
  wire [15:0] n48_O_2_0_1; // @[Top.scala 118:21]
  wire [15:0] n48_O_2_0_2; // @[Top.scala 118:21]
  wire [15:0] n48_O_3_0_0; // @[Top.scala 118:21]
  wire [15:0] n48_O_3_0_1; // @[Top.scala 118:21]
  wire [15:0] n48_O_3_0_2; // @[Top.scala 118:21]
  wire  n55_valid_up; // @[Top.scala 121:21]
  wire  n55_valid_down; // @[Top.scala 121:21]
  wire [15:0] n55_I_0_0_0; // @[Top.scala 121:21]
  wire [15:0] n55_I_0_0_1; // @[Top.scala 121:21]
  wire [15:0] n55_I_0_0_2; // @[Top.scala 121:21]
  wire [15:0] n55_I_1_0_0; // @[Top.scala 121:21]
  wire [15:0] n55_I_1_0_1; // @[Top.scala 121:21]
  wire [15:0] n55_I_1_0_2; // @[Top.scala 121:21]
  wire [15:0] n55_I_2_0_0; // @[Top.scala 121:21]
  wire [15:0] n55_I_2_0_1; // @[Top.scala 121:21]
  wire [15:0] n55_I_2_0_2; // @[Top.scala 121:21]
  wire [15:0] n55_I_3_0_0; // @[Top.scala 121:21]
  wire [15:0] n55_I_3_0_1; // @[Top.scala 121:21]
  wire [15:0] n55_I_3_0_2; // @[Top.scala 121:21]
  wire [15:0] n55_O_0_0; // @[Top.scala 121:21]
  wire [15:0] n55_O_0_1; // @[Top.scala 121:21]
  wire [15:0] n55_O_0_2; // @[Top.scala 121:21]
  wire [15:0] n55_O_1_0; // @[Top.scala 121:21]
  wire [15:0] n55_O_1_1; // @[Top.scala 121:21]
  wire [15:0] n55_O_1_2; // @[Top.scala 121:21]
  wire [15:0] n55_O_2_0; // @[Top.scala 121:21]
  wire [15:0] n55_O_2_1; // @[Top.scala 121:21]
  wire [15:0] n55_O_2_2; // @[Top.scala 121:21]
  wire [15:0] n55_O_3_0; // @[Top.scala 121:21]
  wire [15:0] n55_O_3_1; // @[Top.scala 121:21]
  wire [15:0] n55_O_3_2; // @[Top.scala 121:21]
  wire  n56_valid_up; // @[Top.scala 124:21]
  wire  n56_valid_down; // @[Top.scala 124:21]
  wire [15:0] n56_I0_0_0; // @[Top.scala 124:21]
  wire [15:0] n56_I0_0_1; // @[Top.scala 124:21]
  wire [15:0] n56_I0_0_2; // @[Top.scala 124:21]
  wire [15:0] n56_I0_1_0; // @[Top.scala 124:21]
  wire [15:0] n56_I0_1_1; // @[Top.scala 124:21]
  wire [15:0] n56_I0_1_2; // @[Top.scala 124:21]
  wire [15:0] n56_I0_2_0; // @[Top.scala 124:21]
  wire [15:0] n56_I0_2_1; // @[Top.scala 124:21]
  wire [15:0] n56_I0_2_2; // @[Top.scala 124:21]
  wire [15:0] n56_I0_3_0; // @[Top.scala 124:21]
  wire [15:0] n56_I0_3_1; // @[Top.scala 124:21]
  wire [15:0] n56_I0_3_2; // @[Top.scala 124:21]
  wire [15:0] n56_I1_0_0; // @[Top.scala 124:21]
  wire [15:0] n56_I1_0_1; // @[Top.scala 124:21]
  wire [15:0] n56_I1_0_2; // @[Top.scala 124:21]
  wire [15:0] n56_I1_1_0; // @[Top.scala 124:21]
  wire [15:0] n56_I1_1_1; // @[Top.scala 124:21]
  wire [15:0] n56_I1_1_2; // @[Top.scala 124:21]
  wire [15:0] n56_I1_2_0; // @[Top.scala 124:21]
  wire [15:0] n56_I1_2_1; // @[Top.scala 124:21]
  wire [15:0] n56_I1_2_2; // @[Top.scala 124:21]
  wire [15:0] n56_I1_3_0; // @[Top.scala 124:21]
  wire [15:0] n56_I1_3_1; // @[Top.scala 124:21]
  wire [15:0] n56_I1_3_2; // @[Top.scala 124:21]
  wire [15:0] n56_O_0_0_0; // @[Top.scala 124:21]
  wire [15:0] n56_O_0_0_1; // @[Top.scala 124:21]
  wire [15:0] n56_O_0_0_2; // @[Top.scala 124:21]
  wire [15:0] n56_O_0_1_0; // @[Top.scala 124:21]
  wire [15:0] n56_O_0_1_1; // @[Top.scala 124:21]
  wire [15:0] n56_O_0_1_2; // @[Top.scala 124:21]
  wire [15:0] n56_O_1_0_0; // @[Top.scala 124:21]
  wire [15:0] n56_O_1_0_1; // @[Top.scala 124:21]
  wire [15:0] n56_O_1_0_2; // @[Top.scala 124:21]
  wire [15:0] n56_O_1_1_0; // @[Top.scala 124:21]
  wire [15:0] n56_O_1_1_1; // @[Top.scala 124:21]
  wire [15:0] n56_O_1_1_2; // @[Top.scala 124:21]
  wire [15:0] n56_O_2_0_0; // @[Top.scala 124:21]
  wire [15:0] n56_O_2_0_1; // @[Top.scala 124:21]
  wire [15:0] n56_O_2_0_2; // @[Top.scala 124:21]
  wire [15:0] n56_O_2_1_0; // @[Top.scala 124:21]
  wire [15:0] n56_O_2_1_1; // @[Top.scala 124:21]
  wire [15:0] n56_O_2_1_2; // @[Top.scala 124:21]
  wire [15:0] n56_O_3_0_0; // @[Top.scala 124:21]
  wire [15:0] n56_O_3_0_1; // @[Top.scala 124:21]
  wire [15:0] n56_O_3_0_2; // @[Top.scala 124:21]
  wire [15:0] n56_O_3_1_0; // @[Top.scala 124:21]
  wire [15:0] n56_O_3_1_1; // @[Top.scala 124:21]
  wire [15:0] n56_O_3_1_2; // @[Top.scala 124:21]
  wire  n63_clock; // @[Top.scala 128:21]
  wire  n63_valid_up; // @[Top.scala 128:21]
  wire  n63_valid_down; // @[Top.scala 128:21]
  wire [15:0] n63_I_0; // @[Top.scala 128:21]
  wire [15:0] n63_I_1; // @[Top.scala 128:21]
  wire [15:0] n63_I_2; // @[Top.scala 128:21]
  wire [15:0] n63_I_3; // @[Top.scala 128:21]
  wire [15:0] n63_O_0; // @[Top.scala 128:21]
  wire [15:0] n63_O_1; // @[Top.scala 128:21]
  wire [15:0] n63_O_2; // @[Top.scala 128:21]
  wire [15:0] n63_O_3; // @[Top.scala 128:21]
  wire  n64_clock; // @[Top.scala 131:21]
  wire  n64_valid_up; // @[Top.scala 131:21]
  wire  n64_valid_down; // @[Top.scala 131:21]
  wire [15:0] n64_I_0; // @[Top.scala 131:21]
  wire [15:0] n64_I_1; // @[Top.scala 131:21]
  wire [15:0] n64_I_2; // @[Top.scala 131:21]
  wire [15:0] n64_I_3; // @[Top.scala 131:21]
  wire [15:0] n64_O_0; // @[Top.scala 131:21]
  wire [15:0] n64_O_1; // @[Top.scala 131:21]
  wire [15:0] n64_O_2; // @[Top.scala 131:21]
  wire [15:0] n64_O_3; // @[Top.scala 131:21]
  wire  n65_valid_up; // @[Top.scala 134:21]
  wire  n65_valid_down; // @[Top.scala 134:21]
  wire [15:0] n65_I0_0; // @[Top.scala 134:21]
  wire [15:0] n65_I0_1; // @[Top.scala 134:21]
  wire [15:0] n65_I0_2; // @[Top.scala 134:21]
  wire [15:0] n65_I0_3; // @[Top.scala 134:21]
  wire [15:0] n65_I1_0; // @[Top.scala 134:21]
  wire [15:0] n65_I1_1; // @[Top.scala 134:21]
  wire [15:0] n65_I1_2; // @[Top.scala 134:21]
  wire [15:0] n65_I1_3; // @[Top.scala 134:21]
  wire [15:0] n65_O_0_0; // @[Top.scala 134:21]
  wire [15:0] n65_O_0_1; // @[Top.scala 134:21]
  wire [15:0] n65_O_1_0; // @[Top.scala 134:21]
  wire [15:0] n65_O_1_1; // @[Top.scala 134:21]
  wire [15:0] n65_O_2_0; // @[Top.scala 134:21]
  wire [15:0] n65_O_2_1; // @[Top.scala 134:21]
  wire [15:0] n65_O_3_0; // @[Top.scala 134:21]
  wire [15:0] n65_O_3_1; // @[Top.scala 134:21]
  wire  n72_valid_up; // @[Top.scala 138:21]
  wire  n72_valid_down; // @[Top.scala 138:21]
  wire [15:0] n72_I0_0_0; // @[Top.scala 138:21]
  wire [15:0] n72_I0_0_1; // @[Top.scala 138:21]
  wire [15:0] n72_I0_1_0; // @[Top.scala 138:21]
  wire [15:0] n72_I0_1_1; // @[Top.scala 138:21]
  wire [15:0] n72_I0_2_0; // @[Top.scala 138:21]
  wire [15:0] n72_I0_2_1; // @[Top.scala 138:21]
  wire [15:0] n72_I0_3_0; // @[Top.scala 138:21]
  wire [15:0] n72_I0_3_1; // @[Top.scala 138:21]
  wire [15:0] n72_I1_0; // @[Top.scala 138:21]
  wire [15:0] n72_I1_1; // @[Top.scala 138:21]
  wire [15:0] n72_I1_2; // @[Top.scala 138:21]
  wire [15:0] n72_I1_3; // @[Top.scala 138:21]
  wire [15:0] n72_O_0_0; // @[Top.scala 138:21]
  wire [15:0] n72_O_0_1; // @[Top.scala 138:21]
  wire [15:0] n72_O_0_2; // @[Top.scala 138:21]
  wire [15:0] n72_O_1_0; // @[Top.scala 138:21]
  wire [15:0] n72_O_1_1; // @[Top.scala 138:21]
  wire [15:0] n72_O_1_2; // @[Top.scala 138:21]
  wire [15:0] n72_O_2_0; // @[Top.scala 138:21]
  wire [15:0] n72_O_2_1; // @[Top.scala 138:21]
  wire [15:0] n72_O_2_2; // @[Top.scala 138:21]
  wire [15:0] n72_O_3_0; // @[Top.scala 138:21]
  wire [15:0] n72_O_3_1; // @[Top.scala 138:21]
  wire [15:0] n72_O_3_2; // @[Top.scala 138:21]
  wire  n81_valid_up; // @[Top.scala 142:21]
  wire  n81_valid_down; // @[Top.scala 142:21]
  wire [15:0] n81_I_0_0; // @[Top.scala 142:21]
  wire [15:0] n81_I_0_1; // @[Top.scala 142:21]
  wire [15:0] n81_I_0_2; // @[Top.scala 142:21]
  wire [15:0] n81_I_1_0; // @[Top.scala 142:21]
  wire [15:0] n81_I_1_1; // @[Top.scala 142:21]
  wire [15:0] n81_I_1_2; // @[Top.scala 142:21]
  wire [15:0] n81_I_2_0; // @[Top.scala 142:21]
  wire [15:0] n81_I_2_1; // @[Top.scala 142:21]
  wire [15:0] n81_I_2_2; // @[Top.scala 142:21]
  wire [15:0] n81_I_3_0; // @[Top.scala 142:21]
  wire [15:0] n81_I_3_1; // @[Top.scala 142:21]
  wire [15:0] n81_I_3_2; // @[Top.scala 142:21]
  wire [15:0] n81_O_0_0_0; // @[Top.scala 142:21]
  wire [15:0] n81_O_0_0_1; // @[Top.scala 142:21]
  wire [15:0] n81_O_0_0_2; // @[Top.scala 142:21]
  wire [15:0] n81_O_1_0_0; // @[Top.scala 142:21]
  wire [15:0] n81_O_1_0_1; // @[Top.scala 142:21]
  wire [15:0] n81_O_1_0_2; // @[Top.scala 142:21]
  wire [15:0] n81_O_2_0_0; // @[Top.scala 142:21]
  wire [15:0] n81_O_2_0_1; // @[Top.scala 142:21]
  wire [15:0] n81_O_2_0_2; // @[Top.scala 142:21]
  wire [15:0] n81_O_3_0_0; // @[Top.scala 142:21]
  wire [15:0] n81_O_3_0_1; // @[Top.scala 142:21]
  wire [15:0] n81_O_3_0_2; // @[Top.scala 142:21]
  wire  n88_valid_up; // @[Top.scala 145:21]
  wire  n88_valid_down; // @[Top.scala 145:21]
  wire [15:0] n88_I_0_0_0; // @[Top.scala 145:21]
  wire [15:0] n88_I_0_0_1; // @[Top.scala 145:21]
  wire [15:0] n88_I_0_0_2; // @[Top.scala 145:21]
  wire [15:0] n88_I_1_0_0; // @[Top.scala 145:21]
  wire [15:0] n88_I_1_0_1; // @[Top.scala 145:21]
  wire [15:0] n88_I_1_0_2; // @[Top.scala 145:21]
  wire [15:0] n88_I_2_0_0; // @[Top.scala 145:21]
  wire [15:0] n88_I_2_0_1; // @[Top.scala 145:21]
  wire [15:0] n88_I_2_0_2; // @[Top.scala 145:21]
  wire [15:0] n88_I_3_0_0; // @[Top.scala 145:21]
  wire [15:0] n88_I_3_0_1; // @[Top.scala 145:21]
  wire [15:0] n88_I_3_0_2; // @[Top.scala 145:21]
  wire [15:0] n88_O_0_0; // @[Top.scala 145:21]
  wire [15:0] n88_O_0_1; // @[Top.scala 145:21]
  wire [15:0] n88_O_0_2; // @[Top.scala 145:21]
  wire [15:0] n88_O_1_0; // @[Top.scala 145:21]
  wire [15:0] n88_O_1_1; // @[Top.scala 145:21]
  wire [15:0] n88_O_1_2; // @[Top.scala 145:21]
  wire [15:0] n88_O_2_0; // @[Top.scala 145:21]
  wire [15:0] n88_O_2_1; // @[Top.scala 145:21]
  wire [15:0] n88_O_2_2; // @[Top.scala 145:21]
  wire [15:0] n88_O_3_0; // @[Top.scala 145:21]
  wire [15:0] n88_O_3_1; // @[Top.scala 145:21]
  wire [15:0] n88_O_3_2; // @[Top.scala 145:21]
  wire  n89_valid_up; // @[Top.scala 148:21]
  wire  n89_valid_down; // @[Top.scala 148:21]
  wire [15:0] n89_I0_0_0_0; // @[Top.scala 148:21]
  wire [15:0] n89_I0_0_0_1; // @[Top.scala 148:21]
  wire [15:0] n89_I0_0_0_2; // @[Top.scala 148:21]
  wire [15:0] n89_I0_0_1_0; // @[Top.scala 148:21]
  wire [15:0] n89_I0_0_1_1; // @[Top.scala 148:21]
  wire [15:0] n89_I0_0_1_2; // @[Top.scala 148:21]
  wire [15:0] n89_I0_1_0_0; // @[Top.scala 148:21]
  wire [15:0] n89_I0_1_0_1; // @[Top.scala 148:21]
  wire [15:0] n89_I0_1_0_2; // @[Top.scala 148:21]
  wire [15:0] n89_I0_1_1_0; // @[Top.scala 148:21]
  wire [15:0] n89_I0_1_1_1; // @[Top.scala 148:21]
  wire [15:0] n89_I0_1_1_2; // @[Top.scala 148:21]
  wire [15:0] n89_I0_2_0_0; // @[Top.scala 148:21]
  wire [15:0] n89_I0_2_0_1; // @[Top.scala 148:21]
  wire [15:0] n89_I0_2_0_2; // @[Top.scala 148:21]
  wire [15:0] n89_I0_2_1_0; // @[Top.scala 148:21]
  wire [15:0] n89_I0_2_1_1; // @[Top.scala 148:21]
  wire [15:0] n89_I0_2_1_2; // @[Top.scala 148:21]
  wire [15:0] n89_I0_3_0_0; // @[Top.scala 148:21]
  wire [15:0] n89_I0_3_0_1; // @[Top.scala 148:21]
  wire [15:0] n89_I0_3_0_2; // @[Top.scala 148:21]
  wire [15:0] n89_I0_3_1_0; // @[Top.scala 148:21]
  wire [15:0] n89_I0_3_1_1; // @[Top.scala 148:21]
  wire [15:0] n89_I0_3_1_2; // @[Top.scala 148:21]
  wire [15:0] n89_I1_0_0; // @[Top.scala 148:21]
  wire [15:0] n89_I1_0_1; // @[Top.scala 148:21]
  wire [15:0] n89_I1_0_2; // @[Top.scala 148:21]
  wire [15:0] n89_I1_1_0; // @[Top.scala 148:21]
  wire [15:0] n89_I1_1_1; // @[Top.scala 148:21]
  wire [15:0] n89_I1_1_2; // @[Top.scala 148:21]
  wire [15:0] n89_I1_2_0; // @[Top.scala 148:21]
  wire [15:0] n89_I1_2_1; // @[Top.scala 148:21]
  wire [15:0] n89_I1_2_2; // @[Top.scala 148:21]
  wire [15:0] n89_I1_3_0; // @[Top.scala 148:21]
  wire [15:0] n89_I1_3_1; // @[Top.scala 148:21]
  wire [15:0] n89_I1_3_2; // @[Top.scala 148:21]
  wire [15:0] n89_O_0_0_0; // @[Top.scala 148:21]
  wire [15:0] n89_O_0_0_1; // @[Top.scala 148:21]
  wire [15:0] n89_O_0_0_2; // @[Top.scala 148:21]
  wire [15:0] n89_O_0_1_0; // @[Top.scala 148:21]
  wire [15:0] n89_O_0_1_1; // @[Top.scala 148:21]
  wire [15:0] n89_O_0_1_2; // @[Top.scala 148:21]
  wire [15:0] n89_O_0_2_0; // @[Top.scala 148:21]
  wire [15:0] n89_O_0_2_1; // @[Top.scala 148:21]
  wire [15:0] n89_O_0_2_2; // @[Top.scala 148:21]
  wire [15:0] n89_O_1_0_0; // @[Top.scala 148:21]
  wire [15:0] n89_O_1_0_1; // @[Top.scala 148:21]
  wire [15:0] n89_O_1_0_2; // @[Top.scala 148:21]
  wire [15:0] n89_O_1_1_0; // @[Top.scala 148:21]
  wire [15:0] n89_O_1_1_1; // @[Top.scala 148:21]
  wire [15:0] n89_O_1_1_2; // @[Top.scala 148:21]
  wire [15:0] n89_O_1_2_0; // @[Top.scala 148:21]
  wire [15:0] n89_O_1_2_1; // @[Top.scala 148:21]
  wire [15:0] n89_O_1_2_2; // @[Top.scala 148:21]
  wire [15:0] n89_O_2_0_0; // @[Top.scala 148:21]
  wire [15:0] n89_O_2_0_1; // @[Top.scala 148:21]
  wire [15:0] n89_O_2_0_2; // @[Top.scala 148:21]
  wire [15:0] n89_O_2_1_0; // @[Top.scala 148:21]
  wire [15:0] n89_O_2_1_1; // @[Top.scala 148:21]
  wire [15:0] n89_O_2_1_2; // @[Top.scala 148:21]
  wire [15:0] n89_O_2_2_0; // @[Top.scala 148:21]
  wire [15:0] n89_O_2_2_1; // @[Top.scala 148:21]
  wire [15:0] n89_O_2_2_2; // @[Top.scala 148:21]
  wire [15:0] n89_O_3_0_0; // @[Top.scala 148:21]
  wire [15:0] n89_O_3_0_1; // @[Top.scala 148:21]
  wire [15:0] n89_O_3_0_2; // @[Top.scala 148:21]
  wire [15:0] n89_O_3_1_0; // @[Top.scala 148:21]
  wire [15:0] n89_O_3_1_1; // @[Top.scala 148:21]
  wire [15:0] n89_O_3_1_2; // @[Top.scala 148:21]
  wire [15:0] n89_O_3_2_0; // @[Top.scala 148:21]
  wire [15:0] n89_O_3_2_1; // @[Top.scala 148:21]
  wire [15:0] n89_O_3_2_2; // @[Top.scala 148:21]
  wire  n98_valid_up; // @[Top.scala 152:21]
  wire  n98_valid_down; // @[Top.scala 152:21]
  wire [15:0] n98_I_0_0_0; // @[Top.scala 152:21]
  wire [15:0] n98_I_0_0_1; // @[Top.scala 152:21]
  wire [15:0] n98_I_0_0_2; // @[Top.scala 152:21]
  wire [15:0] n98_I_0_1_0; // @[Top.scala 152:21]
  wire [15:0] n98_I_0_1_1; // @[Top.scala 152:21]
  wire [15:0] n98_I_0_1_2; // @[Top.scala 152:21]
  wire [15:0] n98_I_0_2_0; // @[Top.scala 152:21]
  wire [15:0] n98_I_0_2_1; // @[Top.scala 152:21]
  wire [15:0] n98_I_0_2_2; // @[Top.scala 152:21]
  wire [15:0] n98_I_1_0_0; // @[Top.scala 152:21]
  wire [15:0] n98_I_1_0_1; // @[Top.scala 152:21]
  wire [15:0] n98_I_1_0_2; // @[Top.scala 152:21]
  wire [15:0] n98_I_1_1_0; // @[Top.scala 152:21]
  wire [15:0] n98_I_1_1_1; // @[Top.scala 152:21]
  wire [15:0] n98_I_1_1_2; // @[Top.scala 152:21]
  wire [15:0] n98_I_1_2_0; // @[Top.scala 152:21]
  wire [15:0] n98_I_1_2_1; // @[Top.scala 152:21]
  wire [15:0] n98_I_1_2_2; // @[Top.scala 152:21]
  wire [15:0] n98_I_2_0_0; // @[Top.scala 152:21]
  wire [15:0] n98_I_2_0_1; // @[Top.scala 152:21]
  wire [15:0] n98_I_2_0_2; // @[Top.scala 152:21]
  wire [15:0] n98_I_2_1_0; // @[Top.scala 152:21]
  wire [15:0] n98_I_2_1_1; // @[Top.scala 152:21]
  wire [15:0] n98_I_2_1_2; // @[Top.scala 152:21]
  wire [15:0] n98_I_2_2_0; // @[Top.scala 152:21]
  wire [15:0] n98_I_2_2_1; // @[Top.scala 152:21]
  wire [15:0] n98_I_2_2_2; // @[Top.scala 152:21]
  wire [15:0] n98_I_3_0_0; // @[Top.scala 152:21]
  wire [15:0] n98_I_3_0_1; // @[Top.scala 152:21]
  wire [15:0] n98_I_3_0_2; // @[Top.scala 152:21]
  wire [15:0] n98_I_3_1_0; // @[Top.scala 152:21]
  wire [15:0] n98_I_3_1_1; // @[Top.scala 152:21]
  wire [15:0] n98_I_3_1_2; // @[Top.scala 152:21]
  wire [15:0] n98_I_3_2_0; // @[Top.scala 152:21]
  wire [15:0] n98_I_3_2_1; // @[Top.scala 152:21]
  wire [15:0] n98_I_3_2_2; // @[Top.scala 152:21]
  wire [15:0] n98_O_0_0_0_0; // @[Top.scala 152:21]
  wire [15:0] n98_O_0_0_0_1; // @[Top.scala 152:21]
  wire [15:0] n98_O_0_0_0_2; // @[Top.scala 152:21]
  wire [15:0] n98_O_0_0_1_0; // @[Top.scala 152:21]
  wire [15:0] n98_O_0_0_1_1; // @[Top.scala 152:21]
  wire [15:0] n98_O_0_0_1_2; // @[Top.scala 152:21]
  wire [15:0] n98_O_0_0_2_0; // @[Top.scala 152:21]
  wire [15:0] n98_O_0_0_2_1; // @[Top.scala 152:21]
  wire [15:0] n98_O_0_0_2_2; // @[Top.scala 152:21]
  wire [15:0] n98_O_1_0_0_0; // @[Top.scala 152:21]
  wire [15:0] n98_O_1_0_0_1; // @[Top.scala 152:21]
  wire [15:0] n98_O_1_0_0_2; // @[Top.scala 152:21]
  wire [15:0] n98_O_1_0_1_0; // @[Top.scala 152:21]
  wire [15:0] n98_O_1_0_1_1; // @[Top.scala 152:21]
  wire [15:0] n98_O_1_0_1_2; // @[Top.scala 152:21]
  wire [15:0] n98_O_1_0_2_0; // @[Top.scala 152:21]
  wire [15:0] n98_O_1_0_2_1; // @[Top.scala 152:21]
  wire [15:0] n98_O_1_0_2_2; // @[Top.scala 152:21]
  wire [15:0] n98_O_2_0_0_0; // @[Top.scala 152:21]
  wire [15:0] n98_O_2_0_0_1; // @[Top.scala 152:21]
  wire [15:0] n98_O_2_0_0_2; // @[Top.scala 152:21]
  wire [15:0] n98_O_2_0_1_0; // @[Top.scala 152:21]
  wire [15:0] n98_O_2_0_1_1; // @[Top.scala 152:21]
  wire [15:0] n98_O_2_0_1_2; // @[Top.scala 152:21]
  wire [15:0] n98_O_2_0_2_0; // @[Top.scala 152:21]
  wire [15:0] n98_O_2_0_2_1; // @[Top.scala 152:21]
  wire [15:0] n98_O_2_0_2_2; // @[Top.scala 152:21]
  wire [15:0] n98_O_3_0_0_0; // @[Top.scala 152:21]
  wire [15:0] n98_O_3_0_0_1; // @[Top.scala 152:21]
  wire [15:0] n98_O_3_0_0_2; // @[Top.scala 152:21]
  wire [15:0] n98_O_3_0_1_0; // @[Top.scala 152:21]
  wire [15:0] n98_O_3_0_1_1; // @[Top.scala 152:21]
  wire [15:0] n98_O_3_0_1_2; // @[Top.scala 152:21]
  wire [15:0] n98_O_3_0_2_0; // @[Top.scala 152:21]
  wire [15:0] n98_O_3_0_2_1; // @[Top.scala 152:21]
  wire [15:0] n98_O_3_0_2_2; // @[Top.scala 152:21]
  wire  n105_valid_up; // @[Top.scala 155:22]
  wire  n105_valid_down; // @[Top.scala 155:22]
  wire [15:0] n105_I_0_0_0_0; // @[Top.scala 155:22]
  wire [15:0] n105_I_0_0_0_1; // @[Top.scala 155:22]
  wire [15:0] n105_I_0_0_0_2; // @[Top.scala 155:22]
  wire [15:0] n105_I_0_0_1_0; // @[Top.scala 155:22]
  wire [15:0] n105_I_0_0_1_1; // @[Top.scala 155:22]
  wire [15:0] n105_I_0_0_1_2; // @[Top.scala 155:22]
  wire [15:0] n105_I_0_0_2_0; // @[Top.scala 155:22]
  wire [15:0] n105_I_0_0_2_1; // @[Top.scala 155:22]
  wire [15:0] n105_I_0_0_2_2; // @[Top.scala 155:22]
  wire [15:0] n105_I_1_0_0_0; // @[Top.scala 155:22]
  wire [15:0] n105_I_1_0_0_1; // @[Top.scala 155:22]
  wire [15:0] n105_I_1_0_0_2; // @[Top.scala 155:22]
  wire [15:0] n105_I_1_0_1_0; // @[Top.scala 155:22]
  wire [15:0] n105_I_1_0_1_1; // @[Top.scala 155:22]
  wire [15:0] n105_I_1_0_1_2; // @[Top.scala 155:22]
  wire [15:0] n105_I_1_0_2_0; // @[Top.scala 155:22]
  wire [15:0] n105_I_1_0_2_1; // @[Top.scala 155:22]
  wire [15:0] n105_I_1_0_2_2; // @[Top.scala 155:22]
  wire [15:0] n105_I_2_0_0_0; // @[Top.scala 155:22]
  wire [15:0] n105_I_2_0_0_1; // @[Top.scala 155:22]
  wire [15:0] n105_I_2_0_0_2; // @[Top.scala 155:22]
  wire [15:0] n105_I_2_0_1_0; // @[Top.scala 155:22]
  wire [15:0] n105_I_2_0_1_1; // @[Top.scala 155:22]
  wire [15:0] n105_I_2_0_1_2; // @[Top.scala 155:22]
  wire [15:0] n105_I_2_0_2_0; // @[Top.scala 155:22]
  wire [15:0] n105_I_2_0_2_1; // @[Top.scala 155:22]
  wire [15:0] n105_I_2_0_2_2; // @[Top.scala 155:22]
  wire [15:0] n105_I_3_0_0_0; // @[Top.scala 155:22]
  wire [15:0] n105_I_3_0_0_1; // @[Top.scala 155:22]
  wire [15:0] n105_I_3_0_0_2; // @[Top.scala 155:22]
  wire [15:0] n105_I_3_0_1_0; // @[Top.scala 155:22]
  wire [15:0] n105_I_3_0_1_1; // @[Top.scala 155:22]
  wire [15:0] n105_I_3_0_1_2; // @[Top.scala 155:22]
  wire [15:0] n105_I_3_0_2_0; // @[Top.scala 155:22]
  wire [15:0] n105_I_3_0_2_1; // @[Top.scala 155:22]
  wire [15:0] n105_I_3_0_2_2; // @[Top.scala 155:22]
  wire [15:0] n105_O_0_0_0; // @[Top.scala 155:22]
  wire [15:0] n105_O_0_0_1; // @[Top.scala 155:22]
  wire [15:0] n105_O_0_0_2; // @[Top.scala 155:22]
  wire [15:0] n105_O_0_1_0; // @[Top.scala 155:22]
  wire [15:0] n105_O_0_1_1; // @[Top.scala 155:22]
  wire [15:0] n105_O_0_1_2; // @[Top.scala 155:22]
  wire [15:0] n105_O_0_2_0; // @[Top.scala 155:22]
  wire [15:0] n105_O_0_2_1; // @[Top.scala 155:22]
  wire [15:0] n105_O_0_2_2; // @[Top.scala 155:22]
  wire [15:0] n105_O_1_0_0; // @[Top.scala 155:22]
  wire [15:0] n105_O_1_0_1; // @[Top.scala 155:22]
  wire [15:0] n105_O_1_0_2; // @[Top.scala 155:22]
  wire [15:0] n105_O_1_1_0; // @[Top.scala 155:22]
  wire [15:0] n105_O_1_1_1; // @[Top.scala 155:22]
  wire [15:0] n105_O_1_1_2; // @[Top.scala 155:22]
  wire [15:0] n105_O_1_2_0; // @[Top.scala 155:22]
  wire [15:0] n105_O_1_2_1; // @[Top.scala 155:22]
  wire [15:0] n105_O_1_2_2; // @[Top.scala 155:22]
  wire [15:0] n105_O_2_0_0; // @[Top.scala 155:22]
  wire [15:0] n105_O_2_0_1; // @[Top.scala 155:22]
  wire [15:0] n105_O_2_0_2; // @[Top.scala 155:22]
  wire [15:0] n105_O_2_1_0; // @[Top.scala 155:22]
  wire [15:0] n105_O_2_1_1; // @[Top.scala 155:22]
  wire [15:0] n105_O_2_1_2; // @[Top.scala 155:22]
  wire [15:0] n105_O_2_2_0; // @[Top.scala 155:22]
  wire [15:0] n105_O_2_2_1; // @[Top.scala 155:22]
  wire [15:0] n105_O_2_2_2; // @[Top.scala 155:22]
  wire [15:0] n105_O_3_0_0; // @[Top.scala 155:22]
  wire [15:0] n105_O_3_0_1; // @[Top.scala 155:22]
  wire [15:0] n105_O_3_0_2; // @[Top.scala 155:22]
  wire [15:0] n105_O_3_1_0; // @[Top.scala 155:22]
  wire [15:0] n105_O_3_1_1; // @[Top.scala 155:22]
  wire [15:0] n105_O_3_1_2; // @[Top.scala 155:22]
  wire [15:0] n105_O_3_2_0; // @[Top.scala 155:22]
  wire [15:0] n105_O_3_2_1; // @[Top.scala 155:22]
  wire [15:0] n105_O_3_2_2; // @[Top.scala 155:22]
  wire  n147_clock; // @[Top.scala 158:22]
  wire  n147_reset; // @[Top.scala 158:22]
  wire  n147_valid_up; // @[Top.scala 158:22]
  wire  n147_valid_down; // @[Top.scala 158:22]
  wire [15:0] n147_I_0_0_0; // @[Top.scala 158:22]
  wire [15:0] n147_I_0_0_1; // @[Top.scala 158:22]
  wire [15:0] n147_I_0_0_2; // @[Top.scala 158:22]
  wire [15:0] n147_I_0_1_0; // @[Top.scala 158:22]
  wire [15:0] n147_I_0_1_1; // @[Top.scala 158:22]
  wire [15:0] n147_I_0_1_2; // @[Top.scala 158:22]
  wire [15:0] n147_I_0_2_0; // @[Top.scala 158:22]
  wire [15:0] n147_I_0_2_1; // @[Top.scala 158:22]
  wire [15:0] n147_I_0_2_2; // @[Top.scala 158:22]
  wire [15:0] n147_I_1_0_0; // @[Top.scala 158:22]
  wire [15:0] n147_I_1_0_1; // @[Top.scala 158:22]
  wire [15:0] n147_I_1_0_2; // @[Top.scala 158:22]
  wire [15:0] n147_I_1_1_0; // @[Top.scala 158:22]
  wire [15:0] n147_I_1_1_1; // @[Top.scala 158:22]
  wire [15:0] n147_I_1_1_2; // @[Top.scala 158:22]
  wire [15:0] n147_I_1_2_0; // @[Top.scala 158:22]
  wire [15:0] n147_I_1_2_1; // @[Top.scala 158:22]
  wire [15:0] n147_I_1_2_2; // @[Top.scala 158:22]
  wire [15:0] n147_I_2_0_0; // @[Top.scala 158:22]
  wire [15:0] n147_I_2_0_1; // @[Top.scala 158:22]
  wire [15:0] n147_I_2_0_2; // @[Top.scala 158:22]
  wire [15:0] n147_I_2_1_0; // @[Top.scala 158:22]
  wire [15:0] n147_I_2_1_1; // @[Top.scala 158:22]
  wire [15:0] n147_I_2_1_2; // @[Top.scala 158:22]
  wire [15:0] n147_I_2_2_0; // @[Top.scala 158:22]
  wire [15:0] n147_I_2_2_1; // @[Top.scala 158:22]
  wire [15:0] n147_I_2_2_2; // @[Top.scala 158:22]
  wire [15:0] n147_I_3_0_0; // @[Top.scala 158:22]
  wire [15:0] n147_I_3_0_1; // @[Top.scala 158:22]
  wire [15:0] n147_I_3_0_2; // @[Top.scala 158:22]
  wire [15:0] n147_I_3_1_0; // @[Top.scala 158:22]
  wire [15:0] n147_I_3_1_1; // @[Top.scala 158:22]
  wire [15:0] n147_I_3_1_2; // @[Top.scala 158:22]
  wire [15:0] n147_I_3_2_0; // @[Top.scala 158:22]
  wire [15:0] n147_I_3_2_1; // @[Top.scala 158:22]
  wire [15:0] n147_I_3_2_2; // @[Top.scala 158:22]
  wire [15:0] n147_O_0_0_0; // @[Top.scala 158:22]
  wire [15:0] n147_O_1_0_0; // @[Top.scala 158:22]
  wire [15:0] n147_O_2_0_0; // @[Top.scala 158:22]
  wire [15:0] n147_O_3_0_0; // @[Top.scala 158:22]
  wire  n148_valid_up; // @[Top.scala 161:22]
  wire  n148_valid_down; // @[Top.scala 161:22]
  wire [15:0] n148_I_0_0_0; // @[Top.scala 161:22]
  wire [15:0] n148_I_1_0_0; // @[Top.scala 161:22]
  wire [15:0] n148_I_2_0_0; // @[Top.scala 161:22]
  wire [15:0] n148_I_3_0_0; // @[Top.scala 161:22]
  wire [15:0] n148_O_0_0; // @[Top.scala 161:22]
  wire [15:0] n148_O_1_0; // @[Top.scala 161:22]
  wire [15:0] n148_O_2_0; // @[Top.scala 161:22]
  wire [15:0] n148_O_3_0; // @[Top.scala 161:22]
  wire  n149_valid_up; // @[Top.scala 164:22]
  wire  n149_valid_down; // @[Top.scala 164:22]
  wire [15:0] n149_I_0_0; // @[Top.scala 164:22]
  wire [15:0] n149_I_1_0; // @[Top.scala 164:22]
  wire [15:0] n149_I_2_0; // @[Top.scala 164:22]
  wire [15:0] n149_I_3_0; // @[Top.scala 164:22]
  wire [15:0] n149_O_0; // @[Top.scala 164:22]
  wire [15:0] n149_O_1; // @[Top.scala 164:22]
  wire [15:0] n149_O_2; // @[Top.scala 164:22]
  wire [15:0] n149_O_3; // @[Top.scala 164:22]
  wire  n150_clock; // @[Top.scala 167:22]
  wire  n150_reset; // @[Top.scala 167:22]
  wire  n150_valid_up; // @[Top.scala 167:22]
  wire  n150_valid_down; // @[Top.scala 167:22]
  wire [15:0] n150_I_0; // @[Top.scala 167:22]
  wire [15:0] n150_I_1; // @[Top.scala 167:22]
  wire [15:0] n150_I_2; // @[Top.scala 167:22]
  wire [15:0] n150_I_3; // @[Top.scala 167:22]
  wire [15:0] n150_O_0; // @[Top.scala 167:22]
  wire [15:0] n150_O_1; // @[Top.scala 167:22]
  wire [15:0] n150_O_2; // @[Top.scala 167:22]
  wire [15:0] n150_O_3; // @[Top.scala 167:22]
  wire  n151_clock; // @[Top.scala 170:22]
  wire  n151_valid_up; // @[Top.scala 170:22]
  wire  n151_valid_down; // @[Top.scala 170:22]
  wire [15:0] n151_I_0; // @[Top.scala 170:22]
  wire [15:0] n151_I_1; // @[Top.scala 170:22]
  wire [15:0] n151_I_2; // @[Top.scala 170:22]
  wire [15:0] n151_I_3; // @[Top.scala 170:22]
  wire [15:0] n151_O_0; // @[Top.scala 170:22]
  wire [15:0] n151_O_1; // @[Top.scala 170:22]
  wire [15:0] n151_O_2; // @[Top.scala 170:22]
  wire [15:0] n151_O_3; // @[Top.scala 170:22]
  wire  n152_valid_up; // @[Top.scala 173:22]
  wire  n152_valid_down; // @[Top.scala 173:22]
  wire [15:0] n152_I0_0; // @[Top.scala 173:22]
  wire [15:0] n152_I0_1; // @[Top.scala 173:22]
  wire [15:0] n152_I0_2; // @[Top.scala 173:22]
  wire [15:0] n152_I0_3; // @[Top.scala 173:22]
  wire [15:0] n152_I1_0; // @[Top.scala 173:22]
  wire [15:0] n152_I1_1; // @[Top.scala 173:22]
  wire [15:0] n152_I1_2; // @[Top.scala 173:22]
  wire [15:0] n152_I1_3; // @[Top.scala 173:22]
  wire [15:0] n152_O_0_0; // @[Top.scala 173:22]
  wire [15:0] n152_O_0_1; // @[Top.scala 173:22]
  wire [15:0] n152_O_1_0; // @[Top.scala 173:22]
  wire [15:0] n152_O_1_1; // @[Top.scala 173:22]
  wire [15:0] n152_O_2_0; // @[Top.scala 173:22]
  wire [15:0] n152_O_2_1; // @[Top.scala 173:22]
  wire [15:0] n152_O_3_0; // @[Top.scala 173:22]
  wire [15:0] n152_O_3_1; // @[Top.scala 173:22]
  wire  n161_valid_up; // @[Top.scala 177:22]
  wire  n161_valid_down; // @[Top.scala 177:22]
  wire [15:0] n161_I_0_0; // @[Top.scala 177:22]
  wire [15:0] n161_I_0_1; // @[Top.scala 177:22]
  wire [15:0] n161_I_1_0; // @[Top.scala 177:22]
  wire [15:0] n161_I_1_1; // @[Top.scala 177:22]
  wire [15:0] n161_I_2_0; // @[Top.scala 177:22]
  wire [15:0] n161_I_2_1; // @[Top.scala 177:22]
  wire [15:0] n161_I_3_0; // @[Top.scala 177:22]
  wire [15:0] n161_I_3_1; // @[Top.scala 177:22]
  wire [15:0] n161_O_0_0_0; // @[Top.scala 177:22]
  wire [15:0] n161_O_0_0_1; // @[Top.scala 177:22]
  wire [15:0] n161_O_1_0_0; // @[Top.scala 177:22]
  wire [15:0] n161_O_1_0_1; // @[Top.scala 177:22]
  wire [15:0] n161_O_2_0_0; // @[Top.scala 177:22]
  wire [15:0] n161_O_2_0_1; // @[Top.scala 177:22]
  wire [15:0] n161_O_3_0_0; // @[Top.scala 177:22]
  wire [15:0] n161_O_3_0_1; // @[Top.scala 177:22]
  wire  n168_valid_up; // @[Top.scala 180:22]
  wire  n168_valid_down; // @[Top.scala 180:22]
  wire [15:0] n168_I_0_0_0; // @[Top.scala 180:22]
  wire [15:0] n168_I_0_0_1; // @[Top.scala 180:22]
  wire [15:0] n168_I_1_0_0; // @[Top.scala 180:22]
  wire [15:0] n168_I_1_0_1; // @[Top.scala 180:22]
  wire [15:0] n168_I_2_0_0; // @[Top.scala 180:22]
  wire [15:0] n168_I_2_0_1; // @[Top.scala 180:22]
  wire [15:0] n168_I_3_0_0; // @[Top.scala 180:22]
  wire [15:0] n168_I_3_0_1; // @[Top.scala 180:22]
  wire [15:0] n168_O_0_0; // @[Top.scala 180:22]
  wire [15:0] n168_O_0_1; // @[Top.scala 180:22]
  wire [15:0] n168_O_1_0; // @[Top.scala 180:22]
  wire [15:0] n168_O_1_1; // @[Top.scala 180:22]
  wire [15:0] n168_O_2_0; // @[Top.scala 180:22]
  wire [15:0] n168_O_2_1; // @[Top.scala 180:22]
  wire [15:0] n168_O_3_0; // @[Top.scala 180:22]
  wire [15:0] n168_O_3_1; // @[Top.scala 180:22]
  wire  n169_clock; // @[Top.scala 183:22]
  wire  n169_valid_up; // @[Top.scala 183:22]
  wire  n169_valid_down; // @[Top.scala 183:22]
  wire [15:0] n169_I_0; // @[Top.scala 183:22]
  wire [15:0] n169_I_1; // @[Top.scala 183:22]
  wire [15:0] n169_I_2; // @[Top.scala 183:22]
  wire [15:0] n169_I_3; // @[Top.scala 183:22]
  wire [15:0] n169_O_0; // @[Top.scala 183:22]
  wire [15:0] n169_O_1; // @[Top.scala 183:22]
  wire [15:0] n169_O_2; // @[Top.scala 183:22]
  wire [15:0] n169_O_3; // @[Top.scala 183:22]
  wire  n170_valid_up; // @[Top.scala 186:22]
  wire  n170_valid_down; // @[Top.scala 186:22]
  wire [15:0] n170_I0_0; // @[Top.scala 186:22]
  wire [15:0] n170_I0_1; // @[Top.scala 186:22]
  wire [15:0] n170_I0_2; // @[Top.scala 186:22]
  wire [15:0] n170_I0_3; // @[Top.scala 186:22]
  wire [15:0] n170_I1_0; // @[Top.scala 186:22]
  wire [15:0] n170_I1_1; // @[Top.scala 186:22]
  wire [15:0] n170_I1_2; // @[Top.scala 186:22]
  wire [15:0] n170_I1_3; // @[Top.scala 186:22]
  wire [15:0] n170_O_0_0; // @[Top.scala 186:22]
  wire [15:0] n170_O_0_1; // @[Top.scala 186:22]
  wire [15:0] n170_O_1_0; // @[Top.scala 186:22]
  wire [15:0] n170_O_1_1; // @[Top.scala 186:22]
  wire [15:0] n170_O_2_0; // @[Top.scala 186:22]
  wire [15:0] n170_O_2_1; // @[Top.scala 186:22]
  wire [15:0] n170_O_3_0; // @[Top.scala 186:22]
  wire [15:0] n170_O_3_1; // @[Top.scala 186:22]
  wire  n179_valid_up; // @[Top.scala 190:22]
  wire  n179_valid_down; // @[Top.scala 190:22]
  wire [15:0] n179_I_0_0; // @[Top.scala 190:22]
  wire [15:0] n179_I_0_1; // @[Top.scala 190:22]
  wire [15:0] n179_I_1_0; // @[Top.scala 190:22]
  wire [15:0] n179_I_1_1; // @[Top.scala 190:22]
  wire [15:0] n179_I_2_0; // @[Top.scala 190:22]
  wire [15:0] n179_I_2_1; // @[Top.scala 190:22]
  wire [15:0] n179_I_3_0; // @[Top.scala 190:22]
  wire [15:0] n179_I_3_1; // @[Top.scala 190:22]
  wire [15:0] n179_O_0_0_0; // @[Top.scala 190:22]
  wire [15:0] n179_O_0_0_1; // @[Top.scala 190:22]
  wire [15:0] n179_O_1_0_0; // @[Top.scala 190:22]
  wire [15:0] n179_O_1_0_1; // @[Top.scala 190:22]
  wire [15:0] n179_O_2_0_0; // @[Top.scala 190:22]
  wire [15:0] n179_O_2_0_1; // @[Top.scala 190:22]
  wire [15:0] n179_O_3_0_0; // @[Top.scala 190:22]
  wire [15:0] n179_O_3_0_1; // @[Top.scala 190:22]
  wire  n186_valid_up; // @[Top.scala 193:22]
  wire  n186_valid_down; // @[Top.scala 193:22]
  wire [15:0] n186_I_0_0_0; // @[Top.scala 193:22]
  wire [15:0] n186_I_0_0_1; // @[Top.scala 193:22]
  wire [15:0] n186_I_1_0_0; // @[Top.scala 193:22]
  wire [15:0] n186_I_1_0_1; // @[Top.scala 193:22]
  wire [15:0] n186_I_2_0_0; // @[Top.scala 193:22]
  wire [15:0] n186_I_2_0_1; // @[Top.scala 193:22]
  wire [15:0] n186_I_3_0_0; // @[Top.scala 193:22]
  wire [15:0] n186_I_3_0_1; // @[Top.scala 193:22]
  wire [15:0] n186_O_0_0; // @[Top.scala 193:22]
  wire [15:0] n186_O_0_1; // @[Top.scala 193:22]
  wire [15:0] n186_O_1_0; // @[Top.scala 193:22]
  wire [15:0] n186_O_1_1; // @[Top.scala 193:22]
  wire [15:0] n186_O_2_0; // @[Top.scala 193:22]
  wire [15:0] n186_O_2_1; // @[Top.scala 193:22]
  wire [15:0] n186_O_3_0; // @[Top.scala 193:22]
  wire [15:0] n186_O_3_1; // @[Top.scala 193:22]
  wire  n187_valid_up; // @[Top.scala 196:22]
  wire  n187_valid_down; // @[Top.scala 196:22]
  wire [15:0] n187_I0_0_0; // @[Top.scala 196:22]
  wire [15:0] n187_I0_0_1; // @[Top.scala 196:22]
  wire [15:0] n187_I0_1_0; // @[Top.scala 196:22]
  wire [15:0] n187_I0_1_1; // @[Top.scala 196:22]
  wire [15:0] n187_I0_2_0; // @[Top.scala 196:22]
  wire [15:0] n187_I0_2_1; // @[Top.scala 196:22]
  wire [15:0] n187_I0_3_0; // @[Top.scala 196:22]
  wire [15:0] n187_I0_3_1; // @[Top.scala 196:22]
  wire [15:0] n187_I1_0_0; // @[Top.scala 196:22]
  wire [15:0] n187_I1_0_1; // @[Top.scala 196:22]
  wire [15:0] n187_I1_1_0; // @[Top.scala 196:22]
  wire [15:0] n187_I1_1_1; // @[Top.scala 196:22]
  wire [15:0] n187_I1_2_0; // @[Top.scala 196:22]
  wire [15:0] n187_I1_2_1; // @[Top.scala 196:22]
  wire [15:0] n187_I1_3_0; // @[Top.scala 196:22]
  wire [15:0] n187_I1_3_1; // @[Top.scala 196:22]
  wire [15:0] n187_O_0_0_0; // @[Top.scala 196:22]
  wire [15:0] n187_O_0_0_1; // @[Top.scala 196:22]
  wire [15:0] n187_O_0_1_0; // @[Top.scala 196:22]
  wire [15:0] n187_O_0_1_1; // @[Top.scala 196:22]
  wire [15:0] n187_O_1_0_0; // @[Top.scala 196:22]
  wire [15:0] n187_O_1_0_1; // @[Top.scala 196:22]
  wire [15:0] n187_O_1_1_0; // @[Top.scala 196:22]
  wire [15:0] n187_O_1_1_1; // @[Top.scala 196:22]
  wire [15:0] n187_O_2_0_0; // @[Top.scala 196:22]
  wire [15:0] n187_O_2_0_1; // @[Top.scala 196:22]
  wire [15:0] n187_O_2_1_0; // @[Top.scala 196:22]
  wire [15:0] n187_O_2_1_1; // @[Top.scala 196:22]
  wire [15:0] n187_O_3_0_0; // @[Top.scala 196:22]
  wire [15:0] n187_O_3_0_1; // @[Top.scala 196:22]
  wire [15:0] n187_O_3_1_0; // @[Top.scala 196:22]
  wire [15:0] n187_O_3_1_1; // @[Top.scala 196:22]
  wire  n196_valid_up; // @[Top.scala 200:22]
  wire  n196_valid_down; // @[Top.scala 200:22]
  wire [15:0] n196_I_0_0_0; // @[Top.scala 200:22]
  wire [15:0] n196_I_0_0_1; // @[Top.scala 200:22]
  wire [15:0] n196_I_0_1_0; // @[Top.scala 200:22]
  wire [15:0] n196_I_0_1_1; // @[Top.scala 200:22]
  wire [15:0] n196_I_1_0_0; // @[Top.scala 200:22]
  wire [15:0] n196_I_1_0_1; // @[Top.scala 200:22]
  wire [15:0] n196_I_1_1_0; // @[Top.scala 200:22]
  wire [15:0] n196_I_1_1_1; // @[Top.scala 200:22]
  wire [15:0] n196_I_2_0_0; // @[Top.scala 200:22]
  wire [15:0] n196_I_2_0_1; // @[Top.scala 200:22]
  wire [15:0] n196_I_2_1_0; // @[Top.scala 200:22]
  wire [15:0] n196_I_2_1_1; // @[Top.scala 200:22]
  wire [15:0] n196_I_3_0_0; // @[Top.scala 200:22]
  wire [15:0] n196_I_3_0_1; // @[Top.scala 200:22]
  wire [15:0] n196_I_3_1_0; // @[Top.scala 200:22]
  wire [15:0] n196_I_3_1_1; // @[Top.scala 200:22]
  wire [15:0] n196_O_0_0_0_0; // @[Top.scala 200:22]
  wire [15:0] n196_O_0_0_0_1; // @[Top.scala 200:22]
  wire [15:0] n196_O_0_0_1_0; // @[Top.scala 200:22]
  wire [15:0] n196_O_0_0_1_1; // @[Top.scala 200:22]
  wire [15:0] n196_O_1_0_0_0; // @[Top.scala 200:22]
  wire [15:0] n196_O_1_0_0_1; // @[Top.scala 200:22]
  wire [15:0] n196_O_1_0_1_0; // @[Top.scala 200:22]
  wire [15:0] n196_O_1_0_1_1; // @[Top.scala 200:22]
  wire [15:0] n196_O_2_0_0_0; // @[Top.scala 200:22]
  wire [15:0] n196_O_2_0_0_1; // @[Top.scala 200:22]
  wire [15:0] n196_O_2_0_1_0; // @[Top.scala 200:22]
  wire [15:0] n196_O_2_0_1_1; // @[Top.scala 200:22]
  wire [15:0] n196_O_3_0_0_0; // @[Top.scala 200:22]
  wire [15:0] n196_O_3_0_0_1; // @[Top.scala 200:22]
  wire [15:0] n196_O_3_0_1_0; // @[Top.scala 200:22]
  wire [15:0] n196_O_3_0_1_1; // @[Top.scala 200:22]
  wire  n203_valid_up; // @[Top.scala 203:22]
  wire  n203_valid_down; // @[Top.scala 203:22]
  wire [15:0] n203_I_0_0_0_0; // @[Top.scala 203:22]
  wire [15:0] n203_I_0_0_0_1; // @[Top.scala 203:22]
  wire [15:0] n203_I_0_0_1_0; // @[Top.scala 203:22]
  wire [15:0] n203_I_0_0_1_1; // @[Top.scala 203:22]
  wire [15:0] n203_I_1_0_0_0; // @[Top.scala 203:22]
  wire [15:0] n203_I_1_0_0_1; // @[Top.scala 203:22]
  wire [15:0] n203_I_1_0_1_0; // @[Top.scala 203:22]
  wire [15:0] n203_I_1_0_1_1; // @[Top.scala 203:22]
  wire [15:0] n203_I_2_0_0_0; // @[Top.scala 203:22]
  wire [15:0] n203_I_2_0_0_1; // @[Top.scala 203:22]
  wire [15:0] n203_I_2_0_1_0; // @[Top.scala 203:22]
  wire [15:0] n203_I_2_0_1_1; // @[Top.scala 203:22]
  wire [15:0] n203_I_3_0_0_0; // @[Top.scala 203:22]
  wire [15:0] n203_I_3_0_0_1; // @[Top.scala 203:22]
  wire [15:0] n203_I_3_0_1_0; // @[Top.scala 203:22]
  wire [15:0] n203_I_3_0_1_1; // @[Top.scala 203:22]
  wire [15:0] n203_O_0_0_0; // @[Top.scala 203:22]
  wire [15:0] n203_O_0_0_1; // @[Top.scala 203:22]
  wire [15:0] n203_O_0_1_0; // @[Top.scala 203:22]
  wire [15:0] n203_O_0_1_1; // @[Top.scala 203:22]
  wire [15:0] n203_O_1_0_0; // @[Top.scala 203:22]
  wire [15:0] n203_O_1_0_1; // @[Top.scala 203:22]
  wire [15:0] n203_O_1_1_0; // @[Top.scala 203:22]
  wire [15:0] n203_O_1_1_1; // @[Top.scala 203:22]
  wire [15:0] n203_O_2_0_0; // @[Top.scala 203:22]
  wire [15:0] n203_O_2_0_1; // @[Top.scala 203:22]
  wire [15:0] n203_O_2_1_0; // @[Top.scala 203:22]
  wire [15:0] n203_O_2_1_1; // @[Top.scala 203:22]
  wire [15:0] n203_O_3_0_0; // @[Top.scala 203:22]
  wire [15:0] n203_O_3_0_1; // @[Top.scala 203:22]
  wire [15:0] n203_O_3_1_0; // @[Top.scala 203:22]
  wire [15:0] n203_O_3_1_1; // @[Top.scala 203:22]
  wire  n245_clock; // @[Top.scala 206:22]
  wire  n245_reset; // @[Top.scala 206:22]
  wire  n245_valid_up; // @[Top.scala 206:22]
  wire  n245_valid_down; // @[Top.scala 206:22]
  wire [15:0] n245_I_0_0_0; // @[Top.scala 206:22]
  wire [15:0] n245_I_0_0_1; // @[Top.scala 206:22]
  wire [15:0] n245_I_0_1_0; // @[Top.scala 206:22]
  wire [15:0] n245_I_0_1_1; // @[Top.scala 206:22]
  wire [15:0] n245_I_1_0_0; // @[Top.scala 206:22]
  wire [15:0] n245_I_1_0_1; // @[Top.scala 206:22]
  wire [15:0] n245_I_1_1_0; // @[Top.scala 206:22]
  wire [15:0] n245_I_1_1_1; // @[Top.scala 206:22]
  wire [15:0] n245_I_2_0_0; // @[Top.scala 206:22]
  wire [15:0] n245_I_2_0_1; // @[Top.scala 206:22]
  wire [15:0] n245_I_2_1_0; // @[Top.scala 206:22]
  wire [15:0] n245_I_2_1_1; // @[Top.scala 206:22]
  wire [15:0] n245_I_3_0_0; // @[Top.scala 206:22]
  wire [15:0] n245_I_3_0_1; // @[Top.scala 206:22]
  wire [15:0] n245_I_3_1_0; // @[Top.scala 206:22]
  wire [15:0] n245_I_3_1_1; // @[Top.scala 206:22]
  wire [15:0] n245_O_0_0_0; // @[Top.scala 206:22]
  wire [15:0] n245_O_1_0_0; // @[Top.scala 206:22]
  wire [15:0] n245_O_2_0_0; // @[Top.scala 206:22]
  wire [15:0] n245_O_3_0_0; // @[Top.scala 206:22]
  wire  n246_valid_up; // @[Top.scala 209:22]
  wire  n246_valid_down; // @[Top.scala 209:22]
  wire [15:0] n246_I_0_0_0; // @[Top.scala 209:22]
  wire [15:0] n246_I_1_0_0; // @[Top.scala 209:22]
  wire [15:0] n246_I_2_0_0; // @[Top.scala 209:22]
  wire [15:0] n246_I_3_0_0; // @[Top.scala 209:22]
  wire [15:0] n246_O_0_0; // @[Top.scala 209:22]
  wire [15:0] n246_O_1_0; // @[Top.scala 209:22]
  wire [15:0] n246_O_2_0; // @[Top.scala 209:22]
  wire [15:0] n246_O_3_0; // @[Top.scala 209:22]
  wire  n247_valid_up; // @[Top.scala 212:22]
  wire  n247_valid_down; // @[Top.scala 212:22]
  wire [15:0] n247_I_0_0; // @[Top.scala 212:22]
  wire [15:0] n247_I_1_0; // @[Top.scala 212:22]
  wire [15:0] n247_I_2_0; // @[Top.scala 212:22]
  wire [15:0] n247_I_3_0; // @[Top.scala 212:22]
  wire [15:0] n247_O_0; // @[Top.scala 212:22]
  wire [15:0] n247_O_1; // @[Top.scala 212:22]
  wire [15:0] n247_O_2; // @[Top.scala 212:22]
  wire [15:0] n247_O_3; // @[Top.scala 212:22]
  wire  n248_clock; // @[Top.scala 215:22]
  wire  n248_reset; // @[Top.scala 215:22]
  wire  n248_valid_up; // @[Top.scala 215:22]
  wire  n248_valid_down; // @[Top.scala 215:22]
  wire [15:0] n248_I_0; // @[Top.scala 215:22]
  wire [15:0] n248_I_1; // @[Top.scala 215:22]
  wire [15:0] n248_I_2; // @[Top.scala 215:22]
  wire [15:0] n248_I_3; // @[Top.scala 215:22]
  wire [15:0] n248_O_0; // @[Top.scala 215:22]
  wire [15:0] n248_O_1; // @[Top.scala 215:22]
  wire [15:0] n248_O_2; // @[Top.scala 215:22]
  wire [15:0] n248_O_3; // @[Top.scala 215:22]
  wire  n249_clock; // @[Top.scala 218:22]
  wire  n249_reset; // @[Top.scala 218:22]
  wire  n249_valid_up; // @[Top.scala 218:22]
  wire  n249_valid_down; // @[Top.scala 218:22]
  wire [15:0] n249_I_0; // @[Top.scala 218:22]
  wire [15:0] n249_I_1; // @[Top.scala 218:22]
  wire [15:0] n249_I_2; // @[Top.scala 218:22]
  wire [15:0] n249_I_3; // @[Top.scala 218:22]
  wire [15:0] n249_O_0; // @[Top.scala 218:22]
  wire [15:0] n249_O_1; // @[Top.scala 218:22]
  wire [15:0] n249_O_2; // @[Top.scala 218:22]
  wire [15:0] n249_O_3; // @[Top.scala 218:22]
  wire  n250_clock; // @[Top.scala 221:22]
  wire  n250_reset; // @[Top.scala 221:22]
  wire  n250_valid_up; // @[Top.scala 221:22]
  wire  n250_valid_down; // @[Top.scala 221:22]
  wire [15:0] n250_I_0; // @[Top.scala 221:22]
  wire [15:0] n250_I_1; // @[Top.scala 221:22]
  wire [15:0] n250_I_2; // @[Top.scala 221:22]
  wire [15:0] n250_I_3; // @[Top.scala 221:22]
  wire [15:0] n250_O_0; // @[Top.scala 221:22]
  wire [15:0] n250_O_1; // @[Top.scala 221:22]
  wire [15:0] n250_O_2; // @[Top.scala 221:22]
  wire [15:0] n250_O_3; // @[Top.scala 221:22]
  FIFO n1 ( // @[Top.scala 75:20]
    .clock(n1_clock),
    .reset(n1_reset),
    .valid_up(n1_valid_up),
    .valid_down(n1_valid_down),
    .I_0(n1_I_0),
    .I_1(n1_I_1),
    .I_2(n1_I_2),
    .I_3(n1_I_3),
    .O_0(n1_O_0),
    .O_1(n1_O_1),
    .O_2(n1_O_2),
    .O_3(n1_O_3)
  );
  ShiftTS n2 ( // @[Top.scala 78:20]
    .clock(n2_clock),
    .reset(n2_reset),
    .valid_up(n2_valid_up),
    .valid_down(n2_valid_down),
    .I_0(n2_I_0),
    .I_1(n2_I_1),
    .I_2(n2_I_2),
    .I_3(n2_I_3),
    .O_0(n2_O_0),
    .O_1(n2_O_1),
    .O_2(n2_O_2),
    .O_3(n2_O_3)
  );
  ShiftTS n3 ( // @[Top.scala 81:20]
    .clock(n3_clock),
    .reset(n3_reset),
    .valid_up(n3_valid_up),
    .valid_down(n3_valid_down),
    .I_0(n3_I_0),
    .I_1(n3_I_1),
    .I_2(n3_I_2),
    .I_3(n3_I_3),
    .O_0(n3_O_0),
    .O_1(n3_O_1),
    .O_2(n3_O_2),
    .O_3(n3_O_3)
  );
  ShiftTS_2 n4 ( // @[Top.scala 84:20]
    .clock(n4_clock),
    .valid_up(n4_valid_up),
    .valid_down(n4_valid_down),
    .I_0(n4_I_0),
    .I_1(n4_I_1),
    .I_2(n4_I_2),
    .I_3(n4_I_3),
    .O_0(n4_O_0),
    .O_1(n4_O_1),
    .O_2(n4_O_2),
    .O_3(n4_O_3)
  );
  ShiftTS_2 n5 ( // @[Top.scala 87:20]
    .clock(n5_clock),
    .valid_up(n5_valid_up),
    .valid_down(n5_valid_down),
    .I_0(n5_I_0),
    .I_1(n5_I_1),
    .I_2(n5_I_2),
    .I_3(n5_I_3),
    .O_0(n5_O_0),
    .O_1(n5_O_1),
    .O_2(n5_O_2),
    .O_3(n5_O_3)
  );
  Map2T n6 ( // @[Top.scala 90:20]
    .valid_up(n6_valid_up),
    .valid_down(n6_valid_down),
    .I0_0(n6_I0_0),
    .I0_1(n6_I0_1),
    .I0_2(n6_I0_2),
    .I0_3(n6_I0_3),
    .I1_0(n6_I1_0),
    .I1_1(n6_I1_1),
    .I1_2(n6_I1_2),
    .I1_3(n6_I1_3),
    .O_0_0(n6_O_0_0),
    .O_0_1(n6_O_0_1),
    .O_1_0(n6_O_1_0),
    .O_1_1(n6_O_1_1),
    .O_2_0(n6_O_2_0),
    .O_2_1(n6_O_2_1),
    .O_3_0(n6_O_3_0),
    .O_3_1(n6_O_3_1)
  );
  Map2T_1 n13 ( // @[Top.scala 94:21]
    .valid_up(n13_valid_up),
    .valid_down(n13_valid_down),
    .I0_0_0(n13_I0_0_0),
    .I0_0_1(n13_I0_0_1),
    .I0_1_0(n13_I0_1_0),
    .I0_1_1(n13_I0_1_1),
    .I0_2_0(n13_I0_2_0),
    .I0_2_1(n13_I0_2_1),
    .I0_3_0(n13_I0_3_0),
    .I0_3_1(n13_I0_3_1),
    .I1_0(n13_I1_0),
    .I1_1(n13_I1_1),
    .I1_2(n13_I1_2),
    .I1_3(n13_I1_3),
    .O_0_0(n13_O_0_0),
    .O_0_1(n13_O_0_1),
    .O_0_2(n13_O_0_2),
    .O_1_0(n13_O_1_0),
    .O_1_1(n13_O_1_1),
    .O_1_2(n13_O_1_2),
    .O_2_0(n13_O_2_0),
    .O_2_1(n13_O_2_1),
    .O_2_2(n13_O_2_2),
    .O_3_0(n13_O_3_0),
    .O_3_1(n13_O_3_1),
    .O_3_2(n13_O_3_2)
  );
  MapT n22 ( // @[Top.scala 98:21]
    .valid_up(n22_valid_up),
    .valid_down(n22_valid_down),
    .I_0_0(n22_I_0_0),
    .I_0_1(n22_I_0_1),
    .I_0_2(n22_I_0_2),
    .I_1_0(n22_I_1_0),
    .I_1_1(n22_I_1_1),
    .I_1_2(n22_I_1_2),
    .I_2_0(n22_I_2_0),
    .I_2_1(n22_I_2_1),
    .I_2_2(n22_I_2_2),
    .I_3_0(n22_I_3_0),
    .I_3_1(n22_I_3_1),
    .I_3_2(n22_I_3_2),
    .O_0_0_0(n22_O_0_0_0),
    .O_0_0_1(n22_O_0_0_1),
    .O_0_0_2(n22_O_0_0_2),
    .O_1_0_0(n22_O_1_0_0),
    .O_1_0_1(n22_O_1_0_1),
    .O_1_0_2(n22_O_1_0_2),
    .O_2_0_0(n22_O_2_0_0),
    .O_2_0_1(n22_O_2_0_1),
    .O_2_0_2(n22_O_2_0_2),
    .O_3_0_0(n22_O_3_0_0),
    .O_3_0_1(n22_O_3_0_1),
    .O_3_0_2(n22_O_3_0_2)
  );
  MapT_1 n29 ( // @[Top.scala 101:21]
    .valid_up(n29_valid_up),
    .valid_down(n29_valid_down),
    .I_0_0_0(n29_I_0_0_0),
    .I_0_0_1(n29_I_0_0_1),
    .I_0_0_2(n29_I_0_0_2),
    .I_1_0_0(n29_I_1_0_0),
    .I_1_0_1(n29_I_1_0_1),
    .I_1_0_2(n29_I_1_0_2),
    .I_2_0_0(n29_I_2_0_0),
    .I_2_0_1(n29_I_2_0_1),
    .I_2_0_2(n29_I_2_0_2),
    .I_3_0_0(n29_I_3_0_0),
    .I_3_0_1(n29_I_3_0_1),
    .I_3_0_2(n29_I_3_0_2),
    .O_0_0(n29_O_0_0),
    .O_0_1(n29_O_0_1),
    .O_0_2(n29_O_0_2),
    .O_1_0(n29_O_1_0),
    .O_1_1(n29_O_1_1),
    .O_1_2(n29_O_1_2),
    .O_2_0(n29_O_2_0),
    .O_2_1(n29_O_2_1),
    .O_2_2(n29_O_2_2),
    .O_3_0(n29_O_3_0),
    .O_3_1(n29_O_3_1),
    .O_3_2(n29_O_3_2)
  );
  ShiftTS_2 n30 ( // @[Top.scala 104:21]
    .clock(n30_clock),
    .valid_up(n30_valid_up),
    .valid_down(n30_valid_down),
    .I_0(n30_I_0),
    .I_1(n30_I_1),
    .I_2(n30_I_2),
    .I_3(n30_I_3),
    .O_0(n30_O_0),
    .O_1(n30_O_1),
    .O_2(n30_O_2),
    .O_3(n30_O_3)
  );
  ShiftTS_2 n31 ( // @[Top.scala 107:21]
    .clock(n31_clock),
    .valid_up(n31_valid_up),
    .valid_down(n31_valid_down),
    .I_0(n31_I_0),
    .I_1(n31_I_1),
    .I_2(n31_I_2),
    .I_3(n31_I_3),
    .O_0(n31_O_0),
    .O_1(n31_O_1),
    .O_2(n31_O_2),
    .O_3(n31_O_3)
  );
  Map2T n32 ( // @[Top.scala 110:21]
    .valid_up(n32_valid_up),
    .valid_down(n32_valid_down),
    .I0_0(n32_I0_0),
    .I0_1(n32_I0_1),
    .I0_2(n32_I0_2),
    .I0_3(n32_I0_3),
    .I1_0(n32_I1_0),
    .I1_1(n32_I1_1),
    .I1_2(n32_I1_2),
    .I1_3(n32_I1_3),
    .O_0_0(n32_O_0_0),
    .O_0_1(n32_O_0_1),
    .O_1_0(n32_O_1_0),
    .O_1_1(n32_O_1_1),
    .O_2_0(n32_O_2_0),
    .O_2_1(n32_O_2_1),
    .O_3_0(n32_O_3_0),
    .O_3_1(n32_O_3_1)
  );
  Map2T_1 n39 ( // @[Top.scala 114:21]
    .valid_up(n39_valid_up),
    .valid_down(n39_valid_down),
    .I0_0_0(n39_I0_0_0),
    .I0_0_1(n39_I0_0_1),
    .I0_1_0(n39_I0_1_0),
    .I0_1_1(n39_I0_1_1),
    .I0_2_0(n39_I0_2_0),
    .I0_2_1(n39_I0_2_1),
    .I0_3_0(n39_I0_3_0),
    .I0_3_1(n39_I0_3_1),
    .I1_0(n39_I1_0),
    .I1_1(n39_I1_1),
    .I1_2(n39_I1_2),
    .I1_3(n39_I1_3),
    .O_0_0(n39_O_0_0),
    .O_0_1(n39_O_0_1),
    .O_0_2(n39_O_0_2),
    .O_1_0(n39_O_1_0),
    .O_1_1(n39_O_1_1),
    .O_1_2(n39_O_1_2),
    .O_2_0(n39_O_2_0),
    .O_2_1(n39_O_2_1),
    .O_2_2(n39_O_2_2),
    .O_3_0(n39_O_3_0),
    .O_3_1(n39_O_3_1),
    .O_3_2(n39_O_3_2)
  );
  MapT n48 ( // @[Top.scala 118:21]
    .valid_up(n48_valid_up),
    .valid_down(n48_valid_down),
    .I_0_0(n48_I_0_0),
    .I_0_1(n48_I_0_1),
    .I_0_2(n48_I_0_2),
    .I_1_0(n48_I_1_0),
    .I_1_1(n48_I_1_1),
    .I_1_2(n48_I_1_2),
    .I_2_0(n48_I_2_0),
    .I_2_1(n48_I_2_1),
    .I_2_2(n48_I_2_2),
    .I_3_0(n48_I_3_0),
    .I_3_1(n48_I_3_1),
    .I_3_2(n48_I_3_2),
    .O_0_0_0(n48_O_0_0_0),
    .O_0_0_1(n48_O_0_0_1),
    .O_0_0_2(n48_O_0_0_2),
    .O_1_0_0(n48_O_1_0_0),
    .O_1_0_1(n48_O_1_0_1),
    .O_1_0_2(n48_O_1_0_2),
    .O_2_0_0(n48_O_2_0_0),
    .O_2_0_1(n48_O_2_0_1),
    .O_2_0_2(n48_O_2_0_2),
    .O_3_0_0(n48_O_3_0_0),
    .O_3_0_1(n48_O_3_0_1),
    .O_3_0_2(n48_O_3_0_2)
  );
  MapT_1 n55 ( // @[Top.scala 121:21]
    .valid_up(n55_valid_up),
    .valid_down(n55_valid_down),
    .I_0_0_0(n55_I_0_0_0),
    .I_0_0_1(n55_I_0_0_1),
    .I_0_0_2(n55_I_0_0_2),
    .I_1_0_0(n55_I_1_0_0),
    .I_1_0_1(n55_I_1_0_1),
    .I_1_0_2(n55_I_1_0_2),
    .I_2_0_0(n55_I_2_0_0),
    .I_2_0_1(n55_I_2_0_1),
    .I_2_0_2(n55_I_2_0_2),
    .I_3_0_0(n55_I_3_0_0),
    .I_3_0_1(n55_I_3_0_1),
    .I_3_0_2(n55_I_3_0_2),
    .O_0_0(n55_O_0_0),
    .O_0_1(n55_O_0_1),
    .O_0_2(n55_O_0_2),
    .O_1_0(n55_O_1_0),
    .O_1_1(n55_O_1_1),
    .O_1_2(n55_O_1_2),
    .O_2_0(n55_O_2_0),
    .O_2_1(n55_O_2_1),
    .O_2_2(n55_O_2_2),
    .O_3_0(n55_O_3_0),
    .O_3_1(n55_O_3_1),
    .O_3_2(n55_O_3_2)
  );
  Map2T_4 n56 ( // @[Top.scala 124:21]
    .valid_up(n56_valid_up),
    .valid_down(n56_valid_down),
    .I0_0_0(n56_I0_0_0),
    .I0_0_1(n56_I0_0_1),
    .I0_0_2(n56_I0_0_2),
    .I0_1_0(n56_I0_1_0),
    .I0_1_1(n56_I0_1_1),
    .I0_1_2(n56_I0_1_2),
    .I0_2_0(n56_I0_2_0),
    .I0_2_1(n56_I0_2_1),
    .I0_2_2(n56_I0_2_2),
    .I0_3_0(n56_I0_3_0),
    .I0_3_1(n56_I0_3_1),
    .I0_3_2(n56_I0_3_2),
    .I1_0_0(n56_I1_0_0),
    .I1_0_1(n56_I1_0_1),
    .I1_0_2(n56_I1_0_2),
    .I1_1_0(n56_I1_1_0),
    .I1_1_1(n56_I1_1_1),
    .I1_1_2(n56_I1_1_2),
    .I1_2_0(n56_I1_2_0),
    .I1_2_1(n56_I1_2_1),
    .I1_2_2(n56_I1_2_2),
    .I1_3_0(n56_I1_3_0),
    .I1_3_1(n56_I1_3_1),
    .I1_3_2(n56_I1_3_2),
    .O_0_0_0(n56_O_0_0_0),
    .O_0_0_1(n56_O_0_0_1),
    .O_0_0_2(n56_O_0_0_2),
    .O_0_1_0(n56_O_0_1_0),
    .O_0_1_1(n56_O_0_1_1),
    .O_0_1_2(n56_O_0_1_2),
    .O_1_0_0(n56_O_1_0_0),
    .O_1_0_1(n56_O_1_0_1),
    .O_1_0_2(n56_O_1_0_2),
    .O_1_1_0(n56_O_1_1_0),
    .O_1_1_1(n56_O_1_1_1),
    .O_1_1_2(n56_O_1_1_2),
    .O_2_0_0(n56_O_2_0_0),
    .O_2_0_1(n56_O_2_0_1),
    .O_2_0_2(n56_O_2_0_2),
    .O_2_1_0(n56_O_2_1_0),
    .O_2_1_1(n56_O_2_1_1),
    .O_2_1_2(n56_O_2_1_2),
    .O_3_0_0(n56_O_3_0_0),
    .O_3_0_1(n56_O_3_0_1),
    .O_3_0_2(n56_O_3_0_2),
    .O_3_1_0(n56_O_3_1_0),
    .O_3_1_1(n56_O_3_1_1),
    .O_3_1_2(n56_O_3_1_2)
  );
  ShiftTS_2 n63 ( // @[Top.scala 128:21]
    .clock(n63_clock),
    .valid_up(n63_valid_up),
    .valid_down(n63_valid_down),
    .I_0(n63_I_0),
    .I_1(n63_I_1),
    .I_2(n63_I_2),
    .I_3(n63_I_3),
    .O_0(n63_O_0),
    .O_1(n63_O_1),
    .O_2(n63_O_2),
    .O_3(n63_O_3)
  );
  ShiftTS_2 n64 ( // @[Top.scala 131:21]
    .clock(n64_clock),
    .valid_up(n64_valid_up),
    .valid_down(n64_valid_down),
    .I_0(n64_I_0),
    .I_1(n64_I_1),
    .I_2(n64_I_2),
    .I_3(n64_I_3),
    .O_0(n64_O_0),
    .O_1(n64_O_1),
    .O_2(n64_O_2),
    .O_3(n64_O_3)
  );
  Map2T n65 ( // @[Top.scala 134:21]
    .valid_up(n65_valid_up),
    .valid_down(n65_valid_down),
    .I0_0(n65_I0_0),
    .I0_1(n65_I0_1),
    .I0_2(n65_I0_2),
    .I0_3(n65_I0_3),
    .I1_0(n65_I1_0),
    .I1_1(n65_I1_1),
    .I1_2(n65_I1_2),
    .I1_3(n65_I1_3),
    .O_0_0(n65_O_0_0),
    .O_0_1(n65_O_0_1),
    .O_1_0(n65_O_1_0),
    .O_1_1(n65_O_1_1),
    .O_2_0(n65_O_2_0),
    .O_2_1(n65_O_2_1),
    .O_3_0(n65_O_3_0),
    .O_3_1(n65_O_3_1)
  );
  Map2T_1 n72 ( // @[Top.scala 138:21]
    .valid_up(n72_valid_up),
    .valid_down(n72_valid_down),
    .I0_0_0(n72_I0_0_0),
    .I0_0_1(n72_I0_0_1),
    .I0_1_0(n72_I0_1_0),
    .I0_1_1(n72_I0_1_1),
    .I0_2_0(n72_I0_2_0),
    .I0_2_1(n72_I0_2_1),
    .I0_3_0(n72_I0_3_0),
    .I0_3_1(n72_I0_3_1),
    .I1_0(n72_I1_0),
    .I1_1(n72_I1_1),
    .I1_2(n72_I1_2),
    .I1_3(n72_I1_3),
    .O_0_0(n72_O_0_0),
    .O_0_1(n72_O_0_1),
    .O_0_2(n72_O_0_2),
    .O_1_0(n72_O_1_0),
    .O_1_1(n72_O_1_1),
    .O_1_2(n72_O_1_2),
    .O_2_0(n72_O_2_0),
    .O_2_1(n72_O_2_1),
    .O_2_2(n72_O_2_2),
    .O_3_0(n72_O_3_0),
    .O_3_1(n72_O_3_1),
    .O_3_2(n72_O_3_2)
  );
  MapT n81 ( // @[Top.scala 142:21]
    .valid_up(n81_valid_up),
    .valid_down(n81_valid_down),
    .I_0_0(n81_I_0_0),
    .I_0_1(n81_I_0_1),
    .I_0_2(n81_I_0_2),
    .I_1_0(n81_I_1_0),
    .I_1_1(n81_I_1_1),
    .I_1_2(n81_I_1_2),
    .I_2_0(n81_I_2_0),
    .I_2_1(n81_I_2_1),
    .I_2_2(n81_I_2_2),
    .I_3_0(n81_I_3_0),
    .I_3_1(n81_I_3_1),
    .I_3_2(n81_I_3_2),
    .O_0_0_0(n81_O_0_0_0),
    .O_0_0_1(n81_O_0_0_1),
    .O_0_0_2(n81_O_0_0_2),
    .O_1_0_0(n81_O_1_0_0),
    .O_1_0_1(n81_O_1_0_1),
    .O_1_0_2(n81_O_1_0_2),
    .O_2_0_0(n81_O_2_0_0),
    .O_2_0_1(n81_O_2_0_1),
    .O_2_0_2(n81_O_2_0_2),
    .O_3_0_0(n81_O_3_0_0),
    .O_3_0_1(n81_O_3_0_1),
    .O_3_0_2(n81_O_3_0_2)
  );
  MapT_1 n88 ( // @[Top.scala 145:21]
    .valid_up(n88_valid_up),
    .valid_down(n88_valid_down),
    .I_0_0_0(n88_I_0_0_0),
    .I_0_0_1(n88_I_0_0_1),
    .I_0_0_2(n88_I_0_0_2),
    .I_1_0_0(n88_I_1_0_0),
    .I_1_0_1(n88_I_1_0_1),
    .I_1_0_2(n88_I_1_0_2),
    .I_2_0_0(n88_I_2_0_0),
    .I_2_0_1(n88_I_2_0_1),
    .I_2_0_2(n88_I_2_0_2),
    .I_3_0_0(n88_I_3_0_0),
    .I_3_0_1(n88_I_3_0_1),
    .I_3_0_2(n88_I_3_0_2),
    .O_0_0(n88_O_0_0),
    .O_0_1(n88_O_0_1),
    .O_0_2(n88_O_0_2),
    .O_1_0(n88_O_1_0),
    .O_1_1(n88_O_1_1),
    .O_1_2(n88_O_1_2),
    .O_2_0(n88_O_2_0),
    .O_2_1(n88_O_2_1),
    .O_2_2(n88_O_2_2),
    .O_3_0(n88_O_3_0),
    .O_3_1(n88_O_3_1),
    .O_3_2(n88_O_3_2)
  );
  Map2T_7 n89 ( // @[Top.scala 148:21]
    .valid_up(n89_valid_up),
    .valid_down(n89_valid_down),
    .I0_0_0_0(n89_I0_0_0_0),
    .I0_0_0_1(n89_I0_0_0_1),
    .I0_0_0_2(n89_I0_0_0_2),
    .I0_0_1_0(n89_I0_0_1_0),
    .I0_0_1_1(n89_I0_0_1_1),
    .I0_0_1_2(n89_I0_0_1_2),
    .I0_1_0_0(n89_I0_1_0_0),
    .I0_1_0_1(n89_I0_1_0_1),
    .I0_1_0_2(n89_I0_1_0_2),
    .I0_1_1_0(n89_I0_1_1_0),
    .I0_1_1_1(n89_I0_1_1_1),
    .I0_1_1_2(n89_I0_1_1_2),
    .I0_2_0_0(n89_I0_2_0_0),
    .I0_2_0_1(n89_I0_2_0_1),
    .I0_2_0_2(n89_I0_2_0_2),
    .I0_2_1_0(n89_I0_2_1_0),
    .I0_2_1_1(n89_I0_2_1_1),
    .I0_2_1_2(n89_I0_2_1_2),
    .I0_3_0_0(n89_I0_3_0_0),
    .I0_3_0_1(n89_I0_3_0_1),
    .I0_3_0_2(n89_I0_3_0_2),
    .I0_3_1_0(n89_I0_3_1_0),
    .I0_3_1_1(n89_I0_3_1_1),
    .I0_3_1_2(n89_I0_3_1_2),
    .I1_0_0(n89_I1_0_0),
    .I1_0_1(n89_I1_0_1),
    .I1_0_2(n89_I1_0_2),
    .I1_1_0(n89_I1_1_0),
    .I1_1_1(n89_I1_1_1),
    .I1_1_2(n89_I1_1_2),
    .I1_2_0(n89_I1_2_0),
    .I1_2_1(n89_I1_2_1),
    .I1_2_2(n89_I1_2_2),
    .I1_3_0(n89_I1_3_0),
    .I1_3_1(n89_I1_3_1),
    .I1_3_2(n89_I1_3_2),
    .O_0_0_0(n89_O_0_0_0),
    .O_0_0_1(n89_O_0_0_1),
    .O_0_0_2(n89_O_0_0_2),
    .O_0_1_0(n89_O_0_1_0),
    .O_0_1_1(n89_O_0_1_1),
    .O_0_1_2(n89_O_0_1_2),
    .O_0_2_0(n89_O_0_2_0),
    .O_0_2_1(n89_O_0_2_1),
    .O_0_2_2(n89_O_0_2_2),
    .O_1_0_0(n89_O_1_0_0),
    .O_1_0_1(n89_O_1_0_1),
    .O_1_0_2(n89_O_1_0_2),
    .O_1_1_0(n89_O_1_1_0),
    .O_1_1_1(n89_O_1_1_1),
    .O_1_1_2(n89_O_1_1_2),
    .O_1_2_0(n89_O_1_2_0),
    .O_1_2_1(n89_O_1_2_1),
    .O_1_2_2(n89_O_1_2_2),
    .O_2_0_0(n89_O_2_0_0),
    .O_2_0_1(n89_O_2_0_1),
    .O_2_0_2(n89_O_2_0_2),
    .O_2_1_0(n89_O_2_1_0),
    .O_2_1_1(n89_O_2_1_1),
    .O_2_1_2(n89_O_2_1_2),
    .O_2_2_0(n89_O_2_2_0),
    .O_2_2_1(n89_O_2_2_1),
    .O_2_2_2(n89_O_2_2_2),
    .O_3_0_0(n89_O_3_0_0),
    .O_3_0_1(n89_O_3_0_1),
    .O_3_0_2(n89_O_3_0_2),
    .O_3_1_0(n89_O_3_1_0),
    .O_3_1_1(n89_O_3_1_1),
    .O_3_1_2(n89_O_3_1_2),
    .O_3_2_0(n89_O_3_2_0),
    .O_3_2_1(n89_O_3_2_1),
    .O_3_2_2(n89_O_3_2_2)
  );
  MapT_6 n98 ( // @[Top.scala 152:21]
    .valid_up(n98_valid_up),
    .valid_down(n98_valid_down),
    .I_0_0_0(n98_I_0_0_0),
    .I_0_0_1(n98_I_0_0_1),
    .I_0_0_2(n98_I_0_0_2),
    .I_0_1_0(n98_I_0_1_0),
    .I_0_1_1(n98_I_0_1_1),
    .I_0_1_2(n98_I_0_1_2),
    .I_0_2_0(n98_I_0_2_0),
    .I_0_2_1(n98_I_0_2_1),
    .I_0_2_2(n98_I_0_2_2),
    .I_1_0_0(n98_I_1_0_0),
    .I_1_0_1(n98_I_1_0_1),
    .I_1_0_2(n98_I_1_0_2),
    .I_1_1_0(n98_I_1_1_0),
    .I_1_1_1(n98_I_1_1_1),
    .I_1_1_2(n98_I_1_1_2),
    .I_1_2_0(n98_I_1_2_0),
    .I_1_2_1(n98_I_1_2_1),
    .I_1_2_2(n98_I_1_2_2),
    .I_2_0_0(n98_I_2_0_0),
    .I_2_0_1(n98_I_2_0_1),
    .I_2_0_2(n98_I_2_0_2),
    .I_2_1_0(n98_I_2_1_0),
    .I_2_1_1(n98_I_2_1_1),
    .I_2_1_2(n98_I_2_1_2),
    .I_2_2_0(n98_I_2_2_0),
    .I_2_2_1(n98_I_2_2_1),
    .I_2_2_2(n98_I_2_2_2),
    .I_3_0_0(n98_I_3_0_0),
    .I_3_0_1(n98_I_3_0_1),
    .I_3_0_2(n98_I_3_0_2),
    .I_3_1_0(n98_I_3_1_0),
    .I_3_1_1(n98_I_3_1_1),
    .I_3_1_2(n98_I_3_1_2),
    .I_3_2_0(n98_I_3_2_0),
    .I_3_2_1(n98_I_3_2_1),
    .I_3_2_2(n98_I_3_2_2),
    .O_0_0_0_0(n98_O_0_0_0_0),
    .O_0_0_0_1(n98_O_0_0_0_1),
    .O_0_0_0_2(n98_O_0_0_0_2),
    .O_0_0_1_0(n98_O_0_0_1_0),
    .O_0_0_1_1(n98_O_0_0_1_1),
    .O_0_0_1_2(n98_O_0_0_1_2),
    .O_0_0_2_0(n98_O_0_0_2_0),
    .O_0_0_2_1(n98_O_0_0_2_1),
    .O_0_0_2_2(n98_O_0_0_2_2),
    .O_1_0_0_0(n98_O_1_0_0_0),
    .O_1_0_0_1(n98_O_1_0_0_1),
    .O_1_0_0_2(n98_O_1_0_0_2),
    .O_1_0_1_0(n98_O_1_0_1_0),
    .O_1_0_1_1(n98_O_1_0_1_1),
    .O_1_0_1_2(n98_O_1_0_1_2),
    .O_1_0_2_0(n98_O_1_0_2_0),
    .O_1_0_2_1(n98_O_1_0_2_1),
    .O_1_0_2_2(n98_O_1_0_2_2),
    .O_2_0_0_0(n98_O_2_0_0_0),
    .O_2_0_0_1(n98_O_2_0_0_1),
    .O_2_0_0_2(n98_O_2_0_0_2),
    .O_2_0_1_0(n98_O_2_0_1_0),
    .O_2_0_1_1(n98_O_2_0_1_1),
    .O_2_0_1_2(n98_O_2_0_1_2),
    .O_2_0_2_0(n98_O_2_0_2_0),
    .O_2_0_2_1(n98_O_2_0_2_1),
    .O_2_0_2_2(n98_O_2_0_2_2),
    .O_3_0_0_0(n98_O_3_0_0_0),
    .O_3_0_0_1(n98_O_3_0_0_1),
    .O_3_0_0_2(n98_O_3_0_0_2),
    .O_3_0_1_0(n98_O_3_0_1_0),
    .O_3_0_1_1(n98_O_3_0_1_1),
    .O_3_0_1_2(n98_O_3_0_1_2),
    .O_3_0_2_0(n98_O_3_0_2_0),
    .O_3_0_2_1(n98_O_3_0_2_1),
    .O_3_0_2_2(n98_O_3_0_2_2)
  );
  MapT_7 n105 ( // @[Top.scala 155:22]
    .valid_up(n105_valid_up),
    .valid_down(n105_valid_down),
    .I_0_0_0_0(n105_I_0_0_0_0),
    .I_0_0_0_1(n105_I_0_0_0_1),
    .I_0_0_0_2(n105_I_0_0_0_2),
    .I_0_0_1_0(n105_I_0_0_1_0),
    .I_0_0_1_1(n105_I_0_0_1_1),
    .I_0_0_1_2(n105_I_0_0_1_2),
    .I_0_0_2_0(n105_I_0_0_2_0),
    .I_0_0_2_1(n105_I_0_0_2_1),
    .I_0_0_2_2(n105_I_0_0_2_2),
    .I_1_0_0_0(n105_I_1_0_0_0),
    .I_1_0_0_1(n105_I_1_0_0_1),
    .I_1_0_0_2(n105_I_1_0_0_2),
    .I_1_0_1_0(n105_I_1_0_1_0),
    .I_1_0_1_1(n105_I_1_0_1_1),
    .I_1_0_1_2(n105_I_1_0_1_2),
    .I_1_0_2_0(n105_I_1_0_2_0),
    .I_1_0_2_1(n105_I_1_0_2_1),
    .I_1_0_2_2(n105_I_1_0_2_2),
    .I_2_0_0_0(n105_I_2_0_0_0),
    .I_2_0_0_1(n105_I_2_0_0_1),
    .I_2_0_0_2(n105_I_2_0_0_2),
    .I_2_0_1_0(n105_I_2_0_1_0),
    .I_2_0_1_1(n105_I_2_0_1_1),
    .I_2_0_1_2(n105_I_2_0_1_2),
    .I_2_0_2_0(n105_I_2_0_2_0),
    .I_2_0_2_1(n105_I_2_0_2_1),
    .I_2_0_2_2(n105_I_2_0_2_2),
    .I_3_0_0_0(n105_I_3_0_0_0),
    .I_3_0_0_1(n105_I_3_0_0_1),
    .I_3_0_0_2(n105_I_3_0_0_2),
    .I_3_0_1_0(n105_I_3_0_1_0),
    .I_3_0_1_1(n105_I_3_0_1_1),
    .I_3_0_1_2(n105_I_3_0_1_2),
    .I_3_0_2_0(n105_I_3_0_2_0),
    .I_3_0_2_1(n105_I_3_0_2_1),
    .I_3_0_2_2(n105_I_3_0_2_2),
    .O_0_0_0(n105_O_0_0_0),
    .O_0_0_1(n105_O_0_0_1),
    .O_0_0_2(n105_O_0_0_2),
    .O_0_1_0(n105_O_0_1_0),
    .O_0_1_1(n105_O_0_1_1),
    .O_0_1_2(n105_O_0_1_2),
    .O_0_2_0(n105_O_0_2_0),
    .O_0_2_1(n105_O_0_2_1),
    .O_0_2_2(n105_O_0_2_2),
    .O_1_0_0(n105_O_1_0_0),
    .O_1_0_1(n105_O_1_0_1),
    .O_1_0_2(n105_O_1_0_2),
    .O_1_1_0(n105_O_1_1_0),
    .O_1_1_1(n105_O_1_1_1),
    .O_1_1_2(n105_O_1_1_2),
    .O_1_2_0(n105_O_1_2_0),
    .O_1_2_1(n105_O_1_2_1),
    .O_1_2_2(n105_O_1_2_2),
    .O_2_0_0(n105_O_2_0_0),
    .O_2_0_1(n105_O_2_0_1),
    .O_2_0_2(n105_O_2_0_2),
    .O_2_1_0(n105_O_2_1_0),
    .O_2_1_1(n105_O_2_1_1),
    .O_2_1_2(n105_O_2_1_2),
    .O_2_2_0(n105_O_2_2_0),
    .O_2_2_1(n105_O_2_2_1),
    .O_2_2_2(n105_O_2_2_2),
    .O_3_0_0(n105_O_3_0_0),
    .O_3_0_1(n105_O_3_0_1),
    .O_3_0_2(n105_O_3_0_2),
    .O_3_1_0(n105_O_3_1_0),
    .O_3_1_1(n105_O_3_1_1),
    .O_3_1_2(n105_O_3_1_2),
    .O_3_2_0(n105_O_3_2_0),
    .O_3_2_1(n105_O_3_2_1),
    .O_3_2_2(n105_O_3_2_2)
  );
  MapT_8 n147 ( // @[Top.scala 158:22]
    .clock(n147_clock),
    .reset(n147_reset),
    .valid_up(n147_valid_up),
    .valid_down(n147_valid_down),
    .I_0_0_0(n147_I_0_0_0),
    .I_0_0_1(n147_I_0_0_1),
    .I_0_0_2(n147_I_0_0_2),
    .I_0_1_0(n147_I_0_1_0),
    .I_0_1_1(n147_I_0_1_1),
    .I_0_1_2(n147_I_0_1_2),
    .I_0_2_0(n147_I_0_2_0),
    .I_0_2_1(n147_I_0_2_1),
    .I_0_2_2(n147_I_0_2_2),
    .I_1_0_0(n147_I_1_0_0),
    .I_1_0_1(n147_I_1_0_1),
    .I_1_0_2(n147_I_1_0_2),
    .I_1_1_0(n147_I_1_1_0),
    .I_1_1_1(n147_I_1_1_1),
    .I_1_1_2(n147_I_1_1_2),
    .I_1_2_0(n147_I_1_2_0),
    .I_1_2_1(n147_I_1_2_1),
    .I_1_2_2(n147_I_1_2_2),
    .I_2_0_0(n147_I_2_0_0),
    .I_2_0_1(n147_I_2_0_1),
    .I_2_0_2(n147_I_2_0_2),
    .I_2_1_0(n147_I_2_1_0),
    .I_2_1_1(n147_I_2_1_1),
    .I_2_1_2(n147_I_2_1_2),
    .I_2_2_0(n147_I_2_2_0),
    .I_2_2_1(n147_I_2_2_1),
    .I_2_2_2(n147_I_2_2_2),
    .I_3_0_0(n147_I_3_0_0),
    .I_3_0_1(n147_I_3_0_1),
    .I_3_0_2(n147_I_3_0_2),
    .I_3_1_0(n147_I_3_1_0),
    .I_3_1_1(n147_I_3_1_1),
    .I_3_1_2(n147_I_3_1_2),
    .I_3_2_0(n147_I_3_2_0),
    .I_3_2_1(n147_I_3_2_1),
    .I_3_2_2(n147_I_3_2_2),
    .O_0_0_0(n147_O_0_0_0),
    .O_1_0_0(n147_O_1_0_0),
    .O_2_0_0(n147_O_2_0_0),
    .O_3_0_0(n147_O_3_0_0)
  );
  Passthrough n148 ( // @[Top.scala 161:22]
    .valid_up(n148_valid_up),
    .valid_down(n148_valid_down),
    .I_0_0_0(n148_I_0_0_0),
    .I_1_0_0(n148_I_1_0_0),
    .I_2_0_0(n148_I_2_0_0),
    .I_3_0_0(n148_I_3_0_0),
    .O_0_0(n148_O_0_0),
    .O_1_0(n148_O_1_0),
    .O_2_0(n148_O_2_0),
    .O_3_0(n148_O_3_0)
  );
  Passthrough_1 n149 ( // @[Top.scala 164:22]
    .valid_up(n149_valid_up),
    .valid_down(n149_valid_down),
    .I_0_0(n149_I_0_0),
    .I_1_0(n149_I_1_0),
    .I_2_0(n149_I_2_0),
    .I_3_0(n149_I_3_0),
    .O_0(n149_O_0),
    .O_1(n149_O_1),
    .O_2(n149_O_2),
    .O_3(n149_O_3)
  );
  ShiftTS n150 ( // @[Top.scala 167:22]
    .clock(n150_clock),
    .reset(n150_reset),
    .valid_up(n150_valid_up),
    .valid_down(n150_valid_down),
    .I_0(n150_I_0),
    .I_1(n150_I_1),
    .I_2(n150_I_2),
    .I_3(n150_I_3),
    .O_0(n150_O_0),
    .O_1(n150_O_1),
    .O_2(n150_O_2),
    .O_3(n150_O_3)
  );
  ShiftTS_2 n151 ( // @[Top.scala 170:22]
    .clock(n151_clock),
    .valid_up(n151_valid_up),
    .valid_down(n151_valid_down),
    .I_0(n151_I_0),
    .I_1(n151_I_1),
    .I_2(n151_I_2),
    .I_3(n151_I_3),
    .O_0(n151_O_0),
    .O_1(n151_O_1),
    .O_2(n151_O_2),
    .O_3(n151_O_3)
  );
  Map2T n152 ( // @[Top.scala 173:22]
    .valid_up(n152_valid_up),
    .valid_down(n152_valid_down),
    .I0_0(n152_I0_0),
    .I0_1(n152_I0_1),
    .I0_2(n152_I0_2),
    .I0_3(n152_I0_3),
    .I1_0(n152_I1_0),
    .I1_1(n152_I1_1),
    .I1_2(n152_I1_2),
    .I1_3(n152_I1_3),
    .O_0_0(n152_O_0_0),
    .O_0_1(n152_O_0_1),
    .O_1_0(n152_O_1_0),
    .O_1_1(n152_O_1_1),
    .O_2_0(n152_O_2_0),
    .O_2_1(n152_O_2_1),
    .O_3_0(n152_O_3_0),
    .O_3_1(n152_O_3_1)
  );
  MapT_9 n161 ( // @[Top.scala 177:22]
    .valid_up(n161_valid_up),
    .valid_down(n161_valid_down),
    .I_0_0(n161_I_0_0),
    .I_0_1(n161_I_0_1),
    .I_1_0(n161_I_1_0),
    .I_1_1(n161_I_1_1),
    .I_2_0(n161_I_2_0),
    .I_2_1(n161_I_2_1),
    .I_3_0(n161_I_3_0),
    .I_3_1(n161_I_3_1),
    .O_0_0_0(n161_O_0_0_0),
    .O_0_0_1(n161_O_0_0_1),
    .O_1_0_0(n161_O_1_0_0),
    .O_1_0_1(n161_O_1_0_1),
    .O_2_0_0(n161_O_2_0_0),
    .O_2_0_1(n161_O_2_0_1),
    .O_3_0_0(n161_O_3_0_0),
    .O_3_0_1(n161_O_3_0_1)
  );
  MapT_10 n168 ( // @[Top.scala 180:22]
    .valid_up(n168_valid_up),
    .valid_down(n168_valid_down),
    .I_0_0_0(n168_I_0_0_0),
    .I_0_0_1(n168_I_0_0_1),
    .I_1_0_0(n168_I_1_0_0),
    .I_1_0_1(n168_I_1_0_1),
    .I_2_0_0(n168_I_2_0_0),
    .I_2_0_1(n168_I_2_0_1),
    .I_3_0_0(n168_I_3_0_0),
    .I_3_0_1(n168_I_3_0_1),
    .O_0_0(n168_O_0_0),
    .O_0_1(n168_O_0_1),
    .O_1_0(n168_O_1_0),
    .O_1_1(n168_O_1_1),
    .O_2_0(n168_O_2_0),
    .O_2_1(n168_O_2_1),
    .O_3_0(n168_O_3_0),
    .O_3_1(n168_O_3_1)
  );
  ShiftTS_2 n169 ( // @[Top.scala 183:22]
    .clock(n169_clock),
    .valid_up(n169_valid_up),
    .valid_down(n169_valid_down),
    .I_0(n169_I_0),
    .I_1(n169_I_1),
    .I_2(n169_I_2),
    .I_3(n169_I_3),
    .O_0(n169_O_0),
    .O_1(n169_O_1),
    .O_2(n169_O_2),
    .O_3(n169_O_3)
  );
  Map2T n170 ( // @[Top.scala 186:22]
    .valid_up(n170_valid_up),
    .valid_down(n170_valid_down),
    .I0_0(n170_I0_0),
    .I0_1(n170_I0_1),
    .I0_2(n170_I0_2),
    .I0_3(n170_I0_3),
    .I1_0(n170_I1_0),
    .I1_1(n170_I1_1),
    .I1_2(n170_I1_2),
    .I1_3(n170_I1_3),
    .O_0_0(n170_O_0_0),
    .O_0_1(n170_O_0_1),
    .O_1_0(n170_O_1_0),
    .O_1_1(n170_O_1_1),
    .O_2_0(n170_O_2_0),
    .O_2_1(n170_O_2_1),
    .O_3_0(n170_O_3_0),
    .O_3_1(n170_O_3_1)
  );
  MapT_9 n179 ( // @[Top.scala 190:22]
    .valid_up(n179_valid_up),
    .valid_down(n179_valid_down),
    .I_0_0(n179_I_0_0),
    .I_0_1(n179_I_0_1),
    .I_1_0(n179_I_1_0),
    .I_1_1(n179_I_1_1),
    .I_2_0(n179_I_2_0),
    .I_2_1(n179_I_2_1),
    .I_3_0(n179_I_3_0),
    .I_3_1(n179_I_3_1),
    .O_0_0_0(n179_O_0_0_0),
    .O_0_0_1(n179_O_0_0_1),
    .O_1_0_0(n179_O_1_0_0),
    .O_1_0_1(n179_O_1_0_1),
    .O_2_0_0(n179_O_2_0_0),
    .O_2_0_1(n179_O_2_0_1),
    .O_3_0_0(n179_O_3_0_0),
    .O_3_0_1(n179_O_3_0_1)
  );
  MapT_10 n186 ( // @[Top.scala 193:22]
    .valid_up(n186_valid_up),
    .valid_down(n186_valid_down),
    .I_0_0_0(n186_I_0_0_0),
    .I_0_0_1(n186_I_0_0_1),
    .I_1_0_0(n186_I_1_0_0),
    .I_1_0_1(n186_I_1_0_1),
    .I_2_0_0(n186_I_2_0_0),
    .I_2_0_1(n186_I_2_0_1),
    .I_3_0_0(n186_I_3_0_0),
    .I_3_0_1(n186_I_3_0_1),
    .O_0_0(n186_O_0_0),
    .O_0_1(n186_O_0_1),
    .O_1_0(n186_O_1_0),
    .O_1_1(n186_O_1_1),
    .O_2_0(n186_O_2_0),
    .O_2_1(n186_O_2_1),
    .O_3_0(n186_O_3_0),
    .O_3_1(n186_O_3_1)
  );
  Map2T_10 n187 ( // @[Top.scala 196:22]
    .valid_up(n187_valid_up),
    .valid_down(n187_valid_down),
    .I0_0_0(n187_I0_0_0),
    .I0_0_1(n187_I0_0_1),
    .I0_1_0(n187_I0_1_0),
    .I0_1_1(n187_I0_1_1),
    .I0_2_0(n187_I0_2_0),
    .I0_2_1(n187_I0_2_1),
    .I0_3_0(n187_I0_3_0),
    .I0_3_1(n187_I0_3_1),
    .I1_0_0(n187_I1_0_0),
    .I1_0_1(n187_I1_0_1),
    .I1_1_0(n187_I1_1_0),
    .I1_1_1(n187_I1_1_1),
    .I1_2_0(n187_I1_2_0),
    .I1_2_1(n187_I1_2_1),
    .I1_3_0(n187_I1_3_0),
    .I1_3_1(n187_I1_3_1),
    .O_0_0_0(n187_O_0_0_0),
    .O_0_0_1(n187_O_0_0_1),
    .O_0_1_0(n187_O_0_1_0),
    .O_0_1_1(n187_O_0_1_1),
    .O_1_0_0(n187_O_1_0_0),
    .O_1_0_1(n187_O_1_0_1),
    .O_1_1_0(n187_O_1_1_0),
    .O_1_1_1(n187_O_1_1_1),
    .O_2_0_0(n187_O_2_0_0),
    .O_2_0_1(n187_O_2_0_1),
    .O_2_1_0(n187_O_2_1_0),
    .O_2_1_1(n187_O_2_1_1),
    .O_3_0_0(n187_O_3_0_0),
    .O_3_0_1(n187_O_3_0_1),
    .O_3_1_0(n187_O_3_1_0),
    .O_3_1_1(n187_O_3_1_1)
  );
  MapT_13 n196 ( // @[Top.scala 200:22]
    .valid_up(n196_valid_up),
    .valid_down(n196_valid_down),
    .I_0_0_0(n196_I_0_0_0),
    .I_0_0_1(n196_I_0_0_1),
    .I_0_1_0(n196_I_0_1_0),
    .I_0_1_1(n196_I_0_1_1),
    .I_1_0_0(n196_I_1_0_0),
    .I_1_0_1(n196_I_1_0_1),
    .I_1_1_0(n196_I_1_1_0),
    .I_1_1_1(n196_I_1_1_1),
    .I_2_0_0(n196_I_2_0_0),
    .I_2_0_1(n196_I_2_0_1),
    .I_2_1_0(n196_I_2_1_0),
    .I_2_1_1(n196_I_2_1_1),
    .I_3_0_0(n196_I_3_0_0),
    .I_3_0_1(n196_I_3_0_1),
    .I_3_1_0(n196_I_3_1_0),
    .I_3_1_1(n196_I_3_1_1),
    .O_0_0_0_0(n196_O_0_0_0_0),
    .O_0_0_0_1(n196_O_0_0_0_1),
    .O_0_0_1_0(n196_O_0_0_1_0),
    .O_0_0_1_1(n196_O_0_0_1_1),
    .O_1_0_0_0(n196_O_1_0_0_0),
    .O_1_0_0_1(n196_O_1_0_0_1),
    .O_1_0_1_0(n196_O_1_0_1_0),
    .O_1_0_1_1(n196_O_1_0_1_1),
    .O_2_0_0_0(n196_O_2_0_0_0),
    .O_2_0_0_1(n196_O_2_0_0_1),
    .O_2_0_1_0(n196_O_2_0_1_0),
    .O_2_0_1_1(n196_O_2_0_1_1),
    .O_3_0_0_0(n196_O_3_0_0_0),
    .O_3_0_0_1(n196_O_3_0_0_1),
    .O_3_0_1_0(n196_O_3_0_1_0),
    .O_3_0_1_1(n196_O_3_0_1_1)
  );
  MapT_14 n203 ( // @[Top.scala 203:22]
    .valid_up(n203_valid_up),
    .valid_down(n203_valid_down),
    .I_0_0_0_0(n203_I_0_0_0_0),
    .I_0_0_0_1(n203_I_0_0_0_1),
    .I_0_0_1_0(n203_I_0_0_1_0),
    .I_0_0_1_1(n203_I_0_0_1_1),
    .I_1_0_0_0(n203_I_1_0_0_0),
    .I_1_0_0_1(n203_I_1_0_0_1),
    .I_1_0_1_0(n203_I_1_0_1_0),
    .I_1_0_1_1(n203_I_1_0_1_1),
    .I_2_0_0_0(n203_I_2_0_0_0),
    .I_2_0_0_1(n203_I_2_0_0_1),
    .I_2_0_1_0(n203_I_2_0_1_0),
    .I_2_0_1_1(n203_I_2_0_1_1),
    .I_3_0_0_0(n203_I_3_0_0_0),
    .I_3_0_0_1(n203_I_3_0_0_1),
    .I_3_0_1_0(n203_I_3_0_1_0),
    .I_3_0_1_1(n203_I_3_0_1_1),
    .O_0_0_0(n203_O_0_0_0),
    .O_0_0_1(n203_O_0_0_1),
    .O_0_1_0(n203_O_0_1_0),
    .O_0_1_1(n203_O_0_1_1),
    .O_1_0_0(n203_O_1_0_0),
    .O_1_0_1(n203_O_1_0_1),
    .O_1_1_0(n203_O_1_1_0),
    .O_1_1_1(n203_O_1_1_1),
    .O_2_0_0(n203_O_2_0_0),
    .O_2_0_1(n203_O_2_0_1),
    .O_2_1_0(n203_O_2_1_0),
    .O_2_1_1(n203_O_2_1_1),
    .O_3_0_0(n203_O_3_0_0),
    .O_3_0_1(n203_O_3_0_1),
    .O_3_1_0(n203_O_3_1_0),
    .O_3_1_1(n203_O_3_1_1)
  );
  MapT_15 n245 ( // @[Top.scala 206:22]
    .clock(n245_clock),
    .reset(n245_reset),
    .valid_up(n245_valid_up),
    .valid_down(n245_valid_down),
    .I_0_0_0(n245_I_0_0_0),
    .I_0_0_1(n245_I_0_0_1),
    .I_0_1_0(n245_I_0_1_0),
    .I_0_1_1(n245_I_0_1_1),
    .I_1_0_0(n245_I_1_0_0),
    .I_1_0_1(n245_I_1_0_1),
    .I_1_1_0(n245_I_1_1_0),
    .I_1_1_1(n245_I_1_1_1),
    .I_2_0_0(n245_I_2_0_0),
    .I_2_0_1(n245_I_2_0_1),
    .I_2_1_0(n245_I_2_1_0),
    .I_2_1_1(n245_I_2_1_1),
    .I_3_0_0(n245_I_3_0_0),
    .I_3_0_1(n245_I_3_0_1),
    .I_3_1_0(n245_I_3_1_0),
    .I_3_1_1(n245_I_3_1_1),
    .O_0_0_0(n245_O_0_0_0),
    .O_1_0_0(n245_O_1_0_0),
    .O_2_0_0(n245_O_2_0_0),
    .O_3_0_0(n245_O_3_0_0)
  );
  Passthrough n246 ( // @[Top.scala 209:22]
    .valid_up(n246_valid_up),
    .valid_down(n246_valid_down),
    .I_0_0_0(n246_I_0_0_0),
    .I_1_0_0(n246_I_1_0_0),
    .I_2_0_0(n246_I_2_0_0),
    .I_3_0_0(n246_I_3_0_0),
    .O_0_0(n246_O_0_0),
    .O_1_0(n246_O_1_0),
    .O_2_0(n246_O_2_0),
    .O_3_0(n246_O_3_0)
  );
  Passthrough_1 n247 ( // @[Top.scala 212:22]
    .valid_up(n247_valid_up),
    .valid_down(n247_valid_down),
    .I_0_0(n247_I_0_0),
    .I_1_0(n247_I_1_0),
    .I_2_0(n247_I_2_0),
    .I_3_0(n247_I_3_0),
    .O_0(n247_O_0),
    .O_1(n247_O_1),
    .O_2(n247_O_2),
    .O_3(n247_O_3)
  );
  FIFO n248 ( // @[Top.scala 215:22]
    .clock(n248_clock),
    .reset(n248_reset),
    .valid_up(n248_valid_up),
    .valid_down(n248_valid_down),
    .I_0(n248_I_0),
    .I_1(n248_I_1),
    .I_2(n248_I_2),
    .I_3(n248_I_3),
    .O_0(n248_O_0),
    .O_1(n248_O_1),
    .O_2(n248_O_2),
    .O_3(n248_O_3)
  );
  FIFO n249 ( // @[Top.scala 218:22]
    .clock(n249_clock),
    .reset(n249_reset),
    .valid_up(n249_valid_up),
    .valid_down(n249_valid_down),
    .I_0(n249_I_0),
    .I_1(n249_I_1),
    .I_2(n249_I_2),
    .I_3(n249_I_3),
    .O_0(n249_O_0),
    .O_1(n249_O_1),
    .O_2(n249_O_2),
    .O_3(n249_O_3)
  );
  FIFO n250 ( // @[Top.scala 221:22]
    .clock(n250_clock),
    .reset(n250_reset),
    .valid_up(n250_valid_up),
    .valid_down(n250_valid_down),
    .I_0(n250_I_0),
    .I_1(n250_I_1),
    .I_2(n250_I_2),
    .I_3(n250_I_3),
    .O_0(n250_O_0),
    .O_1(n250_O_1),
    .O_2(n250_O_2),
    .O_3(n250_O_3)
  );
  assign valid_down = n250_valid_down; // @[Top.scala 225:16]
  assign O_0 = n250_O_0; // @[Top.scala 224:7]
  assign O_1 = n250_O_1; // @[Top.scala 224:7]
  assign O_2 = n250_O_2; // @[Top.scala 224:7]
  assign O_3 = n250_O_3; // @[Top.scala 224:7]
  assign n1_clock = clock;
  assign n1_reset = reset;
  assign n1_valid_up = valid_up; // @[Top.scala 77:17]
  assign n1_I_0 = I_0; // @[Top.scala 76:10]
  assign n1_I_1 = I_1; // @[Top.scala 76:10]
  assign n1_I_2 = I_2; // @[Top.scala 76:10]
  assign n1_I_3 = I_3; // @[Top.scala 76:10]
  assign n2_clock = clock;
  assign n2_reset = reset;
  assign n2_valid_up = n1_valid_down; // @[Top.scala 80:17]
  assign n2_I_0 = n1_O_0; // @[Top.scala 79:10]
  assign n2_I_1 = n1_O_1; // @[Top.scala 79:10]
  assign n2_I_2 = n1_O_2; // @[Top.scala 79:10]
  assign n2_I_3 = n1_O_3; // @[Top.scala 79:10]
  assign n3_clock = clock;
  assign n3_reset = reset;
  assign n3_valid_up = n2_valid_down; // @[Top.scala 83:17]
  assign n3_I_0 = n2_O_0; // @[Top.scala 82:10]
  assign n3_I_1 = n2_O_1; // @[Top.scala 82:10]
  assign n3_I_2 = n2_O_2; // @[Top.scala 82:10]
  assign n3_I_3 = n2_O_3; // @[Top.scala 82:10]
  assign n4_clock = clock;
  assign n4_valid_up = n3_valid_down; // @[Top.scala 86:17]
  assign n4_I_0 = n3_O_0; // @[Top.scala 85:10]
  assign n4_I_1 = n3_O_1; // @[Top.scala 85:10]
  assign n4_I_2 = n3_O_2; // @[Top.scala 85:10]
  assign n4_I_3 = n3_O_3; // @[Top.scala 85:10]
  assign n5_clock = clock;
  assign n5_valid_up = n4_valid_down; // @[Top.scala 89:17]
  assign n5_I_0 = n4_O_0; // @[Top.scala 88:10]
  assign n5_I_1 = n4_O_1; // @[Top.scala 88:10]
  assign n5_I_2 = n4_O_2; // @[Top.scala 88:10]
  assign n5_I_3 = n4_O_3; // @[Top.scala 88:10]
  assign n6_valid_up = n5_valid_down & n4_valid_down; // @[Top.scala 93:17]
  assign n6_I0_0 = n5_O_0; // @[Top.scala 91:11]
  assign n6_I0_1 = n5_O_1; // @[Top.scala 91:11]
  assign n6_I0_2 = n5_O_2; // @[Top.scala 91:11]
  assign n6_I0_3 = n5_O_3; // @[Top.scala 91:11]
  assign n6_I1_0 = n4_O_0; // @[Top.scala 92:11]
  assign n6_I1_1 = n4_O_1; // @[Top.scala 92:11]
  assign n6_I1_2 = n4_O_2; // @[Top.scala 92:11]
  assign n6_I1_3 = n4_O_3; // @[Top.scala 92:11]
  assign n13_valid_up = n6_valid_down & n3_valid_down; // @[Top.scala 97:18]
  assign n13_I0_0_0 = n6_O_0_0; // @[Top.scala 95:12]
  assign n13_I0_0_1 = n6_O_0_1; // @[Top.scala 95:12]
  assign n13_I0_1_0 = n6_O_1_0; // @[Top.scala 95:12]
  assign n13_I0_1_1 = n6_O_1_1; // @[Top.scala 95:12]
  assign n13_I0_2_0 = n6_O_2_0; // @[Top.scala 95:12]
  assign n13_I0_2_1 = n6_O_2_1; // @[Top.scala 95:12]
  assign n13_I0_3_0 = n6_O_3_0; // @[Top.scala 95:12]
  assign n13_I0_3_1 = n6_O_3_1; // @[Top.scala 95:12]
  assign n13_I1_0 = n3_O_0; // @[Top.scala 96:12]
  assign n13_I1_1 = n3_O_1; // @[Top.scala 96:12]
  assign n13_I1_2 = n3_O_2; // @[Top.scala 96:12]
  assign n13_I1_3 = n3_O_3; // @[Top.scala 96:12]
  assign n22_valid_up = n13_valid_down; // @[Top.scala 100:18]
  assign n22_I_0_0 = n13_O_0_0; // @[Top.scala 99:11]
  assign n22_I_0_1 = n13_O_0_1; // @[Top.scala 99:11]
  assign n22_I_0_2 = n13_O_0_2; // @[Top.scala 99:11]
  assign n22_I_1_0 = n13_O_1_0; // @[Top.scala 99:11]
  assign n22_I_1_1 = n13_O_1_1; // @[Top.scala 99:11]
  assign n22_I_1_2 = n13_O_1_2; // @[Top.scala 99:11]
  assign n22_I_2_0 = n13_O_2_0; // @[Top.scala 99:11]
  assign n22_I_2_1 = n13_O_2_1; // @[Top.scala 99:11]
  assign n22_I_2_2 = n13_O_2_2; // @[Top.scala 99:11]
  assign n22_I_3_0 = n13_O_3_0; // @[Top.scala 99:11]
  assign n22_I_3_1 = n13_O_3_1; // @[Top.scala 99:11]
  assign n22_I_3_2 = n13_O_3_2; // @[Top.scala 99:11]
  assign n29_valid_up = n22_valid_down; // @[Top.scala 103:18]
  assign n29_I_0_0_0 = n22_O_0_0_0; // @[Top.scala 102:11]
  assign n29_I_0_0_1 = n22_O_0_0_1; // @[Top.scala 102:11]
  assign n29_I_0_0_2 = n22_O_0_0_2; // @[Top.scala 102:11]
  assign n29_I_1_0_0 = n22_O_1_0_0; // @[Top.scala 102:11]
  assign n29_I_1_0_1 = n22_O_1_0_1; // @[Top.scala 102:11]
  assign n29_I_1_0_2 = n22_O_1_0_2; // @[Top.scala 102:11]
  assign n29_I_2_0_0 = n22_O_2_0_0; // @[Top.scala 102:11]
  assign n29_I_2_0_1 = n22_O_2_0_1; // @[Top.scala 102:11]
  assign n29_I_2_0_2 = n22_O_2_0_2; // @[Top.scala 102:11]
  assign n29_I_3_0_0 = n22_O_3_0_0; // @[Top.scala 102:11]
  assign n29_I_3_0_1 = n22_O_3_0_1; // @[Top.scala 102:11]
  assign n29_I_3_0_2 = n22_O_3_0_2; // @[Top.scala 102:11]
  assign n30_clock = clock;
  assign n30_valid_up = n2_valid_down; // @[Top.scala 106:18]
  assign n30_I_0 = n2_O_0; // @[Top.scala 105:11]
  assign n30_I_1 = n2_O_1; // @[Top.scala 105:11]
  assign n30_I_2 = n2_O_2; // @[Top.scala 105:11]
  assign n30_I_3 = n2_O_3; // @[Top.scala 105:11]
  assign n31_clock = clock;
  assign n31_valid_up = n30_valid_down; // @[Top.scala 109:18]
  assign n31_I_0 = n30_O_0; // @[Top.scala 108:11]
  assign n31_I_1 = n30_O_1; // @[Top.scala 108:11]
  assign n31_I_2 = n30_O_2; // @[Top.scala 108:11]
  assign n31_I_3 = n30_O_3; // @[Top.scala 108:11]
  assign n32_valid_up = n31_valid_down & n30_valid_down; // @[Top.scala 113:18]
  assign n32_I0_0 = n31_O_0; // @[Top.scala 111:12]
  assign n32_I0_1 = n31_O_1; // @[Top.scala 111:12]
  assign n32_I0_2 = n31_O_2; // @[Top.scala 111:12]
  assign n32_I0_3 = n31_O_3; // @[Top.scala 111:12]
  assign n32_I1_0 = n30_O_0; // @[Top.scala 112:12]
  assign n32_I1_1 = n30_O_1; // @[Top.scala 112:12]
  assign n32_I1_2 = n30_O_2; // @[Top.scala 112:12]
  assign n32_I1_3 = n30_O_3; // @[Top.scala 112:12]
  assign n39_valid_up = n32_valid_down & n2_valid_down; // @[Top.scala 117:18]
  assign n39_I0_0_0 = n32_O_0_0; // @[Top.scala 115:12]
  assign n39_I0_0_1 = n32_O_0_1; // @[Top.scala 115:12]
  assign n39_I0_1_0 = n32_O_1_0; // @[Top.scala 115:12]
  assign n39_I0_1_1 = n32_O_1_1; // @[Top.scala 115:12]
  assign n39_I0_2_0 = n32_O_2_0; // @[Top.scala 115:12]
  assign n39_I0_2_1 = n32_O_2_1; // @[Top.scala 115:12]
  assign n39_I0_3_0 = n32_O_3_0; // @[Top.scala 115:12]
  assign n39_I0_3_1 = n32_O_3_1; // @[Top.scala 115:12]
  assign n39_I1_0 = n2_O_0; // @[Top.scala 116:12]
  assign n39_I1_1 = n2_O_1; // @[Top.scala 116:12]
  assign n39_I1_2 = n2_O_2; // @[Top.scala 116:12]
  assign n39_I1_3 = n2_O_3; // @[Top.scala 116:12]
  assign n48_valid_up = n39_valid_down; // @[Top.scala 120:18]
  assign n48_I_0_0 = n39_O_0_0; // @[Top.scala 119:11]
  assign n48_I_0_1 = n39_O_0_1; // @[Top.scala 119:11]
  assign n48_I_0_2 = n39_O_0_2; // @[Top.scala 119:11]
  assign n48_I_1_0 = n39_O_1_0; // @[Top.scala 119:11]
  assign n48_I_1_1 = n39_O_1_1; // @[Top.scala 119:11]
  assign n48_I_1_2 = n39_O_1_2; // @[Top.scala 119:11]
  assign n48_I_2_0 = n39_O_2_0; // @[Top.scala 119:11]
  assign n48_I_2_1 = n39_O_2_1; // @[Top.scala 119:11]
  assign n48_I_2_2 = n39_O_2_2; // @[Top.scala 119:11]
  assign n48_I_3_0 = n39_O_3_0; // @[Top.scala 119:11]
  assign n48_I_3_1 = n39_O_3_1; // @[Top.scala 119:11]
  assign n48_I_3_2 = n39_O_3_2; // @[Top.scala 119:11]
  assign n55_valid_up = n48_valid_down; // @[Top.scala 123:18]
  assign n55_I_0_0_0 = n48_O_0_0_0; // @[Top.scala 122:11]
  assign n55_I_0_0_1 = n48_O_0_0_1; // @[Top.scala 122:11]
  assign n55_I_0_0_2 = n48_O_0_0_2; // @[Top.scala 122:11]
  assign n55_I_1_0_0 = n48_O_1_0_0; // @[Top.scala 122:11]
  assign n55_I_1_0_1 = n48_O_1_0_1; // @[Top.scala 122:11]
  assign n55_I_1_0_2 = n48_O_1_0_2; // @[Top.scala 122:11]
  assign n55_I_2_0_0 = n48_O_2_0_0; // @[Top.scala 122:11]
  assign n55_I_2_0_1 = n48_O_2_0_1; // @[Top.scala 122:11]
  assign n55_I_2_0_2 = n48_O_2_0_2; // @[Top.scala 122:11]
  assign n55_I_3_0_0 = n48_O_3_0_0; // @[Top.scala 122:11]
  assign n55_I_3_0_1 = n48_O_3_0_1; // @[Top.scala 122:11]
  assign n55_I_3_0_2 = n48_O_3_0_2; // @[Top.scala 122:11]
  assign n56_valid_up = n29_valid_down & n55_valid_down; // @[Top.scala 127:18]
  assign n56_I0_0_0 = n29_O_0_0; // @[Top.scala 125:12]
  assign n56_I0_0_1 = n29_O_0_1; // @[Top.scala 125:12]
  assign n56_I0_0_2 = n29_O_0_2; // @[Top.scala 125:12]
  assign n56_I0_1_0 = n29_O_1_0; // @[Top.scala 125:12]
  assign n56_I0_1_1 = n29_O_1_1; // @[Top.scala 125:12]
  assign n56_I0_1_2 = n29_O_1_2; // @[Top.scala 125:12]
  assign n56_I0_2_0 = n29_O_2_0; // @[Top.scala 125:12]
  assign n56_I0_2_1 = n29_O_2_1; // @[Top.scala 125:12]
  assign n56_I0_2_2 = n29_O_2_2; // @[Top.scala 125:12]
  assign n56_I0_3_0 = n29_O_3_0; // @[Top.scala 125:12]
  assign n56_I0_3_1 = n29_O_3_1; // @[Top.scala 125:12]
  assign n56_I0_3_2 = n29_O_3_2; // @[Top.scala 125:12]
  assign n56_I1_0_0 = n55_O_0_0; // @[Top.scala 126:12]
  assign n56_I1_0_1 = n55_O_0_1; // @[Top.scala 126:12]
  assign n56_I1_0_2 = n55_O_0_2; // @[Top.scala 126:12]
  assign n56_I1_1_0 = n55_O_1_0; // @[Top.scala 126:12]
  assign n56_I1_1_1 = n55_O_1_1; // @[Top.scala 126:12]
  assign n56_I1_1_2 = n55_O_1_2; // @[Top.scala 126:12]
  assign n56_I1_2_0 = n55_O_2_0; // @[Top.scala 126:12]
  assign n56_I1_2_1 = n55_O_2_1; // @[Top.scala 126:12]
  assign n56_I1_2_2 = n55_O_2_2; // @[Top.scala 126:12]
  assign n56_I1_3_0 = n55_O_3_0; // @[Top.scala 126:12]
  assign n56_I1_3_1 = n55_O_3_1; // @[Top.scala 126:12]
  assign n56_I1_3_2 = n55_O_3_2; // @[Top.scala 126:12]
  assign n63_clock = clock;
  assign n63_valid_up = n1_valid_down; // @[Top.scala 130:18]
  assign n63_I_0 = n1_O_0; // @[Top.scala 129:11]
  assign n63_I_1 = n1_O_1; // @[Top.scala 129:11]
  assign n63_I_2 = n1_O_2; // @[Top.scala 129:11]
  assign n63_I_3 = n1_O_3; // @[Top.scala 129:11]
  assign n64_clock = clock;
  assign n64_valid_up = n63_valid_down; // @[Top.scala 133:18]
  assign n64_I_0 = n63_O_0; // @[Top.scala 132:11]
  assign n64_I_1 = n63_O_1; // @[Top.scala 132:11]
  assign n64_I_2 = n63_O_2; // @[Top.scala 132:11]
  assign n64_I_3 = n63_O_3; // @[Top.scala 132:11]
  assign n65_valid_up = n64_valid_down & n63_valid_down; // @[Top.scala 137:18]
  assign n65_I0_0 = n64_O_0; // @[Top.scala 135:12]
  assign n65_I0_1 = n64_O_1; // @[Top.scala 135:12]
  assign n65_I0_2 = n64_O_2; // @[Top.scala 135:12]
  assign n65_I0_3 = n64_O_3; // @[Top.scala 135:12]
  assign n65_I1_0 = n63_O_0; // @[Top.scala 136:12]
  assign n65_I1_1 = n63_O_1; // @[Top.scala 136:12]
  assign n65_I1_2 = n63_O_2; // @[Top.scala 136:12]
  assign n65_I1_3 = n63_O_3; // @[Top.scala 136:12]
  assign n72_valid_up = n65_valid_down & n1_valid_down; // @[Top.scala 141:18]
  assign n72_I0_0_0 = n65_O_0_0; // @[Top.scala 139:12]
  assign n72_I0_0_1 = n65_O_0_1; // @[Top.scala 139:12]
  assign n72_I0_1_0 = n65_O_1_0; // @[Top.scala 139:12]
  assign n72_I0_1_1 = n65_O_1_1; // @[Top.scala 139:12]
  assign n72_I0_2_0 = n65_O_2_0; // @[Top.scala 139:12]
  assign n72_I0_2_1 = n65_O_2_1; // @[Top.scala 139:12]
  assign n72_I0_3_0 = n65_O_3_0; // @[Top.scala 139:12]
  assign n72_I0_3_1 = n65_O_3_1; // @[Top.scala 139:12]
  assign n72_I1_0 = n1_O_0; // @[Top.scala 140:12]
  assign n72_I1_1 = n1_O_1; // @[Top.scala 140:12]
  assign n72_I1_2 = n1_O_2; // @[Top.scala 140:12]
  assign n72_I1_3 = n1_O_3; // @[Top.scala 140:12]
  assign n81_valid_up = n72_valid_down; // @[Top.scala 144:18]
  assign n81_I_0_0 = n72_O_0_0; // @[Top.scala 143:11]
  assign n81_I_0_1 = n72_O_0_1; // @[Top.scala 143:11]
  assign n81_I_0_2 = n72_O_0_2; // @[Top.scala 143:11]
  assign n81_I_1_0 = n72_O_1_0; // @[Top.scala 143:11]
  assign n81_I_1_1 = n72_O_1_1; // @[Top.scala 143:11]
  assign n81_I_1_2 = n72_O_1_2; // @[Top.scala 143:11]
  assign n81_I_2_0 = n72_O_2_0; // @[Top.scala 143:11]
  assign n81_I_2_1 = n72_O_2_1; // @[Top.scala 143:11]
  assign n81_I_2_2 = n72_O_2_2; // @[Top.scala 143:11]
  assign n81_I_3_0 = n72_O_3_0; // @[Top.scala 143:11]
  assign n81_I_3_1 = n72_O_3_1; // @[Top.scala 143:11]
  assign n81_I_3_2 = n72_O_3_2; // @[Top.scala 143:11]
  assign n88_valid_up = n81_valid_down; // @[Top.scala 147:18]
  assign n88_I_0_0_0 = n81_O_0_0_0; // @[Top.scala 146:11]
  assign n88_I_0_0_1 = n81_O_0_0_1; // @[Top.scala 146:11]
  assign n88_I_0_0_2 = n81_O_0_0_2; // @[Top.scala 146:11]
  assign n88_I_1_0_0 = n81_O_1_0_0; // @[Top.scala 146:11]
  assign n88_I_1_0_1 = n81_O_1_0_1; // @[Top.scala 146:11]
  assign n88_I_1_0_2 = n81_O_1_0_2; // @[Top.scala 146:11]
  assign n88_I_2_0_0 = n81_O_2_0_0; // @[Top.scala 146:11]
  assign n88_I_2_0_1 = n81_O_2_0_1; // @[Top.scala 146:11]
  assign n88_I_2_0_2 = n81_O_2_0_2; // @[Top.scala 146:11]
  assign n88_I_3_0_0 = n81_O_3_0_0; // @[Top.scala 146:11]
  assign n88_I_3_0_1 = n81_O_3_0_1; // @[Top.scala 146:11]
  assign n88_I_3_0_2 = n81_O_3_0_2; // @[Top.scala 146:11]
  assign n89_valid_up = n56_valid_down & n88_valid_down; // @[Top.scala 151:18]
  assign n89_I0_0_0_0 = n56_O_0_0_0; // @[Top.scala 149:12]
  assign n89_I0_0_0_1 = n56_O_0_0_1; // @[Top.scala 149:12]
  assign n89_I0_0_0_2 = n56_O_0_0_2; // @[Top.scala 149:12]
  assign n89_I0_0_1_0 = n56_O_0_1_0; // @[Top.scala 149:12]
  assign n89_I0_0_1_1 = n56_O_0_1_1; // @[Top.scala 149:12]
  assign n89_I0_0_1_2 = n56_O_0_1_2; // @[Top.scala 149:12]
  assign n89_I0_1_0_0 = n56_O_1_0_0; // @[Top.scala 149:12]
  assign n89_I0_1_0_1 = n56_O_1_0_1; // @[Top.scala 149:12]
  assign n89_I0_1_0_2 = n56_O_1_0_2; // @[Top.scala 149:12]
  assign n89_I0_1_1_0 = n56_O_1_1_0; // @[Top.scala 149:12]
  assign n89_I0_1_1_1 = n56_O_1_1_1; // @[Top.scala 149:12]
  assign n89_I0_1_1_2 = n56_O_1_1_2; // @[Top.scala 149:12]
  assign n89_I0_2_0_0 = n56_O_2_0_0; // @[Top.scala 149:12]
  assign n89_I0_2_0_1 = n56_O_2_0_1; // @[Top.scala 149:12]
  assign n89_I0_2_0_2 = n56_O_2_0_2; // @[Top.scala 149:12]
  assign n89_I0_2_1_0 = n56_O_2_1_0; // @[Top.scala 149:12]
  assign n89_I0_2_1_1 = n56_O_2_1_1; // @[Top.scala 149:12]
  assign n89_I0_2_1_2 = n56_O_2_1_2; // @[Top.scala 149:12]
  assign n89_I0_3_0_0 = n56_O_3_0_0; // @[Top.scala 149:12]
  assign n89_I0_3_0_1 = n56_O_3_0_1; // @[Top.scala 149:12]
  assign n89_I0_3_0_2 = n56_O_3_0_2; // @[Top.scala 149:12]
  assign n89_I0_3_1_0 = n56_O_3_1_0; // @[Top.scala 149:12]
  assign n89_I0_3_1_1 = n56_O_3_1_1; // @[Top.scala 149:12]
  assign n89_I0_3_1_2 = n56_O_3_1_2; // @[Top.scala 149:12]
  assign n89_I1_0_0 = n88_O_0_0; // @[Top.scala 150:12]
  assign n89_I1_0_1 = n88_O_0_1; // @[Top.scala 150:12]
  assign n89_I1_0_2 = n88_O_0_2; // @[Top.scala 150:12]
  assign n89_I1_1_0 = n88_O_1_0; // @[Top.scala 150:12]
  assign n89_I1_1_1 = n88_O_1_1; // @[Top.scala 150:12]
  assign n89_I1_1_2 = n88_O_1_2; // @[Top.scala 150:12]
  assign n89_I1_2_0 = n88_O_2_0; // @[Top.scala 150:12]
  assign n89_I1_2_1 = n88_O_2_1; // @[Top.scala 150:12]
  assign n89_I1_2_2 = n88_O_2_2; // @[Top.scala 150:12]
  assign n89_I1_3_0 = n88_O_3_0; // @[Top.scala 150:12]
  assign n89_I1_3_1 = n88_O_3_1; // @[Top.scala 150:12]
  assign n89_I1_3_2 = n88_O_3_2; // @[Top.scala 150:12]
  assign n98_valid_up = n89_valid_down; // @[Top.scala 154:18]
  assign n98_I_0_0_0 = n89_O_0_0_0; // @[Top.scala 153:11]
  assign n98_I_0_0_1 = n89_O_0_0_1; // @[Top.scala 153:11]
  assign n98_I_0_0_2 = n89_O_0_0_2; // @[Top.scala 153:11]
  assign n98_I_0_1_0 = n89_O_0_1_0; // @[Top.scala 153:11]
  assign n98_I_0_1_1 = n89_O_0_1_1; // @[Top.scala 153:11]
  assign n98_I_0_1_2 = n89_O_0_1_2; // @[Top.scala 153:11]
  assign n98_I_0_2_0 = n89_O_0_2_0; // @[Top.scala 153:11]
  assign n98_I_0_2_1 = n89_O_0_2_1; // @[Top.scala 153:11]
  assign n98_I_0_2_2 = n89_O_0_2_2; // @[Top.scala 153:11]
  assign n98_I_1_0_0 = n89_O_1_0_0; // @[Top.scala 153:11]
  assign n98_I_1_0_1 = n89_O_1_0_1; // @[Top.scala 153:11]
  assign n98_I_1_0_2 = n89_O_1_0_2; // @[Top.scala 153:11]
  assign n98_I_1_1_0 = n89_O_1_1_0; // @[Top.scala 153:11]
  assign n98_I_1_1_1 = n89_O_1_1_1; // @[Top.scala 153:11]
  assign n98_I_1_1_2 = n89_O_1_1_2; // @[Top.scala 153:11]
  assign n98_I_1_2_0 = n89_O_1_2_0; // @[Top.scala 153:11]
  assign n98_I_1_2_1 = n89_O_1_2_1; // @[Top.scala 153:11]
  assign n98_I_1_2_2 = n89_O_1_2_2; // @[Top.scala 153:11]
  assign n98_I_2_0_0 = n89_O_2_0_0; // @[Top.scala 153:11]
  assign n98_I_2_0_1 = n89_O_2_0_1; // @[Top.scala 153:11]
  assign n98_I_2_0_2 = n89_O_2_0_2; // @[Top.scala 153:11]
  assign n98_I_2_1_0 = n89_O_2_1_0; // @[Top.scala 153:11]
  assign n98_I_2_1_1 = n89_O_2_1_1; // @[Top.scala 153:11]
  assign n98_I_2_1_2 = n89_O_2_1_2; // @[Top.scala 153:11]
  assign n98_I_2_2_0 = n89_O_2_2_0; // @[Top.scala 153:11]
  assign n98_I_2_2_1 = n89_O_2_2_1; // @[Top.scala 153:11]
  assign n98_I_2_2_2 = n89_O_2_2_2; // @[Top.scala 153:11]
  assign n98_I_3_0_0 = n89_O_3_0_0; // @[Top.scala 153:11]
  assign n98_I_3_0_1 = n89_O_3_0_1; // @[Top.scala 153:11]
  assign n98_I_3_0_2 = n89_O_3_0_2; // @[Top.scala 153:11]
  assign n98_I_3_1_0 = n89_O_3_1_0; // @[Top.scala 153:11]
  assign n98_I_3_1_1 = n89_O_3_1_1; // @[Top.scala 153:11]
  assign n98_I_3_1_2 = n89_O_3_1_2; // @[Top.scala 153:11]
  assign n98_I_3_2_0 = n89_O_3_2_0; // @[Top.scala 153:11]
  assign n98_I_3_2_1 = n89_O_3_2_1; // @[Top.scala 153:11]
  assign n98_I_3_2_2 = n89_O_3_2_2; // @[Top.scala 153:11]
  assign n105_valid_up = n98_valid_down; // @[Top.scala 157:19]
  assign n105_I_0_0_0_0 = n98_O_0_0_0_0; // @[Top.scala 156:12]
  assign n105_I_0_0_0_1 = n98_O_0_0_0_1; // @[Top.scala 156:12]
  assign n105_I_0_0_0_2 = n98_O_0_0_0_2; // @[Top.scala 156:12]
  assign n105_I_0_0_1_0 = n98_O_0_0_1_0; // @[Top.scala 156:12]
  assign n105_I_0_0_1_1 = n98_O_0_0_1_1; // @[Top.scala 156:12]
  assign n105_I_0_0_1_2 = n98_O_0_0_1_2; // @[Top.scala 156:12]
  assign n105_I_0_0_2_0 = n98_O_0_0_2_0; // @[Top.scala 156:12]
  assign n105_I_0_0_2_1 = n98_O_0_0_2_1; // @[Top.scala 156:12]
  assign n105_I_0_0_2_2 = n98_O_0_0_2_2; // @[Top.scala 156:12]
  assign n105_I_1_0_0_0 = n98_O_1_0_0_0; // @[Top.scala 156:12]
  assign n105_I_1_0_0_1 = n98_O_1_0_0_1; // @[Top.scala 156:12]
  assign n105_I_1_0_0_2 = n98_O_1_0_0_2; // @[Top.scala 156:12]
  assign n105_I_1_0_1_0 = n98_O_1_0_1_0; // @[Top.scala 156:12]
  assign n105_I_1_0_1_1 = n98_O_1_0_1_1; // @[Top.scala 156:12]
  assign n105_I_1_0_1_2 = n98_O_1_0_1_2; // @[Top.scala 156:12]
  assign n105_I_1_0_2_0 = n98_O_1_0_2_0; // @[Top.scala 156:12]
  assign n105_I_1_0_2_1 = n98_O_1_0_2_1; // @[Top.scala 156:12]
  assign n105_I_1_0_2_2 = n98_O_1_0_2_2; // @[Top.scala 156:12]
  assign n105_I_2_0_0_0 = n98_O_2_0_0_0; // @[Top.scala 156:12]
  assign n105_I_2_0_0_1 = n98_O_2_0_0_1; // @[Top.scala 156:12]
  assign n105_I_2_0_0_2 = n98_O_2_0_0_2; // @[Top.scala 156:12]
  assign n105_I_2_0_1_0 = n98_O_2_0_1_0; // @[Top.scala 156:12]
  assign n105_I_2_0_1_1 = n98_O_2_0_1_1; // @[Top.scala 156:12]
  assign n105_I_2_0_1_2 = n98_O_2_0_1_2; // @[Top.scala 156:12]
  assign n105_I_2_0_2_0 = n98_O_2_0_2_0; // @[Top.scala 156:12]
  assign n105_I_2_0_2_1 = n98_O_2_0_2_1; // @[Top.scala 156:12]
  assign n105_I_2_0_2_2 = n98_O_2_0_2_2; // @[Top.scala 156:12]
  assign n105_I_3_0_0_0 = n98_O_3_0_0_0; // @[Top.scala 156:12]
  assign n105_I_3_0_0_1 = n98_O_3_0_0_1; // @[Top.scala 156:12]
  assign n105_I_3_0_0_2 = n98_O_3_0_0_2; // @[Top.scala 156:12]
  assign n105_I_3_0_1_0 = n98_O_3_0_1_0; // @[Top.scala 156:12]
  assign n105_I_3_0_1_1 = n98_O_3_0_1_1; // @[Top.scala 156:12]
  assign n105_I_3_0_1_2 = n98_O_3_0_1_2; // @[Top.scala 156:12]
  assign n105_I_3_0_2_0 = n98_O_3_0_2_0; // @[Top.scala 156:12]
  assign n105_I_3_0_2_1 = n98_O_3_0_2_1; // @[Top.scala 156:12]
  assign n105_I_3_0_2_2 = n98_O_3_0_2_2; // @[Top.scala 156:12]
  assign n147_clock = clock;
  assign n147_reset = reset;
  assign n147_valid_up = n105_valid_down; // @[Top.scala 160:19]
  assign n147_I_0_0_0 = n105_O_0_0_0; // @[Top.scala 159:12]
  assign n147_I_0_0_1 = n105_O_0_0_1; // @[Top.scala 159:12]
  assign n147_I_0_0_2 = n105_O_0_0_2; // @[Top.scala 159:12]
  assign n147_I_0_1_0 = n105_O_0_1_0; // @[Top.scala 159:12]
  assign n147_I_0_1_1 = n105_O_0_1_1; // @[Top.scala 159:12]
  assign n147_I_0_1_2 = n105_O_0_1_2; // @[Top.scala 159:12]
  assign n147_I_0_2_0 = n105_O_0_2_0; // @[Top.scala 159:12]
  assign n147_I_0_2_1 = n105_O_0_2_1; // @[Top.scala 159:12]
  assign n147_I_0_2_2 = n105_O_0_2_2; // @[Top.scala 159:12]
  assign n147_I_1_0_0 = n105_O_1_0_0; // @[Top.scala 159:12]
  assign n147_I_1_0_1 = n105_O_1_0_1; // @[Top.scala 159:12]
  assign n147_I_1_0_2 = n105_O_1_0_2; // @[Top.scala 159:12]
  assign n147_I_1_1_0 = n105_O_1_1_0; // @[Top.scala 159:12]
  assign n147_I_1_1_1 = n105_O_1_1_1; // @[Top.scala 159:12]
  assign n147_I_1_1_2 = n105_O_1_1_2; // @[Top.scala 159:12]
  assign n147_I_1_2_0 = n105_O_1_2_0; // @[Top.scala 159:12]
  assign n147_I_1_2_1 = n105_O_1_2_1; // @[Top.scala 159:12]
  assign n147_I_1_2_2 = n105_O_1_2_2; // @[Top.scala 159:12]
  assign n147_I_2_0_0 = n105_O_2_0_0; // @[Top.scala 159:12]
  assign n147_I_2_0_1 = n105_O_2_0_1; // @[Top.scala 159:12]
  assign n147_I_2_0_2 = n105_O_2_0_2; // @[Top.scala 159:12]
  assign n147_I_2_1_0 = n105_O_2_1_0; // @[Top.scala 159:12]
  assign n147_I_2_1_1 = n105_O_2_1_1; // @[Top.scala 159:12]
  assign n147_I_2_1_2 = n105_O_2_1_2; // @[Top.scala 159:12]
  assign n147_I_2_2_0 = n105_O_2_2_0; // @[Top.scala 159:12]
  assign n147_I_2_2_1 = n105_O_2_2_1; // @[Top.scala 159:12]
  assign n147_I_2_2_2 = n105_O_2_2_2; // @[Top.scala 159:12]
  assign n147_I_3_0_0 = n105_O_3_0_0; // @[Top.scala 159:12]
  assign n147_I_3_0_1 = n105_O_3_0_1; // @[Top.scala 159:12]
  assign n147_I_3_0_2 = n105_O_3_0_2; // @[Top.scala 159:12]
  assign n147_I_3_1_0 = n105_O_3_1_0; // @[Top.scala 159:12]
  assign n147_I_3_1_1 = n105_O_3_1_1; // @[Top.scala 159:12]
  assign n147_I_3_1_2 = n105_O_3_1_2; // @[Top.scala 159:12]
  assign n147_I_3_2_0 = n105_O_3_2_0; // @[Top.scala 159:12]
  assign n147_I_3_2_1 = n105_O_3_2_1; // @[Top.scala 159:12]
  assign n147_I_3_2_2 = n105_O_3_2_2; // @[Top.scala 159:12]
  assign n148_valid_up = n147_valid_down; // @[Top.scala 163:19]
  assign n148_I_0_0_0 = n147_O_0_0_0; // @[Top.scala 162:12]
  assign n148_I_1_0_0 = n147_O_1_0_0; // @[Top.scala 162:12]
  assign n148_I_2_0_0 = n147_O_2_0_0; // @[Top.scala 162:12]
  assign n148_I_3_0_0 = n147_O_3_0_0; // @[Top.scala 162:12]
  assign n149_valid_up = n148_valid_down; // @[Top.scala 166:19]
  assign n149_I_0_0 = n148_O_0_0; // @[Top.scala 165:12]
  assign n149_I_1_0 = n148_O_1_0; // @[Top.scala 165:12]
  assign n149_I_2_0 = n148_O_2_0; // @[Top.scala 165:12]
  assign n149_I_3_0 = n148_O_3_0; // @[Top.scala 165:12]
  assign n150_clock = clock;
  assign n150_reset = reset;
  assign n150_valid_up = n149_valid_down; // @[Top.scala 169:19]
  assign n150_I_0 = n149_O_0; // @[Top.scala 168:12]
  assign n150_I_1 = n149_O_1; // @[Top.scala 168:12]
  assign n150_I_2 = n149_O_2; // @[Top.scala 168:12]
  assign n150_I_3 = n149_O_3; // @[Top.scala 168:12]
  assign n151_clock = clock;
  assign n151_valid_up = n150_valid_down; // @[Top.scala 172:19]
  assign n151_I_0 = n150_O_0; // @[Top.scala 171:12]
  assign n151_I_1 = n150_O_1; // @[Top.scala 171:12]
  assign n151_I_2 = n150_O_2; // @[Top.scala 171:12]
  assign n151_I_3 = n150_O_3; // @[Top.scala 171:12]
  assign n152_valid_up = n151_valid_down & n150_valid_down; // @[Top.scala 176:19]
  assign n152_I0_0 = n151_O_0; // @[Top.scala 174:13]
  assign n152_I0_1 = n151_O_1; // @[Top.scala 174:13]
  assign n152_I0_2 = n151_O_2; // @[Top.scala 174:13]
  assign n152_I0_3 = n151_O_3; // @[Top.scala 174:13]
  assign n152_I1_0 = n150_O_0; // @[Top.scala 175:13]
  assign n152_I1_1 = n150_O_1; // @[Top.scala 175:13]
  assign n152_I1_2 = n150_O_2; // @[Top.scala 175:13]
  assign n152_I1_3 = n150_O_3; // @[Top.scala 175:13]
  assign n161_valid_up = n152_valid_down; // @[Top.scala 179:19]
  assign n161_I_0_0 = n152_O_0_0; // @[Top.scala 178:12]
  assign n161_I_0_1 = n152_O_0_1; // @[Top.scala 178:12]
  assign n161_I_1_0 = n152_O_1_0; // @[Top.scala 178:12]
  assign n161_I_1_1 = n152_O_1_1; // @[Top.scala 178:12]
  assign n161_I_2_0 = n152_O_2_0; // @[Top.scala 178:12]
  assign n161_I_2_1 = n152_O_2_1; // @[Top.scala 178:12]
  assign n161_I_3_0 = n152_O_3_0; // @[Top.scala 178:12]
  assign n161_I_3_1 = n152_O_3_1; // @[Top.scala 178:12]
  assign n168_valid_up = n161_valid_down; // @[Top.scala 182:19]
  assign n168_I_0_0_0 = n161_O_0_0_0; // @[Top.scala 181:12]
  assign n168_I_0_0_1 = n161_O_0_0_1; // @[Top.scala 181:12]
  assign n168_I_1_0_0 = n161_O_1_0_0; // @[Top.scala 181:12]
  assign n168_I_1_0_1 = n161_O_1_0_1; // @[Top.scala 181:12]
  assign n168_I_2_0_0 = n161_O_2_0_0; // @[Top.scala 181:12]
  assign n168_I_2_0_1 = n161_O_2_0_1; // @[Top.scala 181:12]
  assign n168_I_3_0_0 = n161_O_3_0_0; // @[Top.scala 181:12]
  assign n168_I_3_0_1 = n161_O_3_0_1; // @[Top.scala 181:12]
  assign n169_clock = clock;
  assign n169_valid_up = n149_valid_down; // @[Top.scala 185:19]
  assign n169_I_0 = n149_O_0; // @[Top.scala 184:12]
  assign n169_I_1 = n149_O_1; // @[Top.scala 184:12]
  assign n169_I_2 = n149_O_2; // @[Top.scala 184:12]
  assign n169_I_3 = n149_O_3; // @[Top.scala 184:12]
  assign n170_valid_up = n169_valid_down & n149_valid_down; // @[Top.scala 189:19]
  assign n170_I0_0 = n169_O_0; // @[Top.scala 187:13]
  assign n170_I0_1 = n169_O_1; // @[Top.scala 187:13]
  assign n170_I0_2 = n169_O_2; // @[Top.scala 187:13]
  assign n170_I0_3 = n169_O_3; // @[Top.scala 187:13]
  assign n170_I1_0 = n149_O_0; // @[Top.scala 188:13]
  assign n170_I1_1 = n149_O_1; // @[Top.scala 188:13]
  assign n170_I1_2 = n149_O_2; // @[Top.scala 188:13]
  assign n170_I1_3 = n149_O_3; // @[Top.scala 188:13]
  assign n179_valid_up = n170_valid_down; // @[Top.scala 192:19]
  assign n179_I_0_0 = n170_O_0_0; // @[Top.scala 191:12]
  assign n179_I_0_1 = n170_O_0_1; // @[Top.scala 191:12]
  assign n179_I_1_0 = n170_O_1_0; // @[Top.scala 191:12]
  assign n179_I_1_1 = n170_O_1_1; // @[Top.scala 191:12]
  assign n179_I_2_0 = n170_O_2_0; // @[Top.scala 191:12]
  assign n179_I_2_1 = n170_O_2_1; // @[Top.scala 191:12]
  assign n179_I_3_0 = n170_O_3_0; // @[Top.scala 191:12]
  assign n179_I_3_1 = n170_O_3_1; // @[Top.scala 191:12]
  assign n186_valid_up = n179_valid_down; // @[Top.scala 195:19]
  assign n186_I_0_0_0 = n179_O_0_0_0; // @[Top.scala 194:12]
  assign n186_I_0_0_1 = n179_O_0_0_1; // @[Top.scala 194:12]
  assign n186_I_1_0_0 = n179_O_1_0_0; // @[Top.scala 194:12]
  assign n186_I_1_0_1 = n179_O_1_0_1; // @[Top.scala 194:12]
  assign n186_I_2_0_0 = n179_O_2_0_0; // @[Top.scala 194:12]
  assign n186_I_2_0_1 = n179_O_2_0_1; // @[Top.scala 194:12]
  assign n186_I_3_0_0 = n179_O_3_0_0; // @[Top.scala 194:12]
  assign n186_I_3_0_1 = n179_O_3_0_1; // @[Top.scala 194:12]
  assign n187_valid_up = n168_valid_down & n186_valid_down; // @[Top.scala 199:19]
  assign n187_I0_0_0 = n168_O_0_0; // @[Top.scala 197:13]
  assign n187_I0_0_1 = n168_O_0_1; // @[Top.scala 197:13]
  assign n187_I0_1_0 = n168_O_1_0; // @[Top.scala 197:13]
  assign n187_I0_1_1 = n168_O_1_1; // @[Top.scala 197:13]
  assign n187_I0_2_0 = n168_O_2_0; // @[Top.scala 197:13]
  assign n187_I0_2_1 = n168_O_2_1; // @[Top.scala 197:13]
  assign n187_I0_3_0 = n168_O_3_0; // @[Top.scala 197:13]
  assign n187_I0_3_1 = n168_O_3_1; // @[Top.scala 197:13]
  assign n187_I1_0_0 = n186_O_0_0; // @[Top.scala 198:13]
  assign n187_I1_0_1 = n186_O_0_1; // @[Top.scala 198:13]
  assign n187_I1_1_0 = n186_O_1_0; // @[Top.scala 198:13]
  assign n187_I1_1_1 = n186_O_1_1; // @[Top.scala 198:13]
  assign n187_I1_2_0 = n186_O_2_0; // @[Top.scala 198:13]
  assign n187_I1_2_1 = n186_O_2_1; // @[Top.scala 198:13]
  assign n187_I1_3_0 = n186_O_3_0; // @[Top.scala 198:13]
  assign n187_I1_3_1 = n186_O_3_1; // @[Top.scala 198:13]
  assign n196_valid_up = n187_valid_down; // @[Top.scala 202:19]
  assign n196_I_0_0_0 = n187_O_0_0_0; // @[Top.scala 201:12]
  assign n196_I_0_0_1 = n187_O_0_0_1; // @[Top.scala 201:12]
  assign n196_I_0_1_0 = n187_O_0_1_0; // @[Top.scala 201:12]
  assign n196_I_0_1_1 = n187_O_0_1_1; // @[Top.scala 201:12]
  assign n196_I_1_0_0 = n187_O_1_0_0; // @[Top.scala 201:12]
  assign n196_I_1_0_1 = n187_O_1_0_1; // @[Top.scala 201:12]
  assign n196_I_1_1_0 = n187_O_1_1_0; // @[Top.scala 201:12]
  assign n196_I_1_1_1 = n187_O_1_1_1; // @[Top.scala 201:12]
  assign n196_I_2_0_0 = n187_O_2_0_0; // @[Top.scala 201:12]
  assign n196_I_2_0_1 = n187_O_2_0_1; // @[Top.scala 201:12]
  assign n196_I_2_1_0 = n187_O_2_1_0; // @[Top.scala 201:12]
  assign n196_I_2_1_1 = n187_O_2_1_1; // @[Top.scala 201:12]
  assign n196_I_3_0_0 = n187_O_3_0_0; // @[Top.scala 201:12]
  assign n196_I_3_0_1 = n187_O_3_0_1; // @[Top.scala 201:12]
  assign n196_I_3_1_0 = n187_O_3_1_0; // @[Top.scala 201:12]
  assign n196_I_3_1_1 = n187_O_3_1_1; // @[Top.scala 201:12]
  assign n203_valid_up = n196_valid_down; // @[Top.scala 205:19]
  assign n203_I_0_0_0_0 = n196_O_0_0_0_0; // @[Top.scala 204:12]
  assign n203_I_0_0_0_1 = n196_O_0_0_0_1; // @[Top.scala 204:12]
  assign n203_I_0_0_1_0 = n196_O_0_0_1_0; // @[Top.scala 204:12]
  assign n203_I_0_0_1_1 = n196_O_0_0_1_1; // @[Top.scala 204:12]
  assign n203_I_1_0_0_0 = n196_O_1_0_0_0; // @[Top.scala 204:12]
  assign n203_I_1_0_0_1 = n196_O_1_0_0_1; // @[Top.scala 204:12]
  assign n203_I_1_0_1_0 = n196_O_1_0_1_0; // @[Top.scala 204:12]
  assign n203_I_1_0_1_1 = n196_O_1_0_1_1; // @[Top.scala 204:12]
  assign n203_I_2_0_0_0 = n196_O_2_0_0_0; // @[Top.scala 204:12]
  assign n203_I_2_0_0_1 = n196_O_2_0_0_1; // @[Top.scala 204:12]
  assign n203_I_2_0_1_0 = n196_O_2_0_1_0; // @[Top.scala 204:12]
  assign n203_I_2_0_1_1 = n196_O_2_0_1_1; // @[Top.scala 204:12]
  assign n203_I_3_0_0_0 = n196_O_3_0_0_0; // @[Top.scala 204:12]
  assign n203_I_3_0_0_1 = n196_O_3_0_0_1; // @[Top.scala 204:12]
  assign n203_I_3_0_1_0 = n196_O_3_0_1_0; // @[Top.scala 204:12]
  assign n203_I_3_0_1_1 = n196_O_3_0_1_1; // @[Top.scala 204:12]
  assign n245_clock = clock;
  assign n245_reset = reset;
  assign n245_valid_up = n203_valid_down; // @[Top.scala 208:19]
  assign n245_I_0_0_0 = n203_O_0_0_0; // @[Top.scala 207:12]
  assign n245_I_0_0_1 = n203_O_0_0_1; // @[Top.scala 207:12]
  assign n245_I_0_1_0 = n203_O_0_1_0; // @[Top.scala 207:12]
  assign n245_I_0_1_1 = n203_O_0_1_1; // @[Top.scala 207:12]
  assign n245_I_1_0_0 = n203_O_1_0_0; // @[Top.scala 207:12]
  assign n245_I_1_0_1 = n203_O_1_0_1; // @[Top.scala 207:12]
  assign n245_I_1_1_0 = n203_O_1_1_0; // @[Top.scala 207:12]
  assign n245_I_1_1_1 = n203_O_1_1_1; // @[Top.scala 207:12]
  assign n245_I_2_0_0 = n203_O_2_0_0; // @[Top.scala 207:12]
  assign n245_I_2_0_1 = n203_O_2_0_1; // @[Top.scala 207:12]
  assign n245_I_2_1_0 = n203_O_2_1_0; // @[Top.scala 207:12]
  assign n245_I_2_1_1 = n203_O_2_1_1; // @[Top.scala 207:12]
  assign n245_I_3_0_0 = n203_O_3_0_0; // @[Top.scala 207:12]
  assign n245_I_3_0_1 = n203_O_3_0_1; // @[Top.scala 207:12]
  assign n245_I_3_1_0 = n203_O_3_1_0; // @[Top.scala 207:12]
  assign n245_I_3_1_1 = n203_O_3_1_1; // @[Top.scala 207:12]
  assign n246_valid_up = n245_valid_down; // @[Top.scala 211:19]
  assign n246_I_0_0_0 = n245_O_0_0_0; // @[Top.scala 210:12]
  assign n246_I_1_0_0 = n245_O_1_0_0; // @[Top.scala 210:12]
  assign n246_I_2_0_0 = n245_O_2_0_0; // @[Top.scala 210:12]
  assign n246_I_3_0_0 = n245_O_3_0_0; // @[Top.scala 210:12]
  assign n247_valid_up = n246_valid_down; // @[Top.scala 214:19]
  assign n247_I_0_0 = n246_O_0_0; // @[Top.scala 213:12]
  assign n247_I_1_0 = n246_O_1_0; // @[Top.scala 213:12]
  assign n247_I_2_0 = n246_O_2_0; // @[Top.scala 213:12]
  assign n247_I_3_0 = n246_O_3_0; // @[Top.scala 213:12]
  assign n248_clock = clock;
  assign n248_reset = reset;
  assign n248_valid_up = n247_valid_down; // @[Top.scala 217:19]
  assign n248_I_0 = n247_O_0; // @[Top.scala 216:12]
  assign n248_I_1 = n247_O_1; // @[Top.scala 216:12]
  assign n248_I_2 = n247_O_2; // @[Top.scala 216:12]
  assign n248_I_3 = n247_O_3; // @[Top.scala 216:12]
  assign n249_clock = clock;
  assign n249_reset = reset;
  assign n249_valid_up = n248_valid_down; // @[Top.scala 220:19]
  assign n249_I_0 = n248_O_0; // @[Top.scala 219:12]
  assign n249_I_1 = n248_O_1; // @[Top.scala 219:12]
  assign n249_I_2 = n248_O_2; // @[Top.scala 219:12]
  assign n249_I_3 = n248_O_3; // @[Top.scala 219:12]
  assign n250_clock = clock;
  assign n250_reset = reset;
  assign n250_valid_up = n249_valid_down; // @[Top.scala 223:19]
  assign n250_I_0 = n249_O_0; // @[Top.scala 222:12]
  assign n250_I_1 = n249_O_1; // @[Top.scala 222:12]
  assign n250_I_2 = n249_O_2; // @[Top.scala 222:12]
  assign n250_I_3 = n249_O_3; // @[Top.scala 222:12]
endmodule
