module FIFO(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I,
  output [7:0] O
);
  reg [7:0] _T; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_1;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O = _T; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= I;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module NestedCounters(
  input   CE,
  output  valid
);
  assign valid = CE; // @[NestedCounters.scala 65:13]
endmodule
module NestedCountersWithNumValid(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 20:44]
  wire  NestedCounters_valid; // @[NestedCounters.scala 20:44]
  NestedCounters NestedCounters ( // @[NestedCounters.scala 20:44]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 22:9]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 21:27]
endmodule
module RAM_ST(
  input         clock,
  input         RE,
  input  [10:0] RADDR,
  output [7:0]  RDATA,
  input         WE,
  input  [10:0] WADDR,
  input  [7:0]  WDATA
);
  wire  write_elem_counter_CE; // @[RAM_ST.scala 20:34]
  wire  write_elem_counter_valid; // @[RAM_ST.scala 20:34]
  wire  read_elem_counter_CE; // @[RAM_ST.scala 21:33]
  wire  read_elem_counter_valid; // @[RAM_ST.scala 21:33]
  reg [7:0] ram [0:1919]; // @[RAM_ST.scala 29:24]
  reg [31:0] _RAND_0;
  wire [7:0] ram__T_8_data; // @[RAM_ST.scala 29:24]
  wire [10:0] ram__T_8_addr; // @[RAM_ST.scala 29:24]
  reg [31:0] _RAND_1;
  wire [7:0] ram__T_2_data; // @[RAM_ST.scala 29:24]
  wire [10:0] ram__T_2_addr; // @[RAM_ST.scala 29:24]
  wire  ram__T_2_mask; // @[RAM_ST.scala 29:24]
  wire  ram__T_2_en; // @[RAM_ST.scala 29:24]
  reg  ram__T_8_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [10:0] ram__T_8_addr_pipe_0;
  reg [31:0] _RAND_3;
  wire [10:0] _GEN_1; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_2; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_3; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_4; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_5; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_6; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_7; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_8; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_9; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_10; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_11; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_12; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_13; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_14; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_15; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_16; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_17; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_18; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_19; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_20; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_21; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_22; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_23; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_24; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_25; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_26; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_27; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_28; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_29; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_30; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_31; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_32; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_33; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_34; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_35; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_36; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_37; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_38; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_39; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_40; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_41; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_42; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_43; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_44; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_45; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_46; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_47; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_48; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_49; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_50; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_51; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_52; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_53; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_54; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_55; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_56; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_57; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_58; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_59; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_60; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_61; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_62; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_63; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_64; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_65; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_66; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_67; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_68; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_69; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_70; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_71; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_72; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_73; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_74; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_75; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_76; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_77; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_78; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_79; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_80; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_81; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_82; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_83; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_84; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_85; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_86; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_87; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_88; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_89; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_90; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_91; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_92; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_93; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_94; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_95; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_96; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_97; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_98; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_99; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_100; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_101; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_102; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_103; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_104; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_105; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_106; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_107; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_108; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_109; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_110; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_111; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_112; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_113; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_114; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_115; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_116; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_117; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_118; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_119; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_120; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_121; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_122; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_123; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_124; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_125; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_126; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_127; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_128; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_129; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_130; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_131; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_132; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_133; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_134; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_135; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_136; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_137; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_138; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_139; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_140; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_141; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_142; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_143; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_144; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_145; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_146; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_147; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_148; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_149; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_150; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_151; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_152; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_153; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_154; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_155; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_156; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_157; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_158; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_159; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_160; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_161; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_162; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_163; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_164; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_165; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_166; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_167; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_168; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_169; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_170; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_171; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_172; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_173; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_174; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_175; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_176; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_177; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_178; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_179; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_180; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_181; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_182; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_183; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_184; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_185; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_186; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_187; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_188; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_189; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_190; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_191; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_192; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_193; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_194; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_195; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_196; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_197; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_198; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_199; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_200; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_201; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_202; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_203; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_204; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_205; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_206; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_207; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_208; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_209; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_210; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_211; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_212; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_213; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_214; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_215; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_216; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_217; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_218; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_219; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_220; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_221; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_222; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_223; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_224; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_225; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_226; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_227; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_228; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_229; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_230; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_231; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_232; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_233; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_234; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_235; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_236; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_237; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_238; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_239; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_240; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_241; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_242; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_243; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_244; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_245; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_246; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_247; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_248; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_249; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_250; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_251; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_252; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_253; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_254; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_255; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_256; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_257; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_258; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_259; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_260; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_261; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_262; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_263; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_264; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_265; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_266; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_267; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_268; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_269; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_270; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_271; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_272; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_273; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_274; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_275; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_276; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_277; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_278; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_279; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_280; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_281; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_282; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_283; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_284; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_285; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_286; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_287; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_288; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_289; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_290; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_291; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_292; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_293; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_294; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_295; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_296; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_297; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_298; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_299; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_300; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_301; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_302; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_303; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_304; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_305; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_306; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_307; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_308; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_309; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_310; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_311; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_312; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_313; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_314; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_315; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_316; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_317; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_318; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_319; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_320; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_321; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_322; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_323; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_324; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_325; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_326; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_327; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_328; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_329; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_330; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_331; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_332; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_333; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_334; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_335; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_336; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_337; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_338; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_339; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_340; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_341; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_342; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_343; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_344; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_345; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_346; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_347; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_348; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_349; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_350; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_351; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_352; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_353; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_354; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_355; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_356; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_357; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_358; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_359; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_360; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_361; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_362; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_363; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_364; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_365; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_366; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_367; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_368; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_369; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_370; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_371; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_372; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_373; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_374; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_375; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_376; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_377; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_378; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_379; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_380; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_381; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_382; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_383; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_384; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_385; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_386; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_387; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_388; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_389; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_390; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_391; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_392; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_393; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_394; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_395; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_396; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_397; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_398; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_399; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_400; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_401; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_402; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_403; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_404; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_405; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_406; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_407; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_408; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_409; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_410; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_411; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_412; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_413; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_414; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_415; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_416; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_417; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_418; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_419; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_420; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_421; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_422; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_423; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_424; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_425; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_426; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_427; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_428; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_429; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_430; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_431; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_432; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_433; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_434; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_435; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_436; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_437; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_438; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_439; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_440; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_441; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_442; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_443; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_444; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_445; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_446; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_447; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_448; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_449; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_450; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_451; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_452; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_453; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_454; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_455; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_456; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_457; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_458; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_459; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_460; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_461; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_462; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_463; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_464; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_465; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_466; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_467; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_468; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_469; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_470; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_471; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_472; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_473; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_474; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_475; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_476; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_477; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_478; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_479; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_480; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_481; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_482; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_483; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_484; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_485; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_486; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_487; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_488; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_489; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_490; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_491; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_492; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_493; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_494; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_495; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_496; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_497; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_498; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_499; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_500; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_501; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_502; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_503; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_504; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_505; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_506; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_507; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_508; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_509; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_510; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_511; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_512; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_513; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_514; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_515; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_516; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_517; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_518; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_519; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_520; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_521; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_522; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_523; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_524; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_525; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_526; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_527; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_528; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_529; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_530; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_531; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_532; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_533; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_534; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_535; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_536; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_537; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_538; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_539; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_540; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_541; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_542; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_543; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_544; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_545; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_546; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_547; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_548; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_549; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_550; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_551; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_552; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_553; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_554; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_555; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_556; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_557; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_558; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_559; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_560; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_561; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_562; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_563; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_564; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_565; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_566; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_567; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_568; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_569; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_570; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_571; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_572; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_573; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_574; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_575; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_576; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_577; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_578; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_579; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_580; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_581; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_582; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_583; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_584; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_585; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_586; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_587; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_588; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_589; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_590; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_591; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_592; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_593; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_594; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_595; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_596; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_597; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_598; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_599; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_600; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_601; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_602; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_603; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_604; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_605; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_606; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_607; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_608; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_609; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_610; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_611; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_612; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_613; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_614; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_615; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_616; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_617; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_618; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_619; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_620; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_621; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_622; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_623; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_624; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_625; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_626; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_627; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_628; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_629; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_630; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_631; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_632; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_633; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_634; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_635; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_636; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_637; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_638; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_639; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_640; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_641; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_642; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_643; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_644; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_645; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_646; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_647; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_648; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_649; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_650; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_651; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_652; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_653; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_654; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_655; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_656; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_657; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_658; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_659; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_660; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_661; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_662; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_663; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_664; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_665; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_666; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_667; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_668; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_669; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_670; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_671; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_672; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_673; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_674; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_675; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_676; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_677; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_678; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_679; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_680; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_681; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_682; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_683; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_684; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_685; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_686; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_687; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_688; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_689; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_690; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_691; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_692; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_693; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_694; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_695; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_696; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_697; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_698; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_699; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_700; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_701; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_702; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_703; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_704; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_705; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_706; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_707; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_708; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_709; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_710; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_711; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_712; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_713; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_714; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_715; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_716; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_717; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_718; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_719; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_720; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_721; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_722; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_723; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_724; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_725; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_726; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_727; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_728; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_729; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_730; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_731; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_732; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_733; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_734; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_735; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_736; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_737; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_738; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_739; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_740; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_741; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_742; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_743; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_744; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_745; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_746; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_747; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_748; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_749; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_750; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_751; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_752; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_753; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_754; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_755; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_756; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_757; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_758; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_759; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_760; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_761; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_762; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_763; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_764; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_765; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_766; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_767; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_768; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_769; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_770; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_771; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_772; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_773; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_774; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_775; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_776; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_777; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_778; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_779; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_780; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_781; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_782; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_783; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_784; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_785; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_786; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_787; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_788; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_789; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_790; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_791; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_792; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_793; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_794; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_795; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_796; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_797; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_798; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_799; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_800; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_801; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_802; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_803; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_804; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_805; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_806; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_807; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_808; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_809; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_810; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_811; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_812; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_813; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_814; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_815; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_816; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_817; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_818; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_819; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_820; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_821; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_822; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_823; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_824; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_825; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_826; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_827; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_828; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_829; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_830; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_831; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_832; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_833; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_834; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_835; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_836; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_837; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_838; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_839; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_840; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_841; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_842; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_843; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_844; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_845; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_846; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_847; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_848; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_849; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_850; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_851; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_852; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_853; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_854; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_855; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_856; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_857; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_858; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_859; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_860; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_861; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_862; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_863; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_864; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_865; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_866; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_867; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_868; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_869; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_870; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_871; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_872; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_873; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_874; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_875; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_876; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_877; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_878; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_879; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_880; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_881; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_882; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_883; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_884; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_885; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_886; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_887; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_888; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_889; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_890; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_891; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_892; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_893; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_894; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_895; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_896; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_897; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_898; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_899; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_900; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_901; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_902; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_903; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_904; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_905; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_906; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_907; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_908; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_909; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_910; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_911; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_912; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_913; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_914; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_915; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_916; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_917; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_918; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_919; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_920; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_921; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_922; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_923; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_924; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_925; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_926; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_927; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_928; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_929; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_930; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_931; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_932; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_933; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_934; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_935; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_936; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_937; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_938; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_939; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_940; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_941; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_942; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_943; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_944; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_945; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_946; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_947; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_948; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_949; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_950; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_951; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_952; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_953; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_954; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_955; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_956; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_957; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_958; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_959; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_960; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_961; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_962; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_963; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_964; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_965; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_966; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_967; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_968; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_969; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_970; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_971; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_972; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_973; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_974; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_975; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_976; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_977; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_978; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_979; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_980; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_981; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_982; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_983; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_984; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_985; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_986; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_987; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_988; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_989; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_990; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_991; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_992; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_993; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_994; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_995; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_996; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_997; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_998; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_999; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1000; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1001; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1002; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1003; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1004; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1005; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1006; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1007; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1008; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1009; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1010; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1011; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1012; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1013; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1014; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1015; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1016; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1017; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1018; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1019; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1020; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1021; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1022; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1023; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1024; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1025; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1026; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1027; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1028; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1029; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1030; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1031; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1032; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1033; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1034; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1035; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1036; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1037; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1038; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1039; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1040; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1041; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1042; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1043; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1044; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1045; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1046; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1047; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1048; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1049; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1050; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1051; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1052; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1053; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1054; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1055; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1056; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1057; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1058; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1059; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1060; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1061; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1062; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1063; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1064; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1065; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1066; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1067; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1068; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1069; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1070; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1071; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1072; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1073; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1074; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1075; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1076; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1077; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1078; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1079; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1080; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1081; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1082; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1083; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1084; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1085; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1086; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1087; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1088; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1089; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1090; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1091; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1092; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1093; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1094; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1095; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1096; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1097; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1098; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1099; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1100; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1101; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1102; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1103; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1104; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1105; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1106; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1107; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1108; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1109; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1110; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1111; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1112; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1113; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1114; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1115; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1116; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1117; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1118; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1119; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1120; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1121; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1122; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1123; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1124; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1125; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1126; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1127; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1128; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1129; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1130; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1131; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1132; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1133; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1134; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1135; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1136; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1137; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1138; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1139; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1140; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1141; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1142; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1143; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1144; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1145; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1146; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1147; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1148; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1149; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1150; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1151; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1152; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1153; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1154; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1155; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1156; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1157; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1158; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1159; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1160; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1161; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1162; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1163; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1164; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1165; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1166; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1167; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1168; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1169; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1170; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1171; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1172; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1173; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1174; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1175; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1176; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1177; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1178; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1179; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1180; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1181; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1182; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1183; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1184; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1185; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1186; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1187; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1188; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1189; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1190; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1191; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1192; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1193; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1194; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1195; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1196; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1197; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1198; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1199; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1200; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1201; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1202; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1203; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1204; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1205; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1206; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1207; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1208; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1209; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1210; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1211; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1212; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1213; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1214; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1215; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1216; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1217; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1218; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1219; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1220; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1221; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1222; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1223; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1224; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1225; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1226; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1227; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1228; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1229; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1230; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1231; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1232; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1233; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1234; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1235; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1236; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1237; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1238; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1239; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1240; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1241; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1242; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1243; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1244; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1245; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1246; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1247; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1248; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1249; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1250; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1251; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1252; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1253; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1254; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1255; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1256; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1257; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1258; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1259; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1260; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1261; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1262; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1263; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1264; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1265; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1266; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1267; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1268; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1269; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1270; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1271; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1272; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1273; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1274; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1275; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1276; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1277; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1278; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1279; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1280; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1281; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1282; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1283; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1284; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1285; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1286; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1287; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1288; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1289; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1290; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1291; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1292; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1293; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1294; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1295; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1296; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1297; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1298; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1299; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1300; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1301; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1302; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1303; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1304; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1305; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1306; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1307; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1308; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1309; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1310; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1311; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1312; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1313; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1314; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1315; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1316; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1317; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1318; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1319; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1320; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1321; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1322; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1323; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1324; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1325; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1326; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1327; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1328; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1329; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1330; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1331; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1332; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1333; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1334; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1335; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1336; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1337; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1338; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1339; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1340; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1341; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1342; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1343; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1344; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1345; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1346; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1347; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1348; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1349; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1350; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1351; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1352; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1353; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1354; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1355; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1356; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1357; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1358; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1359; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1360; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1361; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1362; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1363; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1364; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1365; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1366; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1367; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1368; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1369; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1370; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1371; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1372; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1373; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1374; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1375; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1376; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1377; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1378; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1379; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1380; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1381; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1382; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1383; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1384; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1385; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1386; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1387; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1388; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1389; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1390; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1391; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1392; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1393; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1394; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1395; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1396; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1397; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1398; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1399; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1400; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1401; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1402; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1403; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1404; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1405; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1406; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1407; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1408; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1409; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1410; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1411; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1412; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1413; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1414; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1415; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1416; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1417; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1418; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1419; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1420; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1421; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1422; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1423; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1424; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1425; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1426; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1427; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1428; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1429; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1430; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1431; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1432; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1433; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1434; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1435; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1436; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1437; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1438; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1439; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1440; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1441; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1442; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1443; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1444; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1445; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1446; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1447; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1448; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1449; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1450; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1451; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1452; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1453; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1454; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1455; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1456; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1457; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1458; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1459; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1460; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1461; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1462; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1463; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1464; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1465; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1466; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1467; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1468; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1469; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1470; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1471; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1472; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1473; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1474; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1475; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1476; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1477; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1478; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1479; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1480; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1481; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1482; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1483; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1484; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1485; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1486; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1487; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1488; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1489; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1490; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1491; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1492; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1493; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1494; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1495; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1496; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1497; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1498; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1499; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1500; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1501; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1502; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1503; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1504; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1505; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1506; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1507; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1508; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1509; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1510; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1511; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1512; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1513; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1514; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1515; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1516; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1517; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1518; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1519; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1520; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1521; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1522; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1523; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1524; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1525; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1526; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1527; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1528; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1529; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1530; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1531; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1532; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1533; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1534; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1535; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1536; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1537; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1538; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1539; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1540; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1541; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1542; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1543; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1544; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1545; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1546; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1547; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1548; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1549; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1550; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1551; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1552; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1553; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1554; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1555; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1556; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1557; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1558; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1559; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1560; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1561; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1562; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1563; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1564; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1565; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1566; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1567; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1568; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1569; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1570; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1571; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1572; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1573; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1574; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1575; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1576; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1577; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1578; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1579; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1580; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1581; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1582; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1583; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1584; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1585; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1586; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1587; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1588; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1589; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1590; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1591; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1592; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1593; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1594; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1595; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1596; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1597; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1598; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1599; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1600; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1601; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1602; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1603; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1604; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1605; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1606; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1607; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1608; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1609; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1610; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1611; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1612; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1613; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1614; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1615; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1616; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1617; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1618; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1619; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1620; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1621; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1622; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1623; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1624; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1625; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1626; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1627; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1628; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1629; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1630; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1631; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1632; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1633; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1634; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1635; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1636; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1637; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1638; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1639; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1640; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1641; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1642; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1643; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1644; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1645; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1646; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1647; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1648; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1649; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1650; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1651; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1652; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1653; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1654; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1655; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1656; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1657; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1658; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1659; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1660; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1661; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1662; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1663; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1664; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1665; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1666; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1667; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1668; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1669; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1670; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1671; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1672; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1673; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1674; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1675; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1676; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1677; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1678; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1679; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1680; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1681; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1682; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1683; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1684; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1685; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1686; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1687; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1688; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1689; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1690; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1691; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1692; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1693; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1694; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1695; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1696; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1697; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1698; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1699; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1700; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1701; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1702; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1703; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1704; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1705; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1706; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1707; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1708; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1709; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1710; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1711; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1712; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1713; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1714; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1715; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1716; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1717; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1718; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1719; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1720; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1721; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1722; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1723; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1724; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1725; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1726; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1727; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1728; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1729; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1730; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1731; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1732; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1733; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1734; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1735; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1736; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1737; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1738; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1739; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1740; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1741; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1742; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1743; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1744; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1745; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1746; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1747; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1748; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1749; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1750; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1751; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1752; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1753; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1754; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1755; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1756; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1757; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1758; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1759; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1760; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1761; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1762; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1763; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1764; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1765; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1766; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1767; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1768; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1769; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1770; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1771; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1772; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1773; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1774; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1775; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1776; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1777; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1778; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1779; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1780; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1781; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1782; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1783; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1784; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1785; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1786; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1787; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1788; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1789; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1790; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1791; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1792; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1793; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1794; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1795; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1796; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1797; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1798; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1799; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1800; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1801; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1802; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1803; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1804; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1805; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1806; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1807; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1808; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1809; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1810; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1811; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1812; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1813; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1814; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1815; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1816; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1817; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1818; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1819; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1820; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1821; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1822; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1823; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1824; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1825; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1826; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1827; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1828; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1829; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1830; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1831; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1832; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1833; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1834; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1835; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1836; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1837; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1838; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1839; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1840; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1841; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1842; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1843; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1844; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1845; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1846; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1847; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1848; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1849; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1850; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1851; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1852; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1853; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1854; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1855; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1856; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1857; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1858; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1859; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1860; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1861; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1862; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1863; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1864; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1865; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1866; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1867; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1868; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1869; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1870; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1871; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1872; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1873; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1874; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1875; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1876; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1877; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1878; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1879; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1880; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1881; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1882; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1883; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1884; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1885; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1886; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1887; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1888; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1889; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1890; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1891; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1892; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1893; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1894; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1895; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1896; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1897; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1898; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1899; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1900; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1901; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1902; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1903; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1904; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1905; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1906; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1907; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1908; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1909; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1910; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1911; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1912; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1913; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1914; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1915; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1916; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1917; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1918; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1919; // @[RAM_ST.scala 31:71]
  wire [11:0] _T; // @[RAM_ST.scala 31:71]
  wire [10:0] _GEN_1926; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1927; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1928; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1929; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1930; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1931; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1932; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1933; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1934; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1935; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1936; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1937; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1938; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1939; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1940; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1941; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1942; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1943; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1944; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1945; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1946; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1947; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1948; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1949; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1950; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1951; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1952; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1953; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1954; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1955; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1956; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1957; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1958; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1959; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1960; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1961; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1962; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1963; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1964; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1965; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1966; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1967; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1968; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1969; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1970; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1971; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1972; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1973; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1974; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1975; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1976; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1977; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1978; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1979; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1980; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1981; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1982; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1983; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1984; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1985; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1986; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1987; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1988; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1989; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1990; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1991; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1992; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1993; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1994; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1995; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1996; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1997; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1998; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_1999; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2000; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2001; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2002; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2003; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2004; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2005; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2006; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2007; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2008; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2009; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2010; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2011; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2012; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2013; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2014; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2015; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2016; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2017; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2018; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2019; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2020; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2021; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2022; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2023; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2024; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2025; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2026; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2027; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2028; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2029; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2030; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2031; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2032; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2033; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2034; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2035; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2036; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2037; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2038; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2039; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2040; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2041; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2042; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2043; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2044; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2045; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2046; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2047; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2048; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2049; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2050; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2051; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2052; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2053; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2054; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2055; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2056; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2057; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2058; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2059; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2060; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2061; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2062; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2063; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2064; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2065; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2066; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2067; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2068; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2069; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2070; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2071; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2072; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2073; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2074; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2075; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2076; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2077; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2078; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2079; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2080; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2081; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2082; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2083; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2084; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2085; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2086; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2087; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2088; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2089; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2090; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2091; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2092; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2093; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2094; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2095; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2096; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2097; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2098; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2099; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2100; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2101; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2102; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2103; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2104; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2105; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2106; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2107; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2108; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2109; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2110; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2111; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2112; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2113; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2114; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2115; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2116; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2117; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2118; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2119; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2120; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2121; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2122; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2123; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2124; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2125; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2126; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2127; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2128; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2129; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2130; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2131; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2132; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2133; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2134; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2135; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2136; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2137; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2138; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2139; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2140; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2141; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2142; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2143; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2144; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2145; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2146; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2147; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2148; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2149; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2150; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2151; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2152; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2153; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2154; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2155; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2156; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2157; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2158; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2159; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2160; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2161; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2162; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2163; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2164; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2165; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2166; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2167; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2168; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2169; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2170; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2171; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2172; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2173; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2174; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2175; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2176; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2177; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2178; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2179; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2180; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2181; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2182; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2183; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2184; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2185; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2186; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2187; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2188; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2189; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2190; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2191; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2192; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2193; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2194; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2195; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2196; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2197; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2198; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2199; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2200; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2201; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2202; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2203; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2204; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2205; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2206; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2207; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2208; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2209; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2210; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2211; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2212; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2213; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2214; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2215; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2216; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2217; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2218; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2219; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2220; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2221; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2222; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2223; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2224; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2225; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2226; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2227; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2228; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2229; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2230; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2231; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2232; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2233; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2234; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2235; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2236; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2237; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2238; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2239; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2240; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2241; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2242; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2243; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2244; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2245; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2246; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2247; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2248; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2249; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2250; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2251; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2252; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2253; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2254; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2255; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2256; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2257; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2258; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2259; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2260; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2261; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2262; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2263; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2264; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2265; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2266; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2267; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2268; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2269; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2270; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2271; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2272; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2273; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2274; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2275; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2276; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2277; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2278; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2279; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2280; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2281; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2282; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2283; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2284; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2285; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2286; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2287; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2288; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2289; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2290; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2291; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2292; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2293; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2294; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2295; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2296; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2297; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2298; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2299; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2300; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2301; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2302; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2303; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2304; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2305; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2306; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2307; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2308; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2309; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2310; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2311; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2312; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2313; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2314; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2315; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2316; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2317; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2318; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2319; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2320; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2321; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2322; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2323; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2324; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2325; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2326; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2327; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2328; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2329; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2330; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2331; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2332; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2333; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2334; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2335; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2336; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2337; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2338; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2339; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2340; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2341; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2342; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2343; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2344; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2345; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2346; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2347; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2348; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2349; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2350; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2351; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2352; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2353; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2354; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2355; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2356; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2357; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2358; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2359; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2360; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2361; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2362; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2363; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2364; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2365; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2366; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2367; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2368; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2369; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2370; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2371; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2372; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2373; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2374; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2375; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2376; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2377; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2378; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2379; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2380; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2381; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2382; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2383; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2384; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2385; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2386; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2387; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2388; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2389; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2390; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2391; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2392; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2393; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2394; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2395; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2396; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2397; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2398; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2399; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2400; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2401; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2402; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2403; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2404; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2405; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2406; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2407; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2408; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2409; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2410; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2411; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2412; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2413; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2414; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2415; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2416; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2417; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2418; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2419; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2420; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2421; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2422; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2423; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2424; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2425; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2426; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2427; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2428; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2429; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2430; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2431; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2432; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2433; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2434; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2435; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2436; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2437; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2438; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2439; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2440; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2441; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2442; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2443; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2444; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2445; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2446; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2447; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2448; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2449; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2450; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2451; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2452; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2453; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2454; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2455; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2456; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2457; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2458; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2459; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2460; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2461; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2462; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2463; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2464; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2465; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2466; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2467; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2468; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2469; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2470; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2471; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2472; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2473; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2474; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2475; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2476; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2477; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2478; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2479; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2480; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2481; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2482; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2483; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2484; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2485; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2486; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2487; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2488; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2489; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2490; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2491; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2492; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2493; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2494; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2495; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2496; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2497; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2498; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2499; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2500; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2501; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2502; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2503; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2504; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2505; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2506; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2507; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2508; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2509; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2510; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2511; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2512; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2513; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2514; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2515; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2516; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2517; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2518; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2519; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2520; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2521; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2522; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2523; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2524; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2525; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2526; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2527; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2528; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2529; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2530; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2531; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2532; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2533; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2534; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2535; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2536; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2537; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2538; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2539; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2540; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2541; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2542; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2543; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2544; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2545; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2546; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2547; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2548; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2549; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2550; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2551; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2552; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2553; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2554; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2555; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2556; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2557; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2558; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2559; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2560; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2561; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2562; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2563; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2564; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2565; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2566; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2567; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2568; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2569; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2570; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2571; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2572; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2573; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2574; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2575; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2576; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2577; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2578; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2579; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2580; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2581; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2582; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2583; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2584; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2585; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2586; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2587; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2588; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2589; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2590; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2591; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2592; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2593; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2594; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2595; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2596; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2597; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2598; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2599; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2600; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2601; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2602; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2603; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2604; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2605; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2606; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2607; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2608; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2609; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2610; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2611; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2612; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2613; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2614; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2615; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2616; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2617; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2618; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2619; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2620; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2621; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2622; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2623; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2624; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2625; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2626; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2627; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2628; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2629; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2630; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2631; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2632; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2633; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2634; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2635; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2636; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2637; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2638; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2639; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2640; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2641; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2642; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2643; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2644; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2645; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2646; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2647; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2648; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2649; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2650; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2651; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2652; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2653; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2654; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2655; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2656; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2657; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2658; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2659; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2660; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2661; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2662; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2663; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2664; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2665; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2666; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2667; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2668; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2669; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2670; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2671; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2672; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2673; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2674; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2675; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2676; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2677; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2678; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2679; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2680; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2681; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2682; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2683; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2684; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2685; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2686; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2687; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2688; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2689; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2690; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2691; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2692; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2693; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2694; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2695; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2696; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2697; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2698; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2699; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2700; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2701; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2702; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2703; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2704; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2705; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2706; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2707; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2708; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2709; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2710; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2711; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2712; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2713; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2714; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2715; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2716; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2717; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2718; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2719; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2720; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2721; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2722; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2723; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2724; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2725; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2726; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2727; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2728; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2729; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2730; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2731; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2732; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2733; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2734; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2735; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2736; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2737; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2738; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2739; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2740; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2741; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2742; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2743; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2744; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2745; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2746; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2747; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2748; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2749; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2750; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2751; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2752; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2753; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2754; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2755; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2756; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2757; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2758; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2759; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2760; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2761; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2762; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2763; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2764; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2765; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2766; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2767; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2768; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2769; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2770; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2771; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2772; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2773; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2774; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2775; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2776; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2777; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2778; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2779; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2780; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2781; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2782; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2783; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2784; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2785; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2786; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2787; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2788; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2789; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2790; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2791; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2792; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2793; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2794; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2795; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2796; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2797; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2798; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2799; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2800; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2801; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2802; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2803; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2804; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2805; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2806; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2807; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2808; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2809; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2810; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2811; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2812; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2813; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2814; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2815; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2816; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2817; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2818; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2819; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2820; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2821; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2822; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2823; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2824; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2825; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2826; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2827; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2828; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2829; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2830; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2831; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2832; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2833; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2834; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2835; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2836; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2837; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2838; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2839; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2840; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2841; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2842; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2843; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2844; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2845; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2846; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2847; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2848; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2849; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2850; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2851; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2852; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2853; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2854; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2855; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2856; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2857; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2858; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2859; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2860; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2861; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2862; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2863; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2864; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2865; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2866; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2867; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2868; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2869; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2870; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2871; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2872; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2873; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2874; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2875; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2876; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2877; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2878; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2879; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2880; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2881; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2882; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2883; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2884; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2885; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2886; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2887; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2888; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2889; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2890; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2891; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2892; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2893; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2894; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2895; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2896; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2897; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2898; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2899; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2900; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2901; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2902; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2903; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2904; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2905; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2906; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2907; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2908; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2909; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2910; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2911; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2912; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2913; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2914; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2915; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2916; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2917; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2918; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2919; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2920; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2921; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2922; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2923; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2924; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2925; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2926; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2927; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2928; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2929; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2930; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2931; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2932; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2933; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2934; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2935; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2936; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2937; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2938; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2939; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2940; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2941; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2942; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2943; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2944; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2945; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2946; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2947; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2948; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2949; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2950; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2951; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2952; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2953; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2954; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2955; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2956; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2957; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2958; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2959; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2960; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2961; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2962; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2963; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2964; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2965; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2966; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2967; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2968; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2969; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2970; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2971; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2972; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2973; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2974; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2975; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2976; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2977; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2978; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2979; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2980; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2981; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2982; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2983; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2984; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2985; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2986; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2987; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2988; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2989; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2990; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2991; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2992; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2993; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2994; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2995; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2996; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2997; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2998; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_2999; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3000; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3001; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3002; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3003; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3004; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3005; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3006; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3007; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3008; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3009; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3010; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3011; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3012; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3013; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3014; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3015; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3016; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3017; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3018; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3019; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3020; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3021; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3022; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3023; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3024; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3025; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3026; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3027; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3028; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3029; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3030; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3031; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3032; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3033; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3034; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3035; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3036; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3037; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3038; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3039; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3040; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3041; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3042; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3043; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3044; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3045; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3046; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3047; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3048; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3049; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3050; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3051; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3052; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3053; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3054; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3055; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3056; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3057; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3058; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3059; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3060; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3061; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3062; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3063; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3064; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3065; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3066; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3067; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3068; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3069; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3070; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3071; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3072; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3073; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3074; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3075; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3076; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3077; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3078; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3079; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3080; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3081; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3082; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3083; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3084; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3085; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3086; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3087; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3088; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3089; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3090; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3091; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3092; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3093; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3094; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3095; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3096; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3097; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3098; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3099; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3100; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3101; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3102; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3103; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3104; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3105; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3106; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3107; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3108; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3109; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3110; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3111; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3112; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3113; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3114; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3115; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3116; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3117; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3118; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3119; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3120; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3121; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3122; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3123; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3124; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3125; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3126; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3127; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3128; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3129; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3130; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3131; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3132; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3133; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3134; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3135; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3136; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3137; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3138; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3139; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3140; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3141; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3142; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3143; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3144; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3145; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3146; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3147; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3148; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3149; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3150; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3151; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3152; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3153; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3154; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3155; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3156; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3157; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3158; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3159; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3160; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3161; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3162; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3163; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3164; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3165; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3166; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3167; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3168; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3169; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3170; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3171; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3172; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3173; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3174; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3175; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3176; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3177; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3178; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3179; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3180; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3181; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3182; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3183; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3184; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3185; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3186; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3187; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3188; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3189; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3190; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3191; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3192; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3193; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3194; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3195; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3196; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3197; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3198; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3199; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3200; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3201; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3202; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3203; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3204; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3205; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3206; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3207; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3208; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3209; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3210; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3211; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3212; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3213; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3214; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3215; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3216; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3217; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3218; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3219; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3220; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3221; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3222; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3223; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3224; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3225; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3226; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3227; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3228; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3229; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3230; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3231; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3232; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3233; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3234; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3235; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3236; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3237; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3238; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3239; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3240; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3241; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3242; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3243; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3244; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3245; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3246; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3247; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3248; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3249; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3250; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3251; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3252; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3253; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3254; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3255; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3256; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3257; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3258; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3259; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3260; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3261; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3262; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3263; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3264; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3265; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3266; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3267; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3268; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3269; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3270; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3271; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3272; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3273; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3274; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3275; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3276; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3277; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3278; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3279; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3280; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3281; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3282; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3283; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3284; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3285; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3286; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3287; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3288; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3289; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3290; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3291; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3292; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3293; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3294; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3295; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3296; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3297; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3298; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3299; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3300; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3301; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3302; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3303; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3304; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3305; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3306; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3307; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3308; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3309; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3310; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3311; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3312; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3313; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3314; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3315; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3316; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3317; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3318; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3319; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3320; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3321; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3322; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3323; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3324; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3325; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3326; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3327; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3328; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3329; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3330; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3331; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3332; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3333; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3334; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3335; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3336; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3337; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3338; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3339; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3340; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3341; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3342; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3343; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3344; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3345; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3346; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3347; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3348; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3349; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3350; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3351; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3352; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3353; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3354; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3355; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3356; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3357; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3358; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3359; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3360; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3361; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3362; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3363; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3364; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3365; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3366; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3367; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3368; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3369; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3370; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3371; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3372; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3373; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3374; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3375; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3376; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3377; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3378; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3379; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3380; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3381; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3382; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3383; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3384; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3385; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3386; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3387; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3388; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3389; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3390; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3391; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3392; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3393; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3394; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3395; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3396; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3397; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3398; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3399; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3400; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3401; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3402; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3403; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3404; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3405; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3406; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3407; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3408; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3409; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3410; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3411; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3412; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3413; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3414; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3415; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3416; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3417; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3418; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3419; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3420; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3421; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3422; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3423; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3424; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3425; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3426; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3427; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3428; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3429; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3430; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3431; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3432; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3433; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3434; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3435; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3436; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3437; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3438; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3439; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3440; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3441; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3442; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3443; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3444; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3445; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3446; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3447; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3448; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3449; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3450; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3451; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3452; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3453; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3454; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3455; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3456; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3457; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3458; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3459; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3460; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3461; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3462; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3463; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3464; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3465; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3466; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3467; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3468; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3469; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3470; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3471; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3472; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3473; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3474; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3475; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3476; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3477; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3478; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3479; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3480; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3481; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3482; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3483; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3484; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3485; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3486; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3487; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3488; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3489; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3490; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3491; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3492; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3493; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3494; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3495; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3496; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3497; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3498; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3499; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3500; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3501; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3502; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3503; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3504; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3505; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3506; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3507; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3508; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3509; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3510; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3511; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3512; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3513; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3514; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3515; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3516; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3517; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3518; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3519; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3520; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3521; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3522; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3523; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3524; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3525; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3526; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3527; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3528; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3529; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3530; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3531; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3532; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3533; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3534; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3535; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3536; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3537; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3538; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3539; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3540; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3541; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3542; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3543; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3544; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3545; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3546; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3547; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3548; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3549; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3550; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3551; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3552; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3553; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3554; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3555; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3556; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3557; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3558; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3559; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3560; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3561; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3562; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3563; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3564; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3565; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3566; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3567; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3568; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3569; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3570; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3571; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3572; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3573; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3574; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3575; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3576; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3577; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3578; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3579; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3580; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3581; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3582; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3583; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3584; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3585; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3586; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3587; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3588; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3589; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3590; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3591; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3592; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3593; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3594; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3595; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3596; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3597; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3598; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3599; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3600; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3601; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3602; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3603; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3604; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3605; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3606; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3607; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3608; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3609; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3610; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3611; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3612; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3613; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3614; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3615; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3616; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3617; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3618; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3619; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3620; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3621; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3622; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3623; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3624; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3625; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3626; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3627; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3628; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3629; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3630; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3631; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3632; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3633; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3634; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3635; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3636; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3637; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3638; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3639; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3640; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3641; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3642; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3643; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3644; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3645; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3646; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3647; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3648; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3649; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3650; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3651; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3652; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3653; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3654; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3655; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3656; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3657; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3658; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3659; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3660; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3661; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3662; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3663; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3664; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3665; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3666; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3667; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3668; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3669; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3670; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3671; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3672; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3673; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3674; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3675; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3676; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3677; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3678; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3679; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3680; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3681; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3682; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3683; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3684; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3685; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3686; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3687; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3688; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3689; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3690; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3691; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3692; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3693; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3694; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3695; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3696; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3697; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3698; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3699; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3700; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3701; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3702; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3703; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3704; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3705; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3706; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3707; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3708; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3709; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3710; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3711; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3712; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3713; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3714; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3715; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3716; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3717; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3718; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3719; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3720; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3721; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3722; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3723; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3724; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3725; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3726; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3727; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3728; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3729; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3730; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3731; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3732; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3733; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3734; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3735; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3736; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3737; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3738; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3739; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3740; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3741; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3742; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3743; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3744; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3745; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3746; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3747; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3748; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3749; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3750; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3751; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3752; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3753; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3754; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3755; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3756; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3757; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3758; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3759; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3760; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3761; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3762; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3763; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3764; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3765; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3766; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3767; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3768; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3769; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3770; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3771; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3772; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3773; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3774; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3775; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3776; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3777; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3778; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3779; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3780; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3781; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3782; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3783; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3784; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3785; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3786; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3787; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3788; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3789; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3790; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3791; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3792; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3793; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3794; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3795; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3796; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3797; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3798; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3799; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3800; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3801; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3802; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3803; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3804; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3805; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3806; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3807; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3808; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3809; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3810; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3811; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3812; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3813; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3814; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3815; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3816; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3817; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3818; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3819; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3820; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3821; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3822; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3823; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3824; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3825; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3826; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3827; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3828; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3829; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3830; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3831; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3832; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3833; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3834; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3835; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3836; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3837; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3838; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3839; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3840; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3841; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3842; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3843; // @[RAM_ST.scala 32:46]
  wire [10:0] _GEN_3844; // @[RAM_ST.scala 32:46]
  wire [11:0] _T_3; // @[RAM_ST.scala 32:46]
  NestedCountersWithNumValid write_elem_counter ( // @[RAM_ST.scala 20:34]
    .CE(write_elem_counter_CE),
    .valid(write_elem_counter_valid)
  );
  NestedCountersWithNumValid read_elem_counter ( // @[RAM_ST.scala 21:33]
    .CE(read_elem_counter_CE),
    .valid(read_elem_counter_valid)
  );
  assign ram__T_8_addr = ram__T_8_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_8_data = ram[ram__T_8_addr]; // @[RAM_ST.scala 29:24]
  `else
  assign ram__T_8_data = ram__T_8_addr >= 11'h780 ? _RAND_1[7:0] : ram[ram__T_8_addr]; // @[RAM_ST.scala 29:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_2_data = WDATA;
  assign ram__T_2_addr = _T[10:0];
  assign ram__T_2_mask = 1'h1;
  assign ram__T_2_en = write_elem_counter_valid;
  assign _GEN_1 = 11'h1 == WADDR ? 11'h1 : 11'h0; // @[RAM_ST.scala 31:71]
  assign _GEN_2 = 11'h2 == WADDR ? 11'h2 : _GEN_1; // @[RAM_ST.scala 31:71]
  assign _GEN_3 = 11'h3 == WADDR ? 11'h3 : _GEN_2; // @[RAM_ST.scala 31:71]
  assign _GEN_4 = 11'h4 == WADDR ? 11'h4 : _GEN_3; // @[RAM_ST.scala 31:71]
  assign _GEN_5 = 11'h5 == WADDR ? 11'h5 : _GEN_4; // @[RAM_ST.scala 31:71]
  assign _GEN_6 = 11'h6 == WADDR ? 11'h6 : _GEN_5; // @[RAM_ST.scala 31:71]
  assign _GEN_7 = 11'h7 == WADDR ? 11'h7 : _GEN_6; // @[RAM_ST.scala 31:71]
  assign _GEN_8 = 11'h8 == WADDR ? 11'h8 : _GEN_7; // @[RAM_ST.scala 31:71]
  assign _GEN_9 = 11'h9 == WADDR ? 11'h9 : _GEN_8; // @[RAM_ST.scala 31:71]
  assign _GEN_10 = 11'ha == WADDR ? 11'ha : _GEN_9; // @[RAM_ST.scala 31:71]
  assign _GEN_11 = 11'hb == WADDR ? 11'hb : _GEN_10; // @[RAM_ST.scala 31:71]
  assign _GEN_12 = 11'hc == WADDR ? 11'hc : _GEN_11; // @[RAM_ST.scala 31:71]
  assign _GEN_13 = 11'hd == WADDR ? 11'hd : _GEN_12; // @[RAM_ST.scala 31:71]
  assign _GEN_14 = 11'he == WADDR ? 11'he : _GEN_13; // @[RAM_ST.scala 31:71]
  assign _GEN_15 = 11'hf == WADDR ? 11'hf : _GEN_14; // @[RAM_ST.scala 31:71]
  assign _GEN_16 = 11'h10 == WADDR ? 11'h10 : _GEN_15; // @[RAM_ST.scala 31:71]
  assign _GEN_17 = 11'h11 == WADDR ? 11'h11 : _GEN_16; // @[RAM_ST.scala 31:71]
  assign _GEN_18 = 11'h12 == WADDR ? 11'h12 : _GEN_17; // @[RAM_ST.scala 31:71]
  assign _GEN_19 = 11'h13 == WADDR ? 11'h13 : _GEN_18; // @[RAM_ST.scala 31:71]
  assign _GEN_20 = 11'h14 == WADDR ? 11'h14 : _GEN_19; // @[RAM_ST.scala 31:71]
  assign _GEN_21 = 11'h15 == WADDR ? 11'h15 : _GEN_20; // @[RAM_ST.scala 31:71]
  assign _GEN_22 = 11'h16 == WADDR ? 11'h16 : _GEN_21; // @[RAM_ST.scala 31:71]
  assign _GEN_23 = 11'h17 == WADDR ? 11'h17 : _GEN_22; // @[RAM_ST.scala 31:71]
  assign _GEN_24 = 11'h18 == WADDR ? 11'h18 : _GEN_23; // @[RAM_ST.scala 31:71]
  assign _GEN_25 = 11'h19 == WADDR ? 11'h19 : _GEN_24; // @[RAM_ST.scala 31:71]
  assign _GEN_26 = 11'h1a == WADDR ? 11'h1a : _GEN_25; // @[RAM_ST.scala 31:71]
  assign _GEN_27 = 11'h1b == WADDR ? 11'h1b : _GEN_26; // @[RAM_ST.scala 31:71]
  assign _GEN_28 = 11'h1c == WADDR ? 11'h1c : _GEN_27; // @[RAM_ST.scala 31:71]
  assign _GEN_29 = 11'h1d == WADDR ? 11'h1d : _GEN_28; // @[RAM_ST.scala 31:71]
  assign _GEN_30 = 11'h1e == WADDR ? 11'h1e : _GEN_29; // @[RAM_ST.scala 31:71]
  assign _GEN_31 = 11'h1f == WADDR ? 11'h1f : _GEN_30; // @[RAM_ST.scala 31:71]
  assign _GEN_32 = 11'h20 == WADDR ? 11'h20 : _GEN_31; // @[RAM_ST.scala 31:71]
  assign _GEN_33 = 11'h21 == WADDR ? 11'h21 : _GEN_32; // @[RAM_ST.scala 31:71]
  assign _GEN_34 = 11'h22 == WADDR ? 11'h22 : _GEN_33; // @[RAM_ST.scala 31:71]
  assign _GEN_35 = 11'h23 == WADDR ? 11'h23 : _GEN_34; // @[RAM_ST.scala 31:71]
  assign _GEN_36 = 11'h24 == WADDR ? 11'h24 : _GEN_35; // @[RAM_ST.scala 31:71]
  assign _GEN_37 = 11'h25 == WADDR ? 11'h25 : _GEN_36; // @[RAM_ST.scala 31:71]
  assign _GEN_38 = 11'h26 == WADDR ? 11'h26 : _GEN_37; // @[RAM_ST.scala 31:71]
  assign _GEN_39 = 11'h27 == WADDR ? 11'h27 : _GEN_38; // @[RAM_ST.scala 31:71]
  assign _GEN_40 = 11'h28 == WADDR ? 11'h28 : _GEN_39; // @[RAM_ST.scala 31:71]
  assign _GEN_41 = 11'h29 == WADDR ? 11'h29 : _GEN_40; // @[RAM_ST.scala 31:71]
  assign _GEN_42 = 11'h2a == WADDR ? 11'h2a : _GEN_41; // @[RAM_ST.scala 31:71]
  assign _GEN_43 = 11'h2b == WADDR ? 11'h2b : _GEN_42; // @[RAM_ST.scala 31:71]
  assign _GEN_44 = 11'h2c == WADDR ? 11'h2c : _GEN_43; // @[RAM_ST.scala 31:71]
  assign _GEN_45 = 11'h2d == WADDR ? 11'h2d : _GEN_44; // @[RAM_ST.scala 31:71]
  assign _GEN_46 = 11'h2e == WADDR ? 11'h2e : _GEN_45; // @[RAM_ST.scala 31:71]
  assign _GEN_47 = 11'h2f == WADDR ? 11'h2f : _GEN_46; // @[RAM_ST.scala 31:71]
  assign _GEN_48 = 11'h30 == WADDR ? 11'h30 : _GEN_47; // @[RAM_ST.scala 31:71]
  assign _GEN_49 = 11'h31 == WADDR ? 11'h31 : _GEN_48; // @[RAM_ST.scala 31:71]
  assign _GEN_50 = 11'h32 == WADDR ? 11'h32 : _GEN_49; // @[RAM_ST.scala 31:71]
  assign _GEN_51 = 11'h33 == WADDR ? 11'h33 : _GEN_50; // @[RAM_ST.scala 31:71]
  assign _GEN_52 = 11'h34 == WADDR ? 11'h34 : _GEN_51; // @[RAM_ST.scala 31:71]
  assign _GEN_53 = 11'h35 == WADDR ? 11'h35 : _GEN_52; // @[RAM_ST.scala 31:71]
  assign _GEN_54 = 11'h36 == WADDR ? 11'h36 : _GEN_53; // @[RAM_ST.scala 31:71]
  assign _GEN_55 = 11'h37 == WADDR ? 11'h37 : _GEN_54; // @[RAM_ST.scala 31:71]
  assign _GEN_56 = 11'h38 == WADDR ? 11'h38 : _GEN_55; // @[RAM_ST.scala 31:71]
  assign _GEN_57 = 11'h39 == WADDR ? 11'h39 : _GEN_56; // @[RAM_ST.scala 31:71]
  assign _GEN_58 = 11'h3a == WADDR ? 11'h3a : _GEN_57; // @[RAM_ST.scala 31:71]
  assign _GEN_59 = 11'h3b == WADDR ? 11'h3b : _GEN_58; // @[RAM_ST.scala 31:71]
  assign _GEN_60 = 11'h3c == WADDR ? 11'h3c : _GEN_59; // @[RAM_ST.scala 31:71]
  assign _GEN_61 = 11'h3d == WADDR ? 11'h3d : _GEN_60; // @[RAM_ST.scala 31:71]
  assign _GEN_62 = 11'h3e == WADDR ? 11'h3e : _GEN_61; // @[RAM_ST.scala 31:71]
  assign _GEN_63 = 11'h3f == WADDR ? 11'h3f : _GEN_62; // @[RAM_ST.scala 31:71]
  assign _GEN_64 = 11'h40 == WADDR ? 11'h40 : _GEN_63; // @[RAM_ST.scala 31:71]
  assign _GEN_65 = 11'h41 == WADDR ? 11'h41 : _GEN_64; // @[RAM_ST.scala 31:71]
  assign _GEN_66 = 11'h42 == WADDR ? 11'h42 : _GEN_65; // @[RAM_ST.scala 31:71]
  assign _GEN_67 = 11'h43 == WADDR ? 11'h43 : _GEN_66; // @[RAM_ST.scala 31:71]
  assign _GEN_68 = 11'h44 == WADDR ? 11'h44 : _GEN_67; // @[RAM_ST.scala 31:71]
  assign _GEN_69 = 11'h45 == WADDR ? 11'h45 : _GEN_68; // @[RAM_ST.scala 31:71]
  assign _GEN_70 = 11'h46 == WADDR ? 11'h46 : _GEN_69; // @[RAM_ST.scala 31:71]
  assign _GEN_71 = 11'h47 == WADDR ? 11'h47 : _GEN_70; // @[RAM_ST.scala 31:71]
  assign _GEN_72 = 11'h48 == WADDR ? 11'h48 : _GEN_71; // @[RAM_ST.scala 31:71]
  assign _GEN_73 = 11'h49 == WADDR ? 11'h49 : _GEN_72; // @[RAM_ST.scala 31:71]
  assign _GEN_74 = 11'h4a == WADDR ? 11'h4a : _GEN_73; // @[RAM_ST.scala 31:71]
  assign _GEN_75 = 11'h4b == WADDR ? 11'h4b : _GEN_74; // @[RAM_ST.scala 31:71]
  assign _GEN_76 = 11'h4c == WADDR ? 11'h4c : _GEN_75; // @[RAM_ST.scala 31:71]
  assign _GEN_77 = 11'h4d == WADDR ? 11'h4d : _GEN_76; // @[RAM_ST.scala 31:71]
  assign _GEN_78 = 11'h4e == WADDR ? 11'h4e : _GEN_77; // @[RAM_ST.scala 31:71]
  assign _GEN_79 = 11'h4f == WADDR ? 11'h4f : _GEN_78; // @[RAM_ST.scala 31:71]
  assign _GEN_80 = 11'h50 == WADDR ? 11'h50 : _GEN_79; // @[RAM_ST.scala 31:71]
  assign _GEN_81 = 11'h51 == WADDR ? 11'h51 : _GEN_80; // @[RAM_ST.scala 31:71]
  assign _GEN_82 = 11'h52 == WADDR ? 11'h52 : _GEN_81; // @[RAM_ST.scala 31:71]
  assign _GEN_83 = 11'h53 == WADDR ? 11'h53 : _GEN_82; // @[RAM_ST.scala 31:71]
  assign _GEN_84 = 11'h54 == WADDR ? 11'h54 : _GEN_83; // @[RAM_ST.scala 31:71]
  assign _GEN_85 = 11'h55 == WADDR ? 11'h55 : _GEN_84; // @[RAM_ST.scala 31:71]
  assign _GEN_86 = 11'h56 == WADDR ? 11'h56 : _GEN_85; // @[RAM_ST.scala 31:71]
  assign _GEN_87 = 11'h57 == WADDR ? 11'h57 : _GEN_86; // @[RAM_ST.scala 31:71]
  assign _GEN_88 = 11'h58 == WADDR ? 11'h58 : _GEN_87; // @[RAM_ST.scala 31:71]
  assign _GEN_89 = 11'h59 == WADDR ? 11'h59 : _GEN_88; // @[RAM_ST.scala 31:71]
  assign _GEN_90 = 11'h5a == WADDR ? 11'h5a : _GEN_89; // @[RAM_ST.scala 31:71]
  assign _GEN_91 = 11'h5b == WADDR ? 11'h5b : _GEN_90; // @[RAM_ST.scala 31:71]
  assign _GEN_92 = 11'h5c == WADDR ? 11'h5c : _GEN_91; // @[RAM_ST.scala 31:71]
  assign _GEN_93 = 11'h5d == WADDR ? 11'h5d : _GEN_92; // @[RAM_ST.scala 31:71]
  assign _GEN_94 = 11'h5e == WADDR ? 11'h5e : _GEN_93; // @[RAM_ST.scala 31:71]
  assign _GEN_95 = 11'h5f == WADDR ? 11'h5f : _GEN_94; // @[RAM_ST.scala 31:71]
  assign _GEN_96 = 11'h60 == WADDR ? 11'h60 : _GEN_95; // @[RAM_ST.scala 31:71]
  assign _GEN_97 = 11'h61 == WADDR ? 11'h61 : _GEN_96; // @[RAM_ST.scala 31:71]
  assign _GEN_98 = 11'h62 == WADDR ? 11'h62 : _GEN_97; // @[RAM_ST.scala 31:71]
  assign _GEN_99 = 11'h63 == WADDR ? 11'h63 : _GEN_98; // @[RAM_ST.scala 31:71]
  assign _GEN_100 = 11'h64 == WADDR ? 11'h64 : _GEN_99; // @[RAM_ST.scala 31:71]
  assign _GEN_101 = 11'h65 == WADDR ? 11'h65 : _GEN_100; // @[RAM_ST.scala 31:71]
  assign _GEN_102 = 11'h66 == WADDR ? 11'h66 : _GEN_101; // @[RAM_ST.scala 31:71]
  assign _GEN_103 = 11'h67 == WADDR ? 11'h67 : _GEN_102; // @[RAM_ST.scala 31:71]
  assign _GEN_104 = 11'h68 == WADDR ? 11'h68 : _GEN_103; // @[RAM_ST.scala 31:71]
  assign _GEN_105 = 11'h69 == WADDR ? 11'h69 : _GEN_104; // @[RAM_ST.scala 31:71]
  assign _GEN_106 = 11'h6a == WADDR ? 11'h6a : _GEN_105; // @[RAM_ST.scala 31:71]
  assign _GEN_107 = 11'h6b == WADDR ? 11'h6b : _GEN_106; // @[RAM_ST.scala 31:71]
  assign _GEN_108 = 11'h6c == WADDR ? 11'h6c : _GEN_107; // @[RAM_ST.scala 31:71]
  assign _GEN_109 = 11'h6d == WADDR ? 11'h6d : _GEN_108; // @[RAM_ST.scala 31:71]
  assign _GEN_110 = 11'h6e == WADDR ? 11'h6e : _GEN_109; // @[RAM_ST.scala 31:71]
  assign _GEN_111 = 11'h6f == WADDR ? 11'h6f : _GEN_110; // @[RAM_ST.scala 31:71]
  assign _GEN_112 = 11'h70 == WADDR ? 11'h70 : _GEN_111; // @[RAM_ST.scala 31:71]
  assign _GEN_113 = 11'h71 == WADDR ? 11'h71 : _GEN_112; // @[RAM_ST.scala 31:71]
  assign _GEN_114 = 11'h72 == WADDR ? 11'h72 : _GEN_113; // @[RAM_ST.scala 31:71]
  assign _GEN_115 = 11'h73 == WADDR ? 11'h73 : _GEN_114; // @[RAM_ST.scala 31:71]
  assign _GEN_116 = 11'h74 == WADDR ? 11'h74 : _GEN_115; // @[RAM_ST.scala 31:71]
  assign _GEN_117 = 11'h75 == WADDR ? 11'h75 : _GEN_116; // @[RAM_ST.scala 31:71]
  assign _GEN_118 = 11'h76 == WADDR ? 11'h76 : _GEN_117; // @[RAM_ST.scala 31:71]
  assign _GEN_119 = 11'h77 == WADDR ? 11'h77 : _GEN_118; // @[RAM_ST.scala 31:71]
  assign _GEN_120 = 11'h78 == WADDR ? 11'h78 : _GEN_119; // @[RAM_ST.scala 31:71]
  assign _GEN_121 = 11'h79 == WADDR ? 11'h79 : _GEN_120; // @[RAM_ST.scala 31:71]
  assign _GEN_122 = 11'h7a == WADDR ? 11'h7a : _GEN_121; // @[RAM_ST.scala 31:71]
  assign _GEN_123 = 11'h7b == WADDR ? 11'h7b : _GEN_122; // @[RAM_ST.scala 31:71]
  assign _GEN_124 = 11'h7c == WADDR ? 11'h7c : _GEN_123; // @[RAM_ST.scala 31:71]
  assign _GEN_125 = 11'h7d == WADDR ? 11'h7d : _GEN_124; // @[RAM_ST.scala 31:71]
  assign _GEN_126 = 11'h7e == WADDR ? 11'h7e : _GEN_125; // @[RAM_ST.scala 31:71]
  assign _GEN_127 = 11'h7f == WADDR ? 11'h7f : _GEN_126; // @[RAM_ST.scala 31:71]
  assign _GEN_128 = 11'h80 == WADDR ? 11'h80 : _GEN_127; // @[RAM_ST.scala 31:71]
  assign _GEN_129 = 11'h81 == WADDR ? 11'h81 : _GEN_128; // @[RAM_ST.scala 31:71]
  assign _GEN_130 = 11'h82 == WADDR ? 11'h82 : _GEN_129; // @[RAM_ST.scala 31:71]
  assign _GEN_131 = 11'h83 == WADDR ? 11'h83 : _GEN_130; // @[RAM_ST.scala 31:71]
  assign _GEN_132 = 11'h84 == WADDR ? 11'h84 : _GEN_131; // @[RAM_ST.scala 31:71]
  assign _GEN_133 = 11'h85 == WADDR ? 11'h85 : _GEN_132; // @[RAM_ST.scala 31:71]
  assign _GEN_134 = 11'h86 == WADDR ? 11'h86 : _GEN_133; // @[RAM_ST.scala 31:71]
  assign _GEN_135 = 11'h87 == WADDR ? 11'h87 : _GEN_134; // @[RAM_ST.scala 31:71]
  assign _GEN_136 = 11'h88 == WADDR ? 11'h88 : _GEN_135; // @[RAM_ST.scala 31:71]
  assign _GEN_137 = 11'h89 == WADDR ? 11'h89 : _GEN_136; // @[RAM_ST.scala 31:71]
  assign _GEN_138 = 11'h8a == WADDR ? 11'h8a : _GEN_137; // @[RAM_ST.scala 31:71]
  assign _GEN_139 = 11'h8b == WADDR ? 11'h8b : _GEN_138; // @[RAM_ST.scala 31:71]
  assign _GEN_140 = 11'h8c == WADDR ? 11'h8c : _GEN_139; // @[RAM_ST.scala 31:71]
  assign _GEN_141 = 11'h8d == WADDR ? 11'h8d : _GEN_140; // @[RAM_ST.scala 31:71]
  assign _GEN_142 = 11'h8e == WADDR ? 11'h8e : _GEN_141; // @[RAM_ST.scala 31:71]
  assign _GEN_143 = 11'h8f == WADDR ? 11'h8f : _GEN_142; // @[RAM_ST.scala 31:71]
  assign _GEN_144 = 11'h90 == WADDR ? 11'h90 : _GEN_143; // @[RAM_ST.scala 31:71]
  assign _GEN_145 = 11'h91 == WADDR ? 11'h91 : _GEN_144; // @[RAM_ST.scala 31:71]
  assign _GEN_146 = 11'h92 == WADDR ? 11'h92 : _GEN_145; // @[RAM_ST.scala 31:71]
  assign _GEN_147 = 11'h93 == WADDR ? 11'h93 : _GEN_146; // @[RAM_ST.scala 31:71]
  assign _GEN_148 = 11'h94 == WADDR ? 11'h94 : _GEN_147; // @[RAM_ST.scala 31:71]
  assign _GEN_149 = 11'h95 == WADDR ? 11'h95 : _GEN_148; // @[RAM_ST.scala 31:71]
  assign _GEN_150 = 11'h96 == WADDR ? 11'h96 : _GEN_149; // @[RAM_ST.scala 31:71]
  assign _GEN_151 = 11'h97 == WADDR ? 11'h97 : _GEN_150; // @[RAM_ST.scala 31:71]
  assign _GEN_152 = 11'h98 == WADDR ? 11'h98 : _GEN_151; // @[RAM_ST.scala 31:71]
  assign _GEN_153 = 11'h99 == WADDR ? 11'h99 : _GEN_152; // @[RAM_ST.scala 31:71]
  assign _GEN_154 = 11'h9a == WADDR ? 11'h9a : _GEN_153; // @[RAM_ST.scala 31:71]
  assign _GEN_155 = 11'h9b == WADDR ? 11'h9b : _GEN_154; // @[RAM_ST.scala 31:71]
  assign _GEN_156 = 11'h9c == WADDR ? 11'h9c : _GEN_155; // @[RAM_ST.scala 31:71]
  assign _GEN_157 = 11'h9d == WADDR ? 11'h9d : _GEN_156; // @[RAM_ST.scala 31:71]
  assign _GEN_158 = 11'h9e == WADDR ? 11'h9e : _GEN_157; // @[RAM_ST.scala 31:71]
  assign _GEN_159 = 11'h9f == WADDR ? 11'h9f : _GEN_158; // @[RAM_ST.scala 31:71]
  assign _GEN_160 = 11'ha0 == WADDR ? 11'ha0 : _GEN_159; // @[RAM_ST.scala 31:71]
  assign _GEN_161 = 11'ha1 == WADDR ? 11'ha1 : _GEN_160; // @[RAM_ST.scala 31:71]
  assign _GEN_162 = 11'ha2 == WADDR ? 11'ha2 : _GEN_161; // @[RAM_ST.scala 31:71]
  assign _GEN_163 = 11'ha3 == WADDR ? 11'ha3 : _GEN_162; // @[RAM_ST.scala 31:71]
  assign _GEN_164 = 11'ha4 == WADDR ? 11'ha4 : _GEN_163; // @[RAM_ST.scala 31:71]
  assign _GEN_165 = 11'ha5 == WADDR ? 11'ha5 : _GEN_164; // @[RAM_ST.scala 31:71]
  assign _GEN_166 = 11'ha6 == WADDR ? 11'ha6 : _GEN_165; // @[RAM_ST.scala 31:71]
  assign _GEN_167 = 11'ha7 == WADDR ? 11'ha7 : _GEN_166; // @[RAM_ST.scala 31:71]
  assign _GEN_168 = 11'ha8 == WADDR ? 11'ha8 : _GEN_167; // @[RAM_ST.scala 31:71]
  assign _GEN_169 = 11'ha9 == WADDR ? 11'ha9 : _GEN_168; // @[RAM_ST.scala 31:71]
  assign _GEN_170 = 11'haa == WADDR ? 11'haa : _GEN_169; // @[RAM_ST.scala 31:71]
  assign _GEN_171 = 11'hab == WADDR ? 11'hab : _GEN_170; // @[RAM_ST.scala 31:71]
  assign _GEN_172 = 11'hac == WADDR ? 11'hac : _GEN_171; // @[RAM_ST.scala 31:71]
  assign _GEN_173 = 11'had == WADDR ? 11'had : _GEN_172; // @[RAM_ST.scala 31:71]
  assign _GEN_174 = 11'hae == WADDR ? 11'hae : _GEN_173; // @[RAM_ST.scala 31:71]
  assign _GEN_175 = 11'haf == WADDR ? 11'haf : _GEN_174; // @[RAM_ST.scala 31:71]
  assign _GEN_176 = 11'hb0 == WADDR ? 11'hb0 : _GEN_175; // @[RAM_ST.scala 31:71]
  assign _GEN_177 = 11'hb1 == WADDR ? 11'hb1 : _GEN_176; // @[RAM_ST.scala 31:71]
  assign _GEN_178 = 11'hb2 == WADDR ? 11'hb2 : _GEN_177; // @[RAM_ST.scala 31:71]
  assign _GEN_179 = 11'hb3 == WADDR ? 11'hb3 : _GEN_178; // @[RAM_ST.scala 31:71]
  assign _GEN_180 = 11'hb4 == WADDR ? 11'hb4 : _GEN_179; // @[RAM_ST.scala 31:71]
  assign _GEN_181 = 11'hb5 == WADDR ? 11'hb5 : _GEN_180; // @[RAM_ST.scala 31:71]
  assign _GEN_182 = 11'hb6 == WADDR ? 11'hb6 : _GEN_181; // @[RAM_ST.scala 31:71]
  assign _GEN_183 = 11'hb7 == WADDR ? 11'hb7 : _GEN_182; // @[RAM_ST.scala 31:71]
  assign _GEN_184 = 11'hb8 == WADDR ? 11'hb8 : _GEN_183; // @[RAM_ST.scala 31:71]
  assign _GEN_185 = 11'hb9 == WADDR ? 11'hb9 : _GEN_184; // @[RAM_ST.scala 31:71]
  assign _GEN_186 = 11'hba == WADDR ? 11'hba : _GEN_185; // @[RAM_ST.scala 31:71]
  assign _GEN_187 = 11'hbb == WADDR ? 11'hbb : _GEN_186; // @[RAM_ST.scala 31:71]
  assign _GEN_188 = 11'hbc == WADDR ? 11'hbc : _GEN_187; // @[RAM_ST.scala 31:71]
  assign _GEN_189 = 11'hbd == WADDR ? 11'hbd : _GEN_188; // @[RAM_ST.scala 31:71]
  assign _GEN_190 = 11'hbe == WADDR ? 11'hbe : _GEN_189; // @[RAM_ST.scala 31:71]
  assign _GEN_191 = 11'hbf == WADDR ? 11'hbf : _GEN_190; // @[RAM_ST.scala 31:71]
  assign _GEN_192 = 11'hc0 == WADDR ? 11'hc0 : _GEN_191; // @[RAM_ST.scala 31:71]
  assign _GEN_193 = 11'hc1 == WADDR ? 11'hc1 : _GEN_192; // @[RAM_ST.scala 31:71]
  assign _GEN_194 = 11'hc2 == WADDR ? 11'hc2 : _GEN_193; // @[RAM_ST.scala 31:71]
  assign _GEN_195 = 11'hc3 == WADDR ? 11'hc3 : _GEN_194; // @[RAM_ST.scala 31:71]
  assign _GEN_196 = 11'hc4 == WADDR ? 11'hc4 : _GEN_195; // @[RAM_ST.scala 31:71]
  assign _GEN_197 = 11'hc5 == WADDR ? 11'hc5 : _GEN_196; // @[RAM_ST.scala 31:71]
  assign _GEN_198 = 11'hc6 == WADDR ? 11'hc6 : _GEN_197; // @[RAM_ST.scala 31:71]
  assign _GEN_199 = 11'hc7 == WADDR ? 11'hc7 : _GEN_198; // @[RAM_ST.scala 31:71]
  assign _GEN_200 = 11'hc8 == WADDR ? 11'hc8 : _GEN_199; // @[RAM_ST.scala 31:71]
  assign _GEN_201 = 11'hc9 == WADDR ? 11'hc9 : _GEN_200; // @[RAM_ST.scala 31:71]
  assign _GEN_202 = 11'hca == WADDR ? 11'hca : _GEN_201; // @[RAM_ST.scala 31:71]
  assign _GEN_203 = 11'hcb == WADDR ? 11'hcb : _GEN_202; // @[RAM_ST.scala 31:71]
  assign _GEN_204 = 11'hcc == WADDR ? 11'hcc : _GEN_203; // @[RAM_ST.scala 31:71]
  assign _GEN_205 = 11'hcd == WADDR ? 11'hcd : _GEN_204; // @[RAM_ST.scala 31:71]
  assign _GEN_206 = 11'hce == WADDR ? 11'hce : _GEN_205; // @[RAM_ST.scala 31:71]
  assign _GEN_207 = 11'hcf == WADDR ? 11'hcf : _GEN_206; // @[RAM_ST.scala 31:71]
  assign _GEN_208 = 11'hd0 == WADDR ? 11'hd0 : _GEN_207; // @[RAM_ST.scala 31:71]
  assign _GEN_209 = 11'hd1 == WADDR ? 11'hd1 : _GEN_208; // @[RAM_ST.scala 31:71]
  assign _GEN_210 = 11'hd2 == WADDR ? 11'hd2 : _GEN_209; // @[RAM_ST.scala 31:71]
  assign _GEN_211 = 11'hd3 == WADDR ? 11'hd3 : _GEN_210; // @[RAM_ST.scala 31:71]
  assign _GEN_212 = 11'hd4 == WADDR ? 11'hd4 : _GEN_211; // @[RAM_ST.scala 31:71]
  assign _GEN_213 = 11'hd5 == WADDR ? 11'hd5 : _GEN_212; // @[RAM_ST.scala 31:71]
  assign _GEN_214 = 11'hd6 == WADDR ? 11'hd6 : _GEN_213; // @[RAM_ST.scala 31:71]
  assign _GEN_215 = 11'hd7 == WADDR ? 11'hd7 : _GEN_214; // @[RAM_ST.scala 31:71]
  assign _GEN_216 = 11'hd8 == WADDR ? 11'hd8 : _GEN_215; // @[RAM_ST.scala 31:71]
  assign _GEN_217 = 11'hd9 == WADDR ? 11'hd9 : _GEN_216; // @[RAM_ST.scala 31:71]
  assign _GEN_218 = 11'hda == WADDR ? 11'hda : _GEN_217; // @[RAM_ST.scala 31:71]
  assign _GEN_219 = 11'hdb == WADDR ? 11'hdb : _GEN_218; // @[RAM_ST.scala 31:71]
  assign _GEN_220 = 11'hdc == WADDR ? 11'hdc : _GEN_219; // @[RAM_ST.scala 31:71]
  assign _GEN_221 = 11'hdd == WADDR ? 11'hdd : _GEN_220; // @[RAM_ST.scala 31:71]
  assign _GEN_222 = 11'hde == WADDR ? 11'hde : _GEN_221; // @[RAM_ST.scala 31:71]
  assign _GEN_223 = 11'hdf == WADDR ? 11'hdf : _GEN_222; // @[RAM_ST.scala 31:71]
  assign _GEN_224 = 11'he0 == WADDR ? 11'he0 : _GEN_223; // @[RAM_ST.scala 31:71]
  assign _GEN_225 = 11'he1 == WADDR ? 11'he1 : _GEN_224; // @[RAM_ST.scala 31:71]
  assign _GEN_226 = 11'he2 == WADDR ? 11'he2 : _GEN_225; // @[RAM_ST.scala 31:71]
  assign _GEN_227 = 11'he3 == WADDR ? 11'he3 : _GEN_226; // @[RAM_ST.scala 31:71]
  assign _GEN_228 = 11'he4 == WADDR ? 11'he4 : _GEN_227; // @[RAM_ST.scala 31:71]
  assign _GEN_229 = 11'he5 == WADDR ? 11'he5 : _GEN_228; // @[RAM_ST.scala 31:71]
  assign _GEN_230 = 11'he6 == WADDR ? 11'he6 : _GEN_229; // @[RAM_ST.scala 31:71]
  assign _GEN_231 = 11'he7 == WADDR ? 11'he7 : _GEN_230; // @[RAM_ST.scala 31:71]
  assign _GEN_232 = 11'he8 == WADDR ? 11'he8 : _GEN_231; // @[RAM_ST.scala 31:71]
  assign _GEN_233 = 11'he9 == WADDR ? 11'he9 : _GEN_232; // @[RAM_ST.scala 31:71]
  assign _GEN_234 = 11'hea == WADDR ? 11'hea : _GEN_233; // @[RAM_ST.scala 31:71]
  assign _GEN_235 = 11'heb == WADDR ? 11'heb : _GEN_234; // @[RAM_ST.scala 31:71]
  assign _GEN_236 = 11'hec == WADDR ? 11'hec : _GEN_235; // @[RAM_ST.scala 31:71]
  assign _GEN_237 = 11'hed == WADDR ? 11'hed : _GEN_236; // @[RAM_ST.scala 31:71]
  assign _GEN_238 = 11'hee == WADDR ? 11'hee : _GEN_237; // @[RAM_ST.scala 31:71]
  assign _GEN_239 = 11'hef == WADDR ? 11'hef : _GEN_238; // @[RAM_ST.scala 31:71]
  assign _GEN_240 = 11'hf0 == WADDR ? 11'hf0 : _GEN_239; // @[RAM_ST.scala 31:71]
  assign _GEN_241 = 11'hf1 == WADDR ? 11'hf1 : _GEN_240; // @[RAM_ST.scala 31:71]
  assign _GEN_242 = 11'hf2 == WADDR ? 11'hf2 : _GEN_241; // @[RAM_ST.scala 31:71]
  assign _GEN_243 = 11'hf3 == WADDR ? 11'hf3 : _GEN_242; // @[RAM_ST.scala 31:71]
  assign _GEN_244 = 11'hf4 == WADDR ? 11'hf4 : _GEN_243; // @[RAM_ST.scala 31:71]
  assign _GEN_245 = 11'hf5 == WADDR ? 11'hf5 : _GEN_244; // @[RAM_ST.scala 31:71]
  assign _GEN_246 = 11'hf6 == WADDR ? 11'hf6 : _GEN_245; // @[RAM_ST.scala 31:71]
  assign _GEN_247 = 11'hf7 == WADDR ? 11'hf7 : _GEN_246; // @[RAM_ST.scala 31:71]
  assign _GEN_248 = 11'hf8 == WADDR ? 11'hf8 : _GEN_247; // @[RAM_ST.scala 31:71]
  assign _GEN_249 = 11'hf9 == WADDR ? 11'hf9 : _GEN_248; // @[RAM_ST.scala 31:71]
  assign _GEN_250 = 11'hfa == WADDR ? 11'hfa : _GEN_249; // @[RAM_ST.scala 31:71]
  assign _GEN_251 = 11'hfb == WADDR ? 11'hfb : _GEN_250; // @[RAM_ST.scala 31:71]
  assign _GEN_252 = 11'hfc == WADDR ? 11'hfc : _GEN_251; // @[RAM_ST.scala 31:71]
  assign _GEN_253 = 11'hfd == WADDR ? 11'hfd : _GEN_252; // @[RAM_ST.scala 31:71]
  assign _GEN_254 = 11'hfe == WADDR ? 11'hfe : _GEN_253; // @[RAM_ST.scala 31:71]
  assign _GEN_255 = 11'hff == WADDR ? 11'hff : _GEN_254; // @[RAM_ST.scala 31:71]
  assign _GEN_256 = 11'h100 == WADDR ? 11'h100 : _GEN_255; // @[RAM_ST.scala 31:71]
  assign _GEN_257 = 11'h101 == WADDR ? 11'h101 : _GEN_256; // @[RAM_ST.scala 31:71]
  assign _GEN_258 = 11'h102 == WADDR ? 11'h102 : _GEN_257; // @[RAM_ST.scala 31:71]
  assign _GEN_259 = 11'h103 == WADDR ? 11'h103 : _GEN_258; // @[RAM_ST.scala 31:71]
  assign _GEN_260 = 11'h104 == WADDR ? 11'h104 : _GEN_259; // @[RAM_ST.scala 31:71]
  assign _GEN_261 = 11'h105 == WADDR ? 11'h105 : _GEN_260; // @[RAM_ST.scala 31:71]
  assign _GEN_262 = 11'h106 == WADDR ? 11'h106 : _GEN_261; // @[RAM_ST.scala 31:71]
  assign _GEN_263 = 11'h107 == WADDR ? 11'h107 : _GEN_262; // @[RAM_ST.scala 31:71]
  assign _GEN_264 = 11'h108 == WADDR ? 11'h108 : _GEN_263; // @[RAM_ST.scala 31:71]
  assign _GEN_265 = 11'h109 == WADDR ? 11'h109 : _GEN_264; // @[RAM_ST.scala 31:71]
  assign _GEN_266 = 11'h10a == WADDR ? 11'h10a : _GEN_265; // @[RAM_ST.scala 31:71]
  assign _GEN_267 = 11'h10b == WADDR ? 11'h10b : _GEN_266; // @[RAM_ST.scala 31:71]
  assign _GEN_268 = 11'h10c == WADDR ? 11'h10c : _GEN_267; // @[RAM_ST.scala 31:71]
  assign _GEN_269 = 11'h10d == WADDR ? 11'h10d : _GEN_268; // @[RAM_ST.scala 31:71]
  assign _GEN_270 = 11'h10e == WADDR ? 11'h10e : _GEN_269; // @[RAM_ST.scala 31:71]
  assign _GEN_271 = 11'h10f == WADDR ? 11'h10f : _GEN_270; // @[RAM_ST.scala 31:71]
  assign _GEN_272 = 11'h110 == WADDR ? 11'h110 : _GEN_271; // @[RAM_ST.scala 31:71]
  assign _GEN_273 = 11'h111 == WADDR ? 11'h111 : _GEN_272; // @[RAM_ST.scala 31:71]
  assign _GEN_274 = 11'h112 == WADDR ? 11'h112 : _GEN_273; // @[RAM_ST.scala 31:71]
  assign _GEN_275 = 11'h113 == WADDR ? 11'h113 : _GEN_274; // @[RAM_ST.scala 31:71]
  assign _GEN_276 = 11'h114 == WADDR ? 11'h114 : _GEN_275; // @[RAM_ST.scala 31:71]
  assign _GEN_277 = 11'h115 == WADDR ? 11'h115 : _GEN_276; // @[RAM_ST.scala 31:71]
  assign _GEN_278 = 11'h116 == WADDR ? 11'h116 : _GEN_277; // @[RAM_ST.scala 31:71]
  assign _GEN_279 = 11'h117 == WADDR ? 11'h117 : _GEN_278; // @[RAM_ST.scala 31:71]
  assign _GEN_280 = 11'h118 == WADDR ? 11'h118 : _GEN_279; // @[RAM_ST.scala 31:71]
  assign _GEN_281 = 11'h119 == WADDR ? 11'h119 : _GEN_280; // @[RAM_ST.scala 31:71]
  assign _GEN_282 = 11'h11a == WADDR ? 11'h11a : _GEN_281; // @[RAM_ST.scala 31:71]
  assign _GEN_283 = 11'h11b == WADDR ? 11'h11b : _GEN_282; // @[RAM_ST.scala 31:71]
  assign _GEN_284 = 11'h11c == WADDR ? 11'h11c : _GEN_283; // @[RAM_ST.scala 31:71]
  assign _GEN_285 = 11'h11d == WADDR ? 11'h11d : _GEN_284; // @[RAM_ST.scala 31:71]
  assign _GEN_286 = 11'h11e == WADDR ? 11'h11e : _GEN_285; // @[RAM_ST.scala 31:71]
  assign _GEN_287 = 11'h11f == WADDR ? 11'h11f : _GEN_286; // @[RAM_ST.scala 31:71]
  assign _GEN_288 = 11'h120 == WADDR ? 11'h120 : _GEN_287; // @[RAM_ST.scala 31:71]
  assign _GEN_289 = 11'h121 == WADDR ? 11'h121 : _GEN_288; // @[RAM_ST.scala 31:71]
  assign _GEN_290 = 11'h122 == WADDR ? 11'h122 : _GEN_289; // @[RAM_ST.scala 31:71]
  assign _GEN_291 = 11'h123 == WADDR ? 11'h123 : _GEN_290; // @[RAM_ST.scala 31:71]
  assign _GEN_292 = 11'h124 == WADDR ? 11'h124 : _GEN_291; // @[RAM_ST.scala 31:71]
  assign _GEN_293 = 11'h125 == WADDR ? 11'h125 : _GEN_292; // @[RAM_ST.scala 31:71]
  assign _GEN_294 = 11'h126 == WADDR ? 11'h126 : _GEN_293; // @[RAM_ST.scala 31:71]
  assign _GEN_295 = 11'h127 == WADDR ? 11'h127 : _GEN_294; // @[RAM_ST.scala 31:71]
  assign _GEN_296 = 11'h128 == WADDR ? 11'h128 : _GEN_295; // @[RAM_ST.scala 31:71]
  assign _GEN_297 = 11'h129 == WADDR ? 11'h129 : _GEN_296; // @[RAM_ST.scala 31:71]
  assign _GEN_298 = 11'h12a == WADDR ? 11'h12a : _GEN_297; // @[RAM_ST.scala 31:71]
  assign _GEN_299 = 11'h12b == WADDR ? 11'h12b : _GEN_298; // @[RAM_ST.scala 31:71]
  assign _GEN_300 = 11'h12c == WADDR ? 11'h12c : _GEN_299; // @[RAM_ST.scala 31:71]
  assign _GEN_301 = 11'h12d == WADDR ? 11'h12d : _GEN_300; // @[RAM_ST.scala 31:71]
  assign _GEN_302 = 11'h12e == WADDR ? 11'h12e : _GEN_301; // @[RAM_ST.scala 31:71]
  assign _GEN_303 = 11'h12f == WADDR ? 11'h12f : _GEN_302; // @[RAM_ST.scala 31:71]
  assign _GEN_304 = 11'h130 == WADDR ? 11'h130 : _GEN_303; // @[RAM_ST.scala 31:71]
  assign _GEN_305 = 11'h131 == WADDR ? 11'h131 : _GEN_304; // @[RAM_ST.scala 31:71]
  assign _GEN_306 = 11'h132 == WADDR ? 11'h132 : _GEN_305; // @[RAM_ST.scala 31:71]
  assign _GEN_307 = 11'h133 == WADDR ? 11'h133 : _GEN_306; // @[RAM_ST.scala 31:71]
  assign _GEN_308 = 11'h134 == WADDR ? 11'h134 : _GEN_307; // @[RAM_ST.scala 31:71]
  assign _GEN_309 = 11'h135 == WADDR ? 11'h135 : _GEN_308; // @[RAM_ST.scala 31:71]
  assign _GEN_310 = 11'h136 == WADDR ? 11'h136 : _GEN_309; // @[RAM_ST.scala 31:71]
  assign _GEN_311 = 11'h137 == WADDR ? 11'h137 : _GEN_310; // @[RAM_ST.scala 31:71]
  assign _GEN_312 = 11'h138 == WADDR ? 11'h138 : _GEN_311; // @[RAM_ST.scala 31:71]
  assign _GEN_313 = 11'h139 == WADDR ? 11'h139 : _GEN_312; // @[RAM_ST.scala 31:71]
  assign _GEN_314 = 11'h13a == WADDR ? 11'h13a : _GEN_313; // @[RAM_ST.scala 31:71]
  assign _GEN_315 = 11'h13b == WADDR ? 11'h13b : _GEN_314; // @[RAM_ST.scala 31:71]
  assign _GEN_316 = 11'h13c == WADDR ? 11'h13c : _GEN_315; // @[RAM_ST.scala 31:71]
  assign _GEN_317 = 11'h13d == WADDR ? 11'h13d : _GEN_316; // @[RAM_ST.scala 31:71]
  assign _GEN_318 = 11'h13e == WADDR ? 11'h13e : _GEN_317; // @[RAM_ST.scala 31:71]
  assign _GEN_319 = 11'h13f == WADDR ? 11'h13f : _GEN_318; // @[RAM_ST.scala 31:71]
  assign _GEN_320 = 11'h140 == WADDR ? 11'h140 : _GEN_319; // @[RAM_ST.scala 31:71]
  assign _GEN_321 = 11'h141 == WADDR ? 11'h141 : _GEN_320; // @[RAM_ST.scala 31:71]
  assign _GEN_322 = 11'h142 == WADDR ? 11'h142 : _GEN_321; // @[RAM_ST.scala 31:71]
  assign _GEN_323 = 11'h143 == WADDR ? 11'h143 : _GEN_322; // @[RAM_ST.scala 31:71]
  assign _GEN_324 = 11'h144 == WADDR ? 11'h144 : _GEN_323; // @[RAM_ST.scala 31:71]
  assign _GEN_325 = 11'h145 == WADDR ? 11'h145 : _GEN_324; // @[RAM_ST.scala 31:71]
  assign _GEN_326 = 11'h146 == WADDR ? 11'h146 : _GEN_325; // @[RAM_ST.scala 31:71]
  assign _GEN_327 = 11'h147 == WADDR ? 11'h147 : _GEN_326; // @[RAM_ST.scala 31:71]
  assign _GEN_328 = 11'h148 == WADDR ? 11'h148 : _GEN_327; // @[RAM_ST.scala 31:71]
  assign _GEN_329 = 11'h149 == WADDR ? 11'h149 : _GEN_328; // @[RAM_ST.scala 31:71]
  assign _GEN_330 = 11'h14a == WADDR ? 11'h14a : _GEN_329; // @[RAM_ST.scala 31:71]
  assign _GEN_331 = 11'h14b == WADDR ? 11'h14b : _GEN_330; // @[RAM_ST.scala 31:71]
  assign _GEN_332 = 11'h14c == WADDR ? 11'h14c : _GEN_331; // @[RAM_ST.scala 31:71]
  assign _GEN_333 = 11'h14d == WADDR ? 11'h14d : _GEN_332; // @[RAM_ST.scala 31:71]
  assign _GEN_334 = 11'h14e == WADDR ? 11'h14e : _GEN_333; // @[RAM_ST.scala 31:71]
  assign _GEN_335 = 11'h14f == WADDR ? 11'h14f : _GEN_334; // @[RAM_ST.scala 31:71]
  assign _GEN_336 = 11'h150 == WADDR ? 11'h150 : _GEN_335; // @[RAM_ST.scala 31:71]
  assign _GEN_337 = 11'h151 == WADDR ? 11'h151 : _GEN_336; // @[RAM_ST.scala 31:71]
  assign _GEN_338 = 11'h152 == WADDR ? 11'h152 : _GEN_337; // @[RAM_ST.scala 31:71]
  assign _GEN_339 = 11'h153 == WADDR ? 11'h153 : _GEN_338; // @[RAM_ST.scala 31:71]
  assign _GEN_340 = 11'h154 == WADDR ? 11'h154 : _GEN_339; // @[RAM_ST.scala 31:71]
  assign _GEN_341 = 11'h155 == WADDR ? 11'h155 : _GEN_340; // @[RAM_ST.scala 31:71]
  assign _GEN_342 = 11'h156 == WADDR ? 11'h156 : _GEN_341; // @[RAM_ST.scala 31:71]
  assign _GEN_343 = 11'h157 == WADDR ? 11'h157 : _GEN_342; // @[RAM_ST.scala 31:71]
  assign _GEN_344 = 11'h158 == WADDR ? 11'h158 : _GEN_343; // @[RAM_ST.scala 31:71]
  assign _GEN_345 = 11'h159 == WADDR ? 11'h159 : _GEN_344; // @[RAM_ST.scala 31:71]
  assign _GEN_346 = 11'h15a == WADDR ? 11'h15a : _GEN_345; // @[RAM_ST.scala 31:71]
  assign _GEN_347 = 11'h15b == WADDR ? 11'h15b : _GEN_346; // @[RAM_ST.scala 31:71]
  assign _GEN_348 = 11'h15c == WADDR ? 11'h15c : _GEN_347; // @[RAM_ST.scala 31:71]
  assign _GEN_349 = 11'h15d == WADDR ? 11'h15d : _GEN_348; // @[RAM_ST.scala 31:71]
  assign _GEN_350 = 11'h15e == WADDR ? 11'h15e : _GEN_349; // @[RAM_ST.scala 31:71]
  assign _GEN_351 = 11'h15f == WADDR ? 11'h15f : _GEN_350; // @[RAM_ST.scala 31:71]
  assign _GEN_352 = 11'h160 == WADDR ? 11'h160 : _GEN_351; // @[RAM_ST.scala 31:71]
  assign _GEN_353 = 11'h161 == WADDR ? 11'h161 : _GEN_352; // @[RAM_ST.scala 31:71]
  assign _GEN_354 = 11'h162 == WADDR ? 11'h162 : _GEN_353; // @[RAM_ST.scala 31:71]
  assign _GEN_355 = 11'h163 == WADDR ? 11'h163 : _GEN_354; // @[RAM_ST.scala 31:71]
  assign _GEN_356 = 11'h164 == WADDR ? 11'h164 : _GEN_355; // @[RAM_ST.scala 31:71]
  assign _GEN_357 = 11'h165 == WADDR ? 11'h165 : _GEN_356; // @[RAM_ST.scala 31:71]
  assign _GEN_358 = 11'h166 == WADDR ? 11'h166 : _GEN_357; // @[RAM_ST.scala 31:71]
  assign _GEN_359 = 11'h167 == WADDR ? 11'h167 : _GEN_358; // @[RAM_ST.scala 31:71]
  assign _GEN_360 = 11'h168 == WADDR ? 11'h168 : _GEN_359; // @[RAM_ST.scala 31:71]
  assign _GEN_361 = 11'h169 == WADDR ? 11'h169 : _GEN_360; // @[RAM_ST.scala 31:71]
  assign _GEN_362 = 11'h16a == WADDR ? 11'h16a : _GEN_361; // @[RAM_ST.scala 31:71]
  assign _GEN_363 = 11'h16b == WADDR ? 11'h16b : _GEN_362; // @[RAM_ST.scala 31:71]
  assign _GEN_364 = 11'h16c == WADDR ? 11'h16c : _GEN_363; // @[RAM_ST.scala 31:71]
  assign _GEN_365 = 11'h16d == WADDR ? 11'h16d : _GEN_364; // @[RAM_ST.scala 31:71]
  assign _GEN_366 = 11'h16e == WADDR ? 11'h16e : _GEN_365; // @[RAM_ST.scala 31:71]
  assign _GEN_367 = 11'h16f == WADDR ? 11'h16f : _GEN_366; // @[RAM_ST.scala 31:71]
  assign _GEN_368 = 11'h170 == WADDR ? 11'h170 : _GEN_367; // @[RAM_ST.scala 31:71]
  assign _GEN_369 = 11'h171 == WADDR ? 11'h171 : _GEN_368; // @[RAM_ST.scala 31:71]
  assign _GEN_370 = 11'h172 == WADDR ? 11'h172 : _GEN_369; // @[RAM_ST.scala 31:71]
  assign _GEN_371 = 11'h173 == WADDR ? 11'h173 : _GEN_370; // @[RAM_ST.scala 31:71]
  assign _GEN_372 = 11'h174 == WADDR ? 11'h174 : _GEN_371; // @[RAM_ST.scala 31:71]
  assign _GEN_373 = 11'h175 == WADDR ? 11'h175 : _GEN_372; // @[RAM_ST.scala 31:71]
  assign _GEN_374 = 11'h176 == WADDR ? 11'h176 : _GEN_373; // @[RAM_ST.scala 31:71]
  assign _GEN_375 = 11'h177 == WADDR ? 11'h177 : _GEN_374; // @[RAM_ST.scala 31:71]
  assign _GEN_376 = 11'h178 == WADDR ? 11'h178 : _GEN_375; // @[RAM_ST.scala 31:71]
  assign _GEN_377 = 11'h179 == WADDR ? 11'h179 : _GEN_376; // @[RAM_ST.scala 31:71]
  assign _GEN_378 = 11'h17a == WADDR ? 11'h17a : _GEN_377; // @[RAM_ST.scala 31:71]
  assign _GEN_379 = 11'h17b == WADDR ? 11'h17b : _GEN_378; // @[RAM_ST.scala 31:71]
  assign _GEN_380 = 11'h17c == WADDR ? 11'h17c : _GEN_379; // @[RAM_ST.scala 31:71]
  assign _GEN_381 = 11'h17d == WADDR ? 11'h17d : _GEN_380; // @[RAM_ST.scala 31:71]
  assign _GEN_382 = 11'h17e == WADDR ? 11'h17e : _GEN_381; // @[RAM_ST.scala 31:71]
  assign _GEN_383 = 11'h17f == WADDR ? 11'h17f : _GEN_382; // @[RAM_ST.scala 31:71]
  assign _GEN_384 = 11'h180 == WADDR ? 11'h180 : _GEN_383; // @[RAM_ST.scala 31:71]
  assign _GEN_385 = 11'h181 == WADDR ? 11'h181 : _GEN_384; // @[RAM_ST.scala 31:71]
  assign _GEN_386 = 11'h182 == WADDR ? 11'h182 : _GEN_385; // @[RAM_ST.scala 31:71]
  assign _GEN_387 = 11'h183 == WADDR ? 11'h183 : _GEN_386; // @[RAM_ST.scala 31:71]
  assign _GEN_388 = 11'h184 == WADDR ? 11'h184 : _GEN_387; // @[RAM_ST.scala 31:71]
  assign _GEN_389 = 11'h185 == WADDR ? 11'h185 : _GEN_388; // @[RAM_ST.scala 31:71]
  assign _GEN_390 = 11'h186 == WADDR ? 11'h186 : _GEN_389; // @[RAM_ST.scala 31:71]
  assign _GEN_391 = 11'h187 == WADDR ? 11'h187 : _GEN_390; // @[RAM_ST.scala 31:71]
  assign _GEN_392 = 11'h188 == WADDR ? 11'h188 : _GEN_391; // @[RAM_ST.scala 31:71]
  assign _GEN_393 = 11'h189 == WADDR ? 11'h189 : _GEN_392; // @[RAM_ST.scala 31:71]
  assign _GEN_394 = 11'h18a == WADDR ? 11'h18a : _GEN_393; // @[RAM_ST.scala 31:71]
  assign _GEN_395 = 11'h18b == WADDR ? 11'h18b : _GEN_394; // @[RAM_ST.scala 31:71]
  assign _GEN_396 = 11'h18c == WADDR ? 11'h18c : _GEN_395; // @[RAM_ST.scala 31:71]
  assign _GEN_397 = 11'h18d == WADDR ? 11'h18d : _GEN_396; // @[RAM_ST.scala 31:71]
  assign _GEN_398 = 11'h18e == WADDR ? 11'h18e : _GEN_397; // @[RAM_ST.scala 31:71]
  assign _GEN_399 = 11'h18f == WADDR ? 11'h18f : _GEN_398; // @[RAM_ST.scala 31:71]
  assign _GEN_400 = 11'h190 == WADDR ? 11'h190 : _GEN_399; // @[RAM_ST.scala 31:71]
  assign _GEN_401 = 11'h191 == WADDR ? 11'h191 : _GEN_400; // @[RAM_ST.scala 31:71]
  assign _GEN_402 = 11'h192 == WADDR ? 11'h192 : _GEN_401; // @[RAM_ST.scala 31:71]
  assign _GEN_403 = 11'h193 == WADDR ? 11'h193 : _GEN_402; // @[RAM_ST.scala 31:71]
  assign _GEN_404 = 11'h194 == WADDR ? 11'h194 : _GEN_403; // @[RAM_ST.scala 31:71]
  assign _GEN_405 = 11'h195 == WADDR ? 11'h195 : _GEN_404; // @[RAM_ST.scala 31:71]
  assign _GEN_406 = 11'h196 == WADDR ? 11'h196 : _GEN_405; // @[RAM_ST.scala 31:71]
  assign _GEN_407 = 11'h197 == WADDR ? 11'h197 : _GEN_406; // @[RAM_ST.scala 31:71]
  assign _GEN_408 = 11'h198 == WADDR ? 11'h198 : _GEN_407; // @[RAM_ST.scala 31:71]
  assign _GEN_409 = 11'h199 == WADDR ? 11'h199 : _GEN_408; // @[RAM_ST.scala 31:71]
  assign _GEN_410 = 11'h19a == WADDR ? 11'h19a : _GEN_409; // @[RAM_ST.scala 31:71]
  assign _GEN_411 = 11'h19b == WADDR ? 11'h19b : _GEN_410; // @[RAM_ST.scala 31:71]
  assign _GEN_412 = 11'h19c == WADDR ? 11'h19c : _GEN_411; // @[RAM_ST.scala 31:71]
  assign _GEN_413 = 11'h19d == WADDR ? 11'h19d : _GEN_412; // @[RAM_ST.scala 31:71]
  assign _GEN_414 = 11'h19e == WADDR ? 11'h19e : _GEN_413; // @[RAM_ST.scala 31:71]
  assign _GEN_415 = 11'h19f == WADDR ? 11'h19f : _GEN_414; // @[RAM_ST.scala 31:71]
  assign _GEN_416 = 11'h1a0 == WADDR ? 11'h1a0 : _GEN_415; // @[RAM_ST.scala 31:71]
  assign _GEN_417 = 11'h1a1 == WADDR ? 11'h1a1 : _GEN_416; // @[RAM_ST.scala 31:71]
  assign _GEN_418 = 11'h1a2 == WADDR ? 11'h1a2 : _GEN_417; // @[RAM_ST.scala 31:71]
  assign _GEN_419 = 11'h1a3 == WADDR ? 11'h1a3 : _GEN_418; // @[RAM_ST.scala 31:71]
  assign _GEN_420 = 11'h1a4 == WADDR ? 11'h1a4 : _GEN_419; // @[RAM_ST.scala 31:71]
  assign _GEN_421 = 11'h1a5 == WADDR ? 11'h1a5 : _GEN_420; // @[RAM_ST.scala 31:71]
  assign _GEN_422 = 11'h1a6 == WADDR ? 11'h1a6 : _GEN_421; // @[RAM_ST.scala 31:71]
  assign _GEN_423 = 11'h1a7 == WADDR ? 11'h1a7 : _GEN_422; // @[RAM_ST.scala 31:71]
  assign _GEN_424 = 11'h1a8 == WADDR ? 11'h1a8 : _GEN_423; // @[RAM_ST.scala 31:71]
  assign _GEN_425 = 11'h1a9 == WADDR ? 11'h1a9 : _GEN_424; // @[RAM_ST.scala 31:71]
  assign _GEN_426 = 11'h1aa == WADDR ? 11'h1aa : _GEN_425; // @[RAM_ST.scala 31:71]
  assign _GEN_427 = 11'h1ab == WADDR ? 11'h1ab : _GEN_426; // @[RAM_ST.scala 31:71]
  assign _GEN_428 = 11'h1ac == WADDR ? 11'h1ac : _GEN_427; // @[RAM_ST.scala 31:71]
  assign _GEN_429 = 11'h1ad == WADDR ? 11'h1ad : _GEN_428; // @[RAM_ST.scala 31:71]
  assign _GEN_430 = 11'h1ae == WADDR ? 11'h1ae : _GEN_429; // @[RAM_ST.scala 31:71]
  assign _GEN_431 = 11'h1af == WADDR ? 11'h1af : _GEN_430; // @[RAM_ST.scala 31:71]
  assign _GEN_432 = 11'h1b0 == WADDR ? 11'h1b0 : _GEN_431; // @[RAM_ST.scala 31:71]
  assign _GEN_433 = 11'h1b1 == WADDR ? 11'h1b1 : _GEN_432; // @[RAM_ST.scala 31:71]
  assign _GEN_434 = 11'h1b2 == WADDR ? 11'h1b2 : _GEN_433; // @[RAM_ST.scala 31:71]
  assign _GEN_435 = 11'h1b3 == WADDR ? 11'h1b3 : _GEN_434; // @[RAM_ST.scala 31:71]
  assign _GEN_436 = 11'h1b4 == WADDR ? 11'h1b4 : _GEN_435; // @[RAM_ST.scala 31:71]
  assign _GEN_437 = 11'h1b5 == WADDR ? 11'h1b5 : _GEN_436; // @[RAM_ST.scala 31:71]
  assign _GEN_438 = 11'h1b6 == WADDR ? 11'h1b6 : _GEN_437; // @[RAM_ST.scala 31:71]
  assign _GEN_439 = 11'h1b7 == WADDR ? 11'h1b7 : _GEN_438; // @[RAM_ST.scala 31:71]
  assign _GEN_440 = 11'h1b8 == WADDR ? 11'h1b8 : _GEN_439; // @[RAM_ST.scala 31:71]
  assign _GEN_441 = 11'h1b9 == WADDR ? 11'h1b9 : _GEN_440; // @[RAM_ST.scala 31:71]
  assign _GEN_442 = 11'h1ba == WADDR ? 11'h1ba : _GEN_441; // @[RAM_ST.scala 31:71]
  assign _GEN_443 = 11'h1bb == WADDR ? 11'h1bb : _GEN_442; // @[RAM_ST.scala 31:71]
  assign _GEN_444 = 11'h1bc == WADDR ? 11'h1bc : _GEN_443; // @[RAM_ST.scala 31:71]
  assign _GEN_445 = 11'h1bd == WADDR ? 11'h1bd : _GEN_444; // @[RAM_ST.scala 31:71]
  assign _GEN_446 = 11'h1be == WADDR ? 11'h1be : _GEN_445; // @[RAM_ST.scala 31:71]
  assign _GEN_447 = 11'h1bf == WADDR ? 11'h1bf : _GEN_446; // @[RAM_ST.scala 31:71]
  assign _GEN_448 = 11'h1c0 == WADDR ? 11'h1c0 : _GEN_447; // @[RAM_ST.scala 31:71]
  assign _GEN_449 = 11'h1c1 == WADDR ? 11'h1c1 : _GEN_448; // @[RAM_ST.scala 31:71]
  assign _GEN_450 = 11'h1c2 == WADDR ? 11'h1c2 : _GEN_449; // @[RAM_ST.scala 31:71]
  assign _GEN_451 = 11'h1c3 == WADDR ? 11'h1c3 : _GEN_450; // @[RAM_ST.scala 31:71]
  assign _GEN_452 = 11'h1c4 == WADDR ? 11'h1c4 : _GEN_451; // @[RAM_ST.scala 31:71]
  assign _GEN_453 = 11'h1c5 == WADDR ? 11'h1c5 : _GEN_452; // @[RAM_ST.scala 31:71]
  assign _GEN_454 = 11'h1c6 == WADDR ? 11'h1c6 : _GEN_453; // @[RAM_ST.scala 31:71]
  assign _GEN_455 = 11'h1c7 == WADDR ? 11'h1c7 : _GEN_454; // @[RAM_ST.scala 31:71]
  assign _GEN_456 = 11'h1c8 == WADDR ? 11'h1c8 : _GEN_455; // @[RAM_ST.scala 31:71]
  assign _GEN_457 = 11'h1c9 == WADDR ? 11'h1c9 : _GEN_456; // @[RAM_ST.scala 31:71]
  assign _GEN_458 = 11'h1ca == WADDR ? 11'h1ca : _GEN_457; // @[RAM_ST.scala 31:71]
  assign _GEN_459 = 11'h1cb == WADDR ? 11'h1cb : _GEN_458; // @[RAM_ST.scala 31:71]
  assign _GEN_460 = 11'h1cc == WADDR ? 11'h1cc : _GEN_459; // @[RAM_ST.scala 31:71]
  assign _GEN_461 = 11'h1cd == WADDR ? 11'h1cd : _GEN_460; // @[RAM_ST.scala 31:71]
  assign _GEN_462 = 11'h1ce == WADDR ? 11'h1ce : _GEN_461; // @[RAM_ST.scala 31:71]
  assign _GEN_463 = 11'h1cf == WADDR ? 11'h1cf : _GEN_462; // @[RAM_ST.scala 31:71]
  assign _GEN_464 = 11'h1d0 == WADDR ? 11'h1d0 : _GEN_463; // @[RAM_ST.scala 31:71]
  assign _GEN_465 = 11'h1d1 == WADDR ? 11'h1d1 : _GEN_464; // @[RAM_ST.scala 31:71]
  assign _GEN_466 = 11'h1d2 == WADDR ? 11'h1d2 : _GEN_465; // @[RAM_ST.scala 31:71]
  assign _GEN_467 = 11'h1d3 == WADDR ? 11'h1d3 : _GEN_466; // @[RAM_ST.scala 31:71]
  assign _GEN_468 = 11'h1d4 == WADDR ? 11'h1d4 : _GEN_467; // @[RAM_ST.scala 31:71]
  assign _GEN_469 = 11'h1d5 == WADDR ? 11'h1d5 : _GEN_468; // @[RAM_ST.scala 31:71]
  assign _GEN_470 = 11'h1d6 == WADDR ? 11'h1d6 : _GEN_469; // @[RAM_ST.scala 31:71]
  assign _GEN_471 = 11'h1d7 == WADDR ? 11'h1d7 : _GEN_470; // @[RAM_ST.scala 31:71]
  assign _GEN_472 = 11'h1d8 == WADDR ? 11'h1d8 : _GEN_471; // @[RAM_ST.scala 31:71]
  assign _GEN_473 = 11'h1d9 == WADDR ? 11'h1d9 : _GEN_472; // @[RAM_ST.scala 31:71]
  assign _GEN_474 = 11'h1da == WADDR ? 11'h1da : _GEN_473; // @[RAM_ST.scala 31:71]
  assign _GEN_475 = 11'h1db == WADDR ? 11'h1db : _GEN_474; // @[RAM_ST.scala 31:71]
  assign _GEN_476 = 11'h1dc == WADDR ? 11'h1dc : _GEN_475; // @[RAM_ST.scala 31:71]
  assign _GEN_477 = 11'h1dd == WADDR ? 11'h1dd : _GEN_476; // @[RAM_ST.scala 31:71]
  assign _GEN_478 = 11'h1de == WADDR ? 11'h1de : _GEN_477; // @[RAM_ST.scala 31:71]
  assign _GEN_479 = 11'h1df == WADDR ? 11'h1df : _GEN_478; // @[RAM_ST.scala 31:71]
  assign _GEN_480 = 11'h1e0 == WADDR ? 11'h1e0 : _GEN_479; // @[RAM_ST.scala 31:71]
  assign _GEN_481 = 11'h1e1 == WADDR ? 11'h1e1 : _GEN_480; // @[RAM_ST.scala 31:71]
  assign _GEN_482 = 11'h1e2 == WADDR ? 11'h1e2 : _GEN_481; // @[RAM_ST.scala 31:71]
  assign _GEN_483 = 11'h1e3 == WADDR ? 11'h1e3 : _GEN_482; // @[RAM_ST.scala 31:71]
  assign _GEN_484 = 11'h1e4 == WADDR ? 11'h1e4 : _GEN_483; // @[RAM_ST.scala 31:71]
  assign _GEN_485 = 11'h1e5 == WADDR ? 11'h1e5 : _GEN_484; // @[RAM_ST.scala 31:71]
  assign _GEN_486 = 11'h1e6 == WADDR ? 11'h1e6 : _GEN_485; // @[RAM_ST.scala 31:71]
  assign _GEN_487 = 11'h1e7 == WADDR ? 11'h1e7 : _GEN_486; // @[RAM_ST.scala 31:71]
  assign _GEN_488 = 11'h1e8 == WADDR ? 11'h1e8 : _GEN_487; // @[RAM_ST.scala 31:71]
  assign _GEN_489 = 11'h1e9 == WADDR ? 11'h1e9 : _GEN_488; // @[RAM_ST.scala 31:71]
  assign _GEN_490 = 11'h1ea == WADDR ? 11'h1ea : _GEN_489; // @[RAM_ST.scala 31:71]
  assign _GEN_491 = 11'h1eb == WADDR ? 11'h1eb : _GEN_490; // @[RAM_ST.scala 31:71]
  assign _GEN_492 = 11'h1ec == WADDR ? 11'h1ec : _GEN_491; // @[RAM_ST.scala 31:71]
  assign _GEN_493 = 11'h1ed == WADDR ? 11'h1ed : _GEN_492; // @[RAM_ST.scala 31:71]
  assign _GEN_494 = 11'h1ee == WADDR ? 11'h1ee : _GEN_493; // @[RAM_ST.scala 31:71]
  assign _GEN_495 = 11'h1ef == WADDR ? 11'h1ef : _GEN_494; // @[RAM_ST.scala 31:71]
  assign _GEN_496 = 11'h1f0 == WADDR ? 11'h1f0 : _GEN_495; // @[RAM_ST.scala 31:71]
  assign _GEN_497 = 11'h1f1 == WADDR ? 11'h1f1 : _GEN_496; // @[RAM_ST.scala 31:71]
  assign _GEN_498 = 11'h1f2 == WADDR ? 11'h1f2 : _GEN_497; // @[RAM_ST.scala 31:71]
  assign _GEN_499 = 11'h1f3 == WADDR ? 11'h1f3 : _GEN_498; // @[RAM_ST.scala 31:71]
  assign _GEN_500 = 11'h1f4 == WADDR ? 11'h1f4 : _GEN_499; // @[RAM_ST.scala 31:71]
  assign _GEN_501 = 11'h1f5 == WADDR ? 11'h1f5 : _GEN_500; // @[RAM_ST.scala 31:71]
  assign _GEN_502 = 11'h1f6 == WADDR ? 11'h1f6 : _GEN_501; // @[RAM_ST.scala 31:71]
  assign _GEN_503 = 11'h1f7 == WADDR ? 11'h1f7 : _GEN_502; // @[RAM_ST.scala 31:71]
  assign _GEN_504 = 11'h1f8 == WADDR ? 11'h1f8 : _GEN_503; // @[RAM_ST.scala 31:71]
  assign _GEN_505 = 11'h1f9 == WADDR ? 11'h1f9 : _GEN_504; // @[RAM_ST.scala 31:71]
  assign _GEN_506 = 11'h1fa == WADDR ? 11'h1fa : _GEN_505; // @[RAM_ST.scala 31:71]
  assign _GEN_507 = 11'h1fb == WADDR ? 11'h1fb : _GEN_506; // @[RAM_ST.scala 31:71]
  assign _GEN_508 = 11'h1fc == WADDR ? 11'h1fc : _GEN_507; // @[RAM_ST.scala 31:71]
  assign _GEN_509 = 11'h1fd == WADDR ? 11'h1fd : _GEN_508; // @[RAM_ST.scala 31:71]
  assign _GEN_510 = 11'h1fe == WADDR ? 11'h1fe : _GEN_509; // @[RAM_ST.scala 31:71]
  assign _GEN_511 = 11'h1ff == WADDR ? 11'h1ff : _GEN_510; // @[RAM_ST.scala 31:71]
  assign _GEN_512 = 11'h200 == WADDR ? 11'h200 : _GEN_511; // @[RAM_ST.scala 31:71]
  assign _GEN_513 = 11'h201 == WADDR ? 11'h201 : _GEN_512; // @[RAM_ST.scala 31:71]
  assign _GEN_514 = 11'h202 == WADDR ? 11'h202 : _GEN_513; // @[RAM_ST.scala 31:71]
  assign _GEN_515 = 11'h203 == WADDR ? 11'h203 : _GEN_514; // @[RAM_ST.scala 31:71]
  assign _GEN_516 = 11'h204 == WADDR ? 11'h204 : _GEN_515; // @[RAM_ST.scala 31:71]
  assign _GEN_517 = 11'h205 == WADDR ? 11'h205 : _GEN_516; // @[RAM_ST.scala 31:71]
  assign _GEN_518 = 11'h206 == WADDR ? 11'h206 : _GEN_517; // @[RAM_ST.scala 31:71]
  assign _GEN_519 = 11'h207 == WADDR ? 11'h207 : _GEN_518; // @[RAM_ST.scala 31:71]
  assign _GEN_520 = 11'h208 == WADDR ? 11'h208 : _GEN_519; // @[RAM_ST.scala 31:71]
  assign _GEN_521 = 11'h209 == WADDR ? 11'h209 : _GEN_520; // @[RAM_ST.scala 31:71]
  assign _GEN_522 = 11'h20a == WADDR ? 11'h20a : _GEN_521; // @[RAM_ST.scala 31:71]
  assign _GEN_523 = 11'h20b == WADDR ? 11'h20b : _GEN_522; // @[RAM_ST.scala 31:71]
  assign _GEN_524 = 11'h20c == WADDR ? 11'h20c : _GEN_523; // @[RAM_ST.scala 31:71]
  assign _GEN_525 = 11'h20d == WADDR ? 11'h20d : _GEN_524; // @[RAM_ST.scala 31:71]
  assign _GEN_526 = 11'h20e == WADDR ? 11'h20e : _GEN_525; // @[RAM_ST.scala 31:71]
  assign _GEN_527 = 11'h20f == WADDR ? 11'h20f : _GEN_526; // @[RAM_ST.scala 31:71]
  assign _GEN_528 = 11'h210 == WADDR ? 11'h210 : _GEN_527; // @[RAM_ST.scala 31:71]
  assign _GEN_529 = 11'h211 == WADDR ? 11'h211 : _GEN_528; // @[RAM_ST.scala 31:71]
  assign _GEN_530 = 11'h212 == WADDR ? 11'h212 : _GEN_529; // @[RAM_ST.scala 31:71]
  assign _GEN_531 = 11'h213 == WADDR ? 11'h213 : _GEN_530; // @[RAM_ST.scala 31:71]
  assign _GEN_532 = 11'h214 == WADDR ? 11'h214 : _GEN_531; // @[RAM_ST.scala 31:71]
  assign _GEN_533 = 11'h215 == WADDR ? 11'h215 : _GEN_532; // @[RAM_ST.scala 31:71]
  assign _GEN_534 = 11'h216 == WADDR ? 11'h216 : _GEN_533; // @[RAM_ST.scala 31:71]
  assign _GEN_535 = 11'h217 == WADDR ? 11'h217 : _GEN_534; // @[RAM_ST.scala 31:71]
  assign _GEN_536 = 11'h218 == WADDR ? 11'h218 : _GEN_535; // @[RAM_ST.scala 31:71]
  assign _GEN_537 = 11'h219 == WADDR ? 11'h219 : _GEN_536; // @[RAM_ST.scala 31:71]
  assign _GEN_538 = 11'h21a == WADDR ? 11'h21a : _GEN_537; // @[RAM_ST.scala 31:71]
  assign _GEN_539 = 11'h21b == WADDR ? 11'h21b : _GEN_538; // @[RAM_ST.scala 31:71]
  assign _GEN_540 = 11'h21c == WADDR ? 11'h21c : _GEN_539; // @[RAM_ST.scala 31:71]
  assign _GEN_541 = 11'h21d == WADDR ? 11'h21d : _GEN_540; // @[RAM_ST.scala 31:71]
  assign _GEN_542 = 11'h21e == WADDR ? 11'h21e : _GEN_541; // @[RAM_ST.scala 31:71]
  assign _GEN_543 = 11'h21f == WADDR ? 11'h21f : _GEN_542; // @[RAM_ST.scala 31:71]
  assign _GEN_544 = 11'h220 == WADDR ? 11'h220 : _GEN_543; // @[RAM_ST.scala 31:71]
  assign _GEN_545 = 11'h221 == WADDR ? 11'h221 : _GEN_544; // @[RAM_ST.scala 31:71]
  assign _GEN_546 = 11'h222 == WADDR ? 11'h222 : _GEN_545; // @[RAM_ST.scala 31:71]
  assign _GEN_547 = 11'h223 == WADDR ? 11'h223 : _GEN_546; // @[RAM_ST.scala 31:71]
  assign _GEN_548 = 11'h224 == WADDR ? 11'h224 : _GEN_547; // @[RAM_ST.scala 31:71]
  assign _GEN_549 = 11'h225 == WADDR ? 11'h225 : _GEN_548; // @[RAM_ST.scala 31:71]
  assign _GEN_550 = 11'h226 == WADDR ? 11'h226 : _GEN_549; // @[RAM_ST.scala 31:71]
  assign _GEN_551 = 11'h227 == WADDR ? 11'h227 : _GEN_550; // @[RAM_ST.scala 31:71]
  assign _GEN_552 = 11'h228 == WADDR ? 11'h228 : _GEN_551; // @[RAM_ST.scala 31:71]
  assign _GEN_553 = 11'h229 == WADDR ? 11'h229 : _GEN_552; // @[RAM_ST.scala 31:71]
  assign _GEN_554 = 11'h22a == WADDR ? 11'h22a : _GEN_553; // @[RAM_ST.scala 31:71]
  assign _GEN_555 = 11'h22b == WADDR ? 11'h22b : _GEN_554; // @[RAM_ST.scala 31:71]
  assign _GEN_556 = 11'h22c == WADDR ? 11'h22c : _GEN_555; // @[RAM_ST.scala 31:71]
  assign _GEN_557 = 11'h22d == WADDR ? 11'h22d : _GEN_556; // @[RAM_ST.scala 31:71]
  assign _GEN_558 = 11'h22e == WADDR ? 11'h22e : _GEN_557; // @[RAM_ST.scala 31:71]
  assign _GEN_559 = 11'h22f == WADDR ? 11'h22f : _GEN_558; // @[RAM_ST.scala 31:71]
  assign _GEN_560 = 11'h230 == WADDR ? 11'h230 : _GEN_559; // @[RAM_ST.scala 31:71]
  assign _GEN_561 = 11'h231 == WADDR ? 11'h231 : _GEN_560; // @[RAM_ST.scala 31:71]
  assign _GEN_562 = 11'h232 == WADDR ? 11'h232 : _GEN_561; // @[RAM_ST.scala 31:71]
  assign _GEN_563 = 11'h233 == WADDR ? 11'h233 : _GEN_562; // @[RAM_ST.scala 31:71]
  assign _GEN_564 = 11'h234 == WADDR ? 11'h234 : _GEN_563; // @[RAM_ST.scala 31:71]
  assign _GEN_565 = 11'h235 == WADDR ? 11'h235 : _GEN_564; // @[RAM_ST.scala 31:71]
  assign _GEN_566 = 11'h236 == WADDR ? 11'h236 : _GEN_565; // @[RAM_ST.scala 31:71]
  assign _GEN_567 = 11'h237 == WADDR ? 11'h237 : _GEN_566; // @[RAM_ST.scala 31:71]
  assign _GEN_568 = 11'h238 == WADDR ? 11'h238 : _GEN_567; // @[RAM_ST.scala 31:71]
  assign _GEN_569 = 11'h239 == WADDR ? 11'h239 : _GEN_568; // @[RAM_ST.scala 31:71]
  assign _GEN_570 = 11'h23a == WADDR ? 11'h23a : _GEN_569; // @[RAM_ST.scala 31:71]
  assign _GEN_571 = 11'h23b == WADDR ? 11'h23b : _GEN_570; // @[RAM_ST.scala 31:71]
  assign _GEN_572 = 11'h23c == WADDR ? 11'h23c : _GEN_571; // @[RAM_ST.scala 31:71]
  assign _GEN_573 = 11'h23d == WADDR ? 11'h23d : _GEN_572; // @[RAM_ST.scala 31:71]
  assign _GEN_574 = 11'h23e == WADDR ? 11'h23e : _GEN_573; // @[RAM_ST.scala 31:71]
  assign _GEN_575 = 11'h23f == WADDR ? 11'h23f : _GEN_574; // @[RAM_ST.scala 31:71]
  assign _GEN_576 = 11'h240 == WADDR ? 11'h240 : _GEN_575; // @[RAM_ST.scala 31:71]
  assign _GEN_577 = 11'h241 == WADDR ? 11'h241 : _GEN_576; // @[RAM_ST.scala 31:71]
  assign _GEN_578 = 11'h242 == WADDR ? 11'h242 : _GEN_577; // @[RAM_ST.scala 31:71]
  assign _GEN_579 = 11'h243 == WADDR ? 11'h243 : _GEN_578; // @[RAM_ST.scala 31:71]
  assign _GEN_580 = 11'h244 == WADDR ? 11'h244 : _GEN_579; // @[RAM_ST.scala 31:71]
  assign _GEN_581 = 11'h245 == WADDR ? 11'h245 : _GEN_580; // @[RAM_ST.scala 31:71]
  assign _GEN_582 = 11'h246 == WADDR ? 11'h246 : _GEN_581; // @[RAM_ST.scala 31:71]
  assign _GEN_583 = 11'h247 == WADDR ? 11'h247 : _GEN_582; // @[RAM_ST.scala 31:71]
  assign _GEN_584 = 11'h248 == WADDR ? 11'h248 : _GEN_583; // @[RAM_ST.scala 31:71]
  assign _GEN_585 = 11'h249 == WADDR ? 11'h249 : _GEN_584; // @[RAM_ST.scala 31:71]
  assign _GEN_586 = 11'h24a == WADDR ? 11'h24a : _GEN_585; // @[RAM_ST.scala 31:71]
  assign _GEN_587 = 11'h24b == WADDR ? 11'h24b : _GEN_586; // @[RAM_ST.scala 31:71]
  assign _GEN_588 = 11'h24c == WADDR ? 11'h24c : _GEN_587; // @[RAM_ST.scala 31:71]
  assign _GEN_589 = 11'h24d == WADDR ? 11'h24d : _GEN_588; // @[RAM_ST.scala 31:71]
  assign _GEN_590 = 11'h24e == WADDR ? 11'h24e : _GEN_589; // @[RAM_ST.scala 31:71]
  assign _GEN_591 = 11'h24f == WADDR ? 11'h24f : _GEN_590; // @[RAM_ST.scala 31:71]
  assign _GEN_592 = 11'h250 == WADDR ? 11'h250 : _GEN_591; // @[RAM_ST.scala 31:71]
  assign _GEN_593 = 11'h251 == WADDR ? 11'h251 : _GEN_592; // @[RAM_ST.scala 31:71]
  assign _GEN_594 = 11'h252 == WADDR ? 11'h252 : _GEN_593; // @[RAM_ST.scala 31:71]
  assign _GEN_595 = 11'h253 == WADDR ? 11'h253 : _GEN_594; // @[RAM_ST.scala 31:71]
  assign _GEN_596 = 11'h254 == WADDR ? 11'h254 : _GEN_595; // @[RAM_ST.scala 31:71]
  assign _GEN_597 = 11'h255 == WADDR ? 11'h255 : _GEN_596; // @[RAM_ST.scala 31:71]
  assign _GEN_598 = 11'h256 == WADDR ? 11'h256 : _GEN_597; // @[RAM_ST.scala 31:71]
  assign _GEN_599 = 11'h257 == WADDR ? 11'h257 : _GEN_598; // @[RAM_ST.scala 31:71]
  assign _GEN_600 = 11'h258 == WADDR ? 11'h258 : _GEN_599; // @[RAM_ST.scala 31:71]
  assign _GEN_601 = 11'h259 == WADDR ? 11'h259 : _GEN_600; // @[RAM_ST.scala 31:71]
  assign _GEN_602 = 11'h25a == WADDR ? 11'h25a : _GEN_601; // @[RAM_ST.scala 31:71]
  assign _GEN_603 = 11'h25b == WADDR ? 11'h25b : _GEN_602; // @[RAM_ST.scala 31:71]
  assign _GEN_604 = 11'h25c == WADDR ? 11'h25c : _GEN_603; // @[RAM_ST.scala 31:71]
  assign _GEN_605 = 11'h25d == WADDR ? 11'h25d : _GEN_604; // @[RAM_ST.scala 31:71]
  assign _GEN_606 = 11'h25e == WADDR ? 11'h25e : _GEN_605; // @[RAM_ST.scala 31:71]
  assign _GEN_607 = 11'h25f == WADDR ? 11'h25f : _GEN_606; // @[RAM_ST.scala 31:71]
  assign _GEN_608 = 11'h260 == WADDR ? 11'h260 : _GEN_607; // @[RAM_ST.scala 31:71]
  assign _GEN_609 = 11'h261 == WADDR ? 11'h261 : _GEN_608; // @[RAM_ST.scala 31:71]
  assign _GEN_610 = 11'h262 == WADDR ? 11'h262 : _GEN_609; // @[RAM_ST.scala 31:71]
  assign _GEN_611 = 11'h263 == WADDR ? 11'h263 : _GEN_610; // @[RAM_ST.scala 31:71]
  assign _GEN_612 = 11'h264 == WADDR ? 11'h264 : _GEN_611; // @[RAM_ST.scala 31:71]
  assign _GEN_613 = 11'h265 == WADDR ? 11'h265 : _GEN_612; // @[RAM_ST.scala 31:71]
  assign _GEN_614 = 11'h266 == WADDR ? 11'h266 : _GEN_613; // @[RAM_ST.scala 31:71]
  assign _GEN_615 = 11'h267 == WADDR ? 11'h267 : _GEN_614; // @[RAM_ST.scala 31:71]
  assign _GEN_616 = 11'h268 == WADDR ? 11'h268 : _GEN_615; // @[RAM_ST.scala 31:71]
  assign _GEN_617 = 11'h269 == WADDR ? 11'h269 : _GEN_616; // @[RAM_ST.scala 31:71]
  assign _GEN_618 = 11'h26a == WADDR ? 11'h26a : _GEN_617; // @[RAM_ST.scala 31:71]
  assign _GEN_619 = 11'h26b == WADDR ? 11'h26b : _GEN_618; // @[RAM_ST.scala 31:71]
  assign _GEN_620 = 11'h26c == WADDR ? 11'h26c : _GEN_619; // @[RAM_ST.scala 31:71]
  assign _GEN_621 = 11'h26d == WADDR ? 11'h26d : _GEN_620; // @[RAM_ST.scala 31:71]
  assign _GEN_622 = 11'h26e == WADDR ? 11'h26e : _GEN_621; // @[RAM_ST.scala 31:71]
  assign _GEN_623 = 11'h26f == WADDR ? 11'h26f : _GEN_622; // @[RAM_ST.scala 31:71]
  assign _GEN_624 = 11'h270 == WADDR ? 11'h270 : _GEN_623; // @[RAM_ST.scala 31:71]
  assign _GEN_625 = 11'h271 == WADDR ? 11'h271 : _GEN_624; // @[RAM_ST.scala 31:71]
  assign _GEN_626 = 11'h272 == WADDR ? 11'h272 : _GEN_625; // @[RAM_ST.scala 31:71]
  assign _GEN_627 = 11'h273 == WADDR ? 11'h273 : _GEN_626; // @[RAM_ST.scala 31:71]
  assign _GEN_628 = 11'h274 == WADDR ? 11'h274 : _GEN_627; // @[RAM_ST.scala 31:71]
  assign _GEN_629 = 11'h275 == WADDR ? 11'h275 : _GEN_628; // @[RAM_ST.scala 31:71]
  assign _GEN_630 = 11'h276 == WADDR ? 11'h276 : _GEN_629; // @[RAM_ST.scala 31:71]
  assign _GEN_631 = 11'h277 == WADDR ? 11'h277 : _GEN_630; // @[RAM_ST.scala 31:71]
  assign _GEN_632 = 11'h278 == WADDR ? 11'h278 : _GEN_631; // @[RAM_ST.scala 31:71]
  assign _GEN_633 = 11'h279 == WADDR ? 11'h279 : _GEN_632; // @[RAM_ST.scala 31:71]
  assign _GEN_634 = 11'h27a == WADDR ? 11'h27a : _GEN_633; // @[RAM_ST.scala 31:71]
  assign _GEN_635 = 11'h27b == WADDR ? 11'h27b : _GEN_634; // @[RAM_ST.scala 31:71]
  assign _GEN_636 = 11'h27c == WADDR ? 11'h27c : _GEN_635; // @[RAM_ST.scala 31:71]
  assign _GEN_637 = 11'h27d == WADDR ? 11'h27d : _GEN_636; // @[RAM_ST.scala 31:71]
  assign _GEN_638 = 11'h27e == WADDR ? 11'h27e : _GEN_637; // @[RAM_ST.scala 31:71]
  assign _GEN_639 = 11'h27f == WADDR ? 11'h27f : _GEN_638; // @[RAM_ST.scala 31:71]
  assign _GEN_640 = 11'h280 == WADDR ? 11'h280 : _GEN_639; // @[RAM_ST.scala 31:71]
  assign _GEN_641 = 11'h281 == WADDR ? 11'h281 : _GEN_640; // @[RAM_ST.scala 31:71]
  assign _GEN_642 = 11'h282 == WADDR ? 11'h282 : _GEN_641; // @[RAM_ST.scala 31:71]
  assign _GEN_643 = 11'h283 == WADDR ? 11'h283 : _GEN_642; // @[RAM_ST.scala 31:71]
  assign _GEN_644 = 11'h284 == WADDR ? 11'h284 : _GEN_643; // @[RAM_ST.scala 31:71]
  assign _GEN_645 = 11'h285 == WADDR ? 11'h285 : _GEN_644; // @[RAM_ST.scala 31:71]
  assign _GEN_646 = 11'h286 == WADDR ? 11'h286 : _GEN_645; // @[RAM_ST.scala 31:71]
  assign _GEN_647 = 11'h287 == WADDR ? 11'h287 : _GEN_646; // @[RAM_ST.scala 31:71]
  assign _GEN_648 = 11'h288 == WADDR ? 11'h288 : _GEN_647; // @[RAM_ST.scala 31:71]
  assign _GEN_649 = 11'h289 == WADDR ? 11'h289 : _GEN_648; // @[RAM_ST.scala 31:71]
  assign _GEN_650 = 11'h28a == WADDR ? 11'h28a : _GEN_649; // @[RAM_ST.scala 31:71]
  assign _GEN_651 = 11'h28b == WADDR ? 11'h28b : _GEN_650; // @[RAM_ST.scala 31:71]
  assign _GEN_652 = 11'h28c == WADDR ? 11'h28c : _GEN_651; // @[RAM_ST.scala 31:71]
  assign _GEN_653 = 11'h28d == WADDR ? 11'h28d : _GEN_652; // @[RAM_ST.scala 31:71]
  assign _GEN_654 = 11'h28e == WADDR ? 11'h28e : _GEN_653; // @[RAM_ST.scala 31:71]
  assign _GEN_655 = 11'h28f == WADDR ? 11'h28f : _GEN_654; // @[RAM_ST.scala 31:71]
  assign _GEN_656 = 11'h290 == WADDR ? 11'h290 : _GEN_655; // @[RAM_ST.scala 31:71]
  assign _GEN_657 = 11'h291 == WADDR ? 11'h291 : _GEN_656; // @[RAM_ST.scala 31:71]
  assign _GEN_658 = 11'h292 == WADDR ? 11'h292 : _GEN_657; // @[RAM_ST.scala 31:71]
  assign _GEN_659 = 11'h293 == WADDR ? 11'h293 : _GEN_658; // @[RAM_ST.scala 31:71]
  assign _GEN_660 = 11'h294 == WADDR ? 11'h294 : _GEN_659; // @[RAM_ST.scala 31:71]
  assign _GEN_661 = 11'h295 == WADDR ? 11'h295 : _GEN_660; // @[RAM_ST.scala 31:71]
  assign _GEN_662 = 11'h296 == WADDR ? 11'h296 : _GEN_661; // @[RAM_ST.scala 31:71]
  assign _GEN_663 = 11'h297 == WADDR ? 11'h297 : _GEN_662; // @[RAM_ST.scala 31:71]
  assign _GEN_664 = 11'h298 == WADDR ? 11'h298 : _GEN_663; // @[RAM_ST.scala 31:71]
  assign _GEN_665 = 11'h299 == WADDR ? 11'h299 : _GEN_664; // @[RAM_ST.scala 31:71]
  assign _GEN_666 = 11'h29a == WADDR ? 11'h29a : _GEN_665; // @[RAM_ST.scala 31:71]
  assign _GEN_667 = 11'h29b == WADDR ? 11'h29b : _GEN_666; // @[RAM_ST.scala 31:71]
  assign _GEN_668 = 11'h29c == WADDR ? 11'h29c : _GEN_667; // @[RAM_ST.scala 31:71]
  assign _GEN_669 = 11'h29d == WADDR ? 11'h29d : _GEN_668; // @[RAM_ST.scala 31:71]
  assign _GEN_670 = 11'h29e == WADDR ? 11'h29e : _GEN_669; // @[RAM_ST.scala 31:71]
  assign _GEN_671 = 11'h29f == WADDR ? 11'h29f : _GEN_670; // @[RAM_ST.scala 31:71]
  assign _GEN_672 = 11'h2a0 == WADDR ? 11'h2a0 : _GEN_671; // @[RAM_ST.scala 31:71]
  assign _GEN_673 = 11'h2a1 == WADDR ? 11'h2a1 : _GEN_672; // @[RAM_ST.scala 31:71]
  assign _GEN_674 = 11'h2a2 == WADDR ? 11'h2a2 : _GEN_673; // @[RAM_ST.scala 31:71]
  assign _GEN_675 = 11'h2a3 == WADDR ? 11'h2a3 : _GEN_674; // @[RAM_ST.scala 31:71]
  assign _GEN_676 = 11'h2a4 == WADDR ? 11'h2a4 : _GEN_675; // @[RAM_ST.scala 31:71]
  assign _GEN_677 = 11'h2a5 == WADDR ? 11'h2a5 : _GEN_676; // @[RAM_ST.scala 31:71]
  assign _GEN_678 = 11'h2a6 == WADDR ? 11'h2a6 : _GEN_677; // @[RAM_ST.scala 31:71]
  assign _GEN_679 = 11'h2a7 == WADDR ? 11'h2a7 : _GEN_678; // @[RAM_ST.scala 31:71]
  assign _GEN_680 = 11'h2a8 == WADDR ? 11'h2a8 : _GEN_679; // @[RAM_ST.scala 31:71]
  assign _GEN_681 = 11'h2a9 == WADDR ? 11'h2a9 : _GEN_680; // @[RAM_ST.scala 31:71]
  assign _GEN_682 = 11'h2aa == WADDR ? 11'h2aa : _GEN_681; // @[RAM_ST.scala 31:71]
  assign _GEN_683 = 11'h2ab == WADDR ? 11'h2ab : _GEN_682; // @[RAM_ST.scala 31:71]
  assign _GEN_684 = 11'h2ac == WADDR ? 11'h2ac : _GEN_683; // @[RAM_ST.scala 31:71]
  assign _GEN_685 = 11'h2ad == WADDR ? 11'h2ad : _GEN_684; // @[RAM_ST.scala 31:71]
  assign _GEN_686 = 11'h2ae == WADDR ? 11'h2ae : _GEN_685; // @[RAM_ST.scala 31:71]
  assign _GEN_687 = 11'h2af == WADDR ? 11'h2af : _GEN_686; // @[RAM_ST.scala 31:71]
  assign _GEN_688 = 11'h2b0 == WADDR ? 11'h2b0 : _GEN_687; // @[RAM_ST.scala 31:71]
  assign _GEN_689 = 11'h2b1 == WADDR ? 11'h2b1 : _GEN_688; // @[RAM_ST.scala 31:71]
  assign _GEN_690 = 11'h2b2 == WADDR ? 11'h2b2 : _GEN_689; // @[RAM_ST.scala 31:71]
  assign _GEN_691 = 11'h2b3 == WADDR ? 11'h2b3 : _GEN_690; // @[RAM_ST.scala 31:71]
  assign _GEN_692 = 11'h2b4 == WADDR ? 11'h2b4 : _GEN_691; // @[RAM_ST.scala 31:71]
  assign _GEN_693 = 11'h2b5 == WADDR ? 11'h2b5 : _GEN_692; // @[RAM_ST.scala 31:71]
  assign _GEN_694 = 11'h2b6 == WADDR ? 11'h2b6 : _GEN_693; // @[RAM_ST.scala 31:71]
  assign _GEN_695 = 11'h2b7 == WADDR ? 11'h2b7 : _GEN_694; // @[RAM_ST.scala 31:71]
  assign _GEN_696 = 11'h2b8 == WADDR ? 11'h2b8 : _GEN_695; // @[RAM_ST.scala 31:71]
  assign _GEN_697 = 11'h2b9 == WADDR ? 11'h2b9 : _GEN_696; // @[RAM_ST.scala 31:71]
  assign _GEN_698 = 11'h2ba == WADDR ? 11'h2ba : _GEN_697; // @[RAM_ST.scala 31:71]
  assign _GEN_699 = 11'h2bb == WADDR ? 11'h2bb : _GEN_698; // @[RAM_ST.scala 31:71]
  assign _GEN_700 = 11'h2bc == WADDR ? 11'h2bc : _GEN_699; // @[RAM_ST.scala 31:71]
  assign _GEN_701 = 11'h2bd == WADDR ? 11'h2bd : _GEN_700; // @[RAM_ST.scala 31:71]
  assign _GEN_702 = 11'h2be == WADDR ? 11'h2be : _GEN_701; // @[RAM_ST.scala 31:71]
  assign _GEN_703 = 11'h2bf == WADDR ? 11'h2bf : _GEN_702; // @[RAM_ST.scala 31:71]
  assign _GEN_704 = 11'h2c0 == WADDR ? 11'h2c0 : _GEN_703; // @[RAM_ST.scala 31:71]
  assign _GEN_705 = 11'h2c1 == WADDR ? 11'h2c1 : _GEN_704; // @[RAM_ST.scala 31:71]
  assign _GEN_706 = 11'h2c2 == WADDR ? 11'h2c2 : _GEN_705; // @[RAM_ST.scala 31:71]
  assign _GEN_707 = 11'h2c3 == WADDR ? 11'h2c3 : _GEN_706; // @[RAM_ST.scala 31:71]
  assign _GEN_708 = 11'h2c4 == WADDR ? 11'h2c4 : _GEN_707; // @[RAM_ST.scala 31:71]
  assign _GEN_709 = 11'h2c5 == WADDR ? 11'h2c5 : _GEN_708; // @[RAM_ST.scala 31:71]
  assign _GEN_710 = 11'h2c6 == WADDR ? 11'h2c6 : _GEN_709; // @[RAM_ST.scala 31:71]
  assign _GEN_711 = 11'h2c7 == WADDR ? 11'h2c7 : _GEN_710; // @[RAM_ST.scala 31:71]
  assign _GEN_712 = 11'h2c8 == WADDR ? 11'h2c8 : _GEN_711; // @[RAM_ST.scala 31:71]
  assign _GEN_713 = 11'h2c9 == WADDR ? 11'h2c9 : _GEN_712; // @[RAM_ST.scala 31:71]
  assign _GEN_714 = 11'h2ca == WADDR ? 11'h2ca : _GEN_713; // @[RAM_ST.scala 31:71]
  assign _GEN_715 = 11'h2cb == WADDR ? 11'h2cb : _GEN_714; // @[RAM_ST.scala 31:71]
  assign _GEN_716 = 11'h2cc == WADDR ? 11'h2cc : _GEN_715; // @[RAM_ST.scala 31:71]
  assign _GEN_717 = 11'h2cd == WADDR ? 11'h2cd : _GEN_716; // @[RAM_ST.scala 31:71]
  assign _GEN_718 = 11'h2ce == WADDR ? 11'h2ce : _GEN_717; // @[RAM_ST.scala 31:71]
  assign _GEN_719 = 11'h2cf == WADDR ? 11'h2cf : _GEN_718; // @[RAM_ST.scala 31:71]
  assign _GEN_720 = 11'h2d0 == WADDR ? 11'h2d0 : _GEN_719; // @[RAM_ST.scala 31:71]
  assign _GEN_721 = 11'h2d1 == WADDR ? 11'h2d1 : _GEN_720; // @[RAM_ST.scala 31:71]
  assign _GEN_722 = 11'h2d2 == WADDR ? 11'h2d2 : _GEN_721; // @[RAM_ST.scala 31:71]
  assign _GEN_723 = 11'h2d3 == WADDR ? 11'h2d3 : _GEN_722; // @[RAM_ST.scala 31:71]
  assign _GEN_724 = 11'h2d4 == WADDR ? 11'h2d4 : _GEN_723; // @[RAM_ST.scala 31:71]
  assign _GEN_725 = 11'h2d5 == WADDR ? 11'h2d5 : _GEN_724; // @[RAM_ST.scala 31:71]
  assign _GEN_726 = 11'h2d6 == WADDR ? 11'h2d6 : _GEN_725; // @[RAM_ST.scala 31:71]
  assign _GEN_727 = 11'h2d7 == WADDR ? 11'h2d7 : _GEN_726; // @[RAM_ST.scala 31:71]
  assign _GEN_728 = 11'h2d8 == WADDR ? 11'h2d8 : _GEN_727; // @[RAM_ST.scala 31:71]
  assign _GEN_729 = 11'h2d9 == WADDR ? 11'h2d9 : _GEN_728; // @[RAM_ST.scala 31:71]
  assign _GEN_730 = 11'h2da == WADDR ? 11'h2da : _GEN_729; // @[RAM_ST.scala 31:71]
  assign _GEN_731 = 11'h2db == WADDR ? 11'h2db : _GEN_730; // @[RAM_ST.scala 31:71]
  assign _GEN_732 = 11'h2dc == WADDR ? 11'h2dc : _GEN_731; // @[RAM_ST.scala 31:71]
  assign _GEN_733 = 11'h2dd == WADDR ? 11'h2dd : _GEN_732; // @[RAM_ST.scala 31:71]
  assign _GEN_734 = 11'h2de == WADDR ? 11'h2de : _GEN_733; // @[RAM_ST.scala 31:71]
  assign _GEN_735 = 11'h2df == WADDR ? 11'h2df : _GEN_734; // @[RAM_ST.scala 31:71]
  assign _GEN_736 = 11'h2e0 == WADDR ? 11'h2e0 : _GEN_735; // @[RAM_ST.scala 31:71]
  assign _GEN_737 = 11'h2e1 == WADDR ? 11'h2e1 : _GEN_736; // @[RAM_ST.scala 31:71]
  assign _GEN_738 = 11'h2e2 == WADDR ? 11'h2e2 : _GEN_737; // @[RAM_ST.scala 31:71]
  assign _GEN_739 = 11'h2e3 == WADDR ? 11'h2e3 : _GEN_738; // @[RAM_ST.scala 31:71]
  assign _GEN_740 = 11'h2e4 == WADDR ? 11'h2e4 : _GEN_739; // @[RAM_ST.scala 31:71]
  assign _GEN_741 = 11'h2e5 == WADDR ? 11'h2e5 : _GEN_740; // @[RAM_ST.scala 31:71]
  assign _GEN_742 = 11'h2e6 == WADDR ? 11'h2e6 : _GEN_741; // @[RAM_ST.scala 31:71]
  assign _GEN_743 = 11'h2e7 == WADDR ? 11'h2e7 : _GEN_742; // @[RAM_ST.scala 31:71]
  assign _GEN_744 = 11'h2e8 == WADDR ? 11'h2e8 : _GEN_743; // @[RAM_ST.scala 31:71]
  assign _GEN_745 = 11'h2e9 == WADDR ? 11'h2e9 : _GEN_744; // @[RAM_ST.scala 31:71]
  assign _GEN_746 = 11'h2ea == WADDR ? 11'h2ea : _GEN_745; // @[RAM_ST.scala 31:71]
  assign _GEN_747 = 11'h2eb == WADDR ? 11'h2eb : _GEN_746; // @[RAM_ST.scala 31:71]
  assign _GEN_748 = 11'h2ec == WADDR ? 11'h2ec : _GEN_747; // @[RAM_ST.scala 31:71]
  assign _GEN_749 = 11'h2ed == WADDR ? 11'h2ed : _GEN_748; // @[RAM_ST.scala 31:71]
  assign _GEN_750 = 11'h2ee == WADDR ? 11'h2ee : _GEN_749; // @[RAM_ST.scala 31:71]
  assign _GEN_751 = 11'h2ef == WADDR ? 11'h2ef : _GEN_750; // @[RAM_ST.scala 31:71]
  assign _GEN_752 = 11'h2f0 == WADDR ? 11'h2f0 : _GEN_751; // @[RAM_ST.scala 31:71]
  assign _GEN_753 = 11'h2f1 == WADDR ? 11'h2f1 : _GEN_752; // @[RAM_ST.scala 31:71]
  assign _GEN_754 = 11'h2f2 == WADDR ? 11'h2f2 : _GEN_753; // @[RAM_ST.scala 31:71]
  assign _GEN_755 = 11'h2f3 == WADDR ? 11'h2f3 : _GEN_754; // @[RAM_ST.scala 31:71]
  assign _GEN_756 = 11'h2f4 == WADDR ? 11'h2f4 : _GEN_755; // @[RAM_ST.scala 31:71]
  assign _GEN_757 = 11'h2f5 == WADDR ? 11'h2f5 : _GEN_756; // @[RAM_ST.scala 31:71]
  assign _GEN_758 = 11'h2f6 == WADDR ? 11'h2f6 : _GEN_757; // @[RAM_ST.scala 31:71]
  assign _GEN_759 = 11'h2f7 == WADDR ? 11'h2f7 : _GEN_758; // @[RAM_ST.scala 31:71]
  assign _GEN_760 = 11'h2f8 == WADDR ? 11'h2f8 : _GEN_759; // @[RAM_ST.scala 31:71]
  assign _GEN_761 = 11'h2f9 == WADDR ? 11'h2f9 : _GEN_760; // @[RAM_ST.scala 31:71]
  assign _GEN_762 = 11'h2fa == WADDR ? 11'h2fa : _GEN_761; // @[RAM_ST.scala 31:71]
  assign _GEN_763 = 11'h2fb == WADDR ? 11'h2fb : _GEN_762; // @[RAM_ST.scala 31:71]
  assign _GEN_764 = 11'h2fc == WADDR ? 11'h2fc : _GEN_763; // @[RAM_ST.scala 31:71]
  assign _GEN_765 = 11'h2fd == WADDR ? 11'h2fd : _GEN_764; // @[RAM_ST.scala 31:71]
  assign _GEN_766 = 11'h2fe == WADDR ? 11'h2fe : _GEN_765; // @[RAM_ST.scala 31:71]
  assign _GEN_767 = 11'h2ff == WADDR ? 11'h2ff : _GEN_766; // @[RAM_ST.scala 31:71]
  assign _GEN_768 = 11'h300 == WADDR ? 11'h300 : _GEN_767; // @[RAM_ST.scala 31:71]
  assign _GEN_769 = 11'h301 == WADDR ? 11'h301 : _GEN_768; // @[RAM_ST.scala 31:71]
  assign _GEN_770 = 11'h302 == WADDR ? 11'h302 : _GEN_769; // @[RAM_ST.scala 31:71]
  assign _GEN_771 = 11'h303 == WADDR ? 11'h303 : _GEN_770; // @[RAM_ST.scala 31:71]
  assign _GEN_772 = 11'h304 == WADDR ? 11'h304 : _GEN_771; // @[RAM_ST.scala 31:71]
  assign _GEN_773 = 11'h305 == WADDR ? 11'h305 : _GEN_772; // @[RAM_ST.scala 31:71]
  assign _GEN_774 = 11'h306 == WADDR ? 11'h306 : _GEN_773; // @[RAM_ST.scala 31:71]
  assign _GEN_775 = 11'h307 == WADDR ? 11'h307 : _GEN_774; // @[RAM_ST.scala 31:71]
  assign _GEN_776 = 11'h308 == WADDR ? 11'h308 : _GEN_775; // @[RAM_ST.scala 31:71]
  assign _GEN_777 = 11'h309 == WADDR ? 11'h309 : _GEN_776; // @[RAM_ST.scala 31:71]
  assign _GEN_778 = 11'h30a == WADDR ? 11'h30a : _GEN_777; // @[RAM_ST.scala 31:71]
  assign _GEN_779 = 11'h30b == WADDR ? 11'h30b : _GEN_778; // @[RAM_ST.scala 31:71]
  assign _GEN_780 = 11'h30c == WADDR ? 11'h30c : _GEN_779; // @[RAM_ST.scala 31:71]
  assign _GEN_781 = 11'h30d == WADDR ? 11'h30d : _GEN_780; // @[RAM_ST.scala 31:71]
  assign _GEN_782 = 11'h30e == WADDR ? 11'h30e : _GEN_781; // @[RAM_ST.scala 31:71]
  assign _GEN_783 = 11'h30f == WADDR ? 11'h30f : _GEN_782; // @[RAM_ST.scala 31:71]
  assign _GEN_784 = 11'h310 == WADDR ? 11'h310 : _GEN_783; // @[RAM_ST.scala 31:71]
  assign _GEN_785 = 11'h311 == WADDR ? 11'h311 : _GEN_784; // @[RAM_ST.scala 31:71]
  assign _GEN_786 = 11'h312 == WADDR ? 11'h312 : _GEN_785; // @[RAM_ST.scala 31:71]
  assign _GEN_787 = 11'h313 == WADDR ? 11'h313 : _GEN_786; // @[RAM_ST.scala 31:71]
  assign _GEN_788 = 11'h314 == WADDR ? 11'h314 : _GEN_787; // @[RAM_ST.scala 31:71]
  assign _GEN_789 = 11'h315 == WADDR ? 11'h315 : _GEN_788; // @[RAM_ST.scala 31:71]
  assign _GEN_790 = 11'h316 == WADDR ? 11'h316 : _GEN_789; // @[RAM_ST.scala 31:71]
  assign _GEN_791 = 11'h317 == WADDR ? 11'h317 : _GEN_790; // @[RAM_ST.scala 31:71]
  assign _GEN_792 = 11'h318 == WADDR ? 11'h318 : _GEN_791; // @[RAM_ST.scala 31:71]
  assign _GEN_793 = 11'h319 == WADDR ? 11'h319 : _GEN_792; // @[RAM_ST.scala 31:71]
  assign _GEN_794 = 11'h31a == WADDR ? 11'h31a : _GEN_793; // @[RAM_ST.scala 31:71]
  assign _GEN_795 = 11'h31b == WADDR ? 11'h31b : _GEN_794; // @[RAM_ST.scala 31:71]
  assign _GEN_796 = 11'h31c == WADDR ? 11'h31c : _GEN_795; // @[RAM_ST.scala 31:71]
  assign _GEN_797 = 11'h31d == WADDR ? 11'h31d : _GEN_796; // @[RAM_ST.scala 31:71]
  assign _GEN_798 = 11'h31e == WADDR ? 11'h31e : _GEN_797; // @[RAM_ST.scala 31:71]
  assign _GEN_799 = 11'h31f == WADDR ? 11'h31f : _GEN_798; // @[RAM_ST.scala 31:71]
  assign _GEN_800 = 11'h320 == WADDR ? 11'h320 : _GEN_799; // @[RAM_ST.scala 31:71]
  assign _GEN_801 = 11'h321 == WADDR ? 11'h321 : _GEN_800; // @[RAM_ST.scala 31:71]
  assign _GEN_802 = 11'h322 == WADDR ? 11'h322 : _GEN_801; // @[RAM_ST.scala 31:71]
  assign _GEN_803 = 11'h323 == WADDR ? 11'h323 : _GEN_802; // @[RAM_ST.scala 31:71]
  assign _GEN_804 = 11'h324 == WADDR ? 11'h324 : _GEN_803; // @[RAM_ST.scala 31:71]
  assign _GEN_805 = 11'h325 == WADDR ? 11'h325 : _GEN_804; // @[RAM_ST.scala 31:71]
  assign _GEN_806 = 11'h326 == WADDR ? 11'h326 : _GEN_805; // @[RAM_ST.scala 31:71]
  assign _GEN_807 = 11'h327 == WADDR ? 11'h327 : _GEN_806; // @[RAM_ST.scala 31:71]
  assign _GEN_808 = 11'h328 == WADDR ? 11'h328 : _GEN_807; // @[RAM_ST.scala 31:71]
  assign _GEN_809 = 11'h329 == WADDR ? 11'h329 : _GEN_808; // @[RAM_ST.scala 31:71]
  assign _GEN_810 = 11'h32a == WADDR ? 11'h32a : _GEN_809; // @[RAM_ST.scala 31:71]
  assign _GEN_811 = 11'h32b == WADDR ? 11'h32b : _GEN_810; // @[RAM_ST.scala 31:71]
  assign _GEN_812 = 11'h32c == WADDR ? 11'h32c : _GEN_811; // @[RAM_ST.scala 31:71]
  assign _GEN_813 = 11'h32d == WADDR ? 11'h32d : _GEN_812; // @[RAM_ST.scala 31:71]
  assign _GEN_814 = 11'h32e == WADDR ? 11'h32e : _GEN_813; // @[RAM_ST.scala 31:71]
  assign _GEN_815 = 11'h32f == WADDR ? 11'h32f : _GEN_814; // @[RAM_ST.scala 31:71]
  assign _GEN_816 = 11'h330 == WADDR ? 11'h330 : _GEN_815; // @[RAM_ST.scala 31:71]
  assign _GEN_817 = 11'h331 == WADDR ? 11'h331 : _GEN_816; // @[RAM_ST.scala 31:71]
  assign _GEN_818 = 11'h332 == WADDR ? 11'h332 : _GEN_817; // @[RAM_ST.scala 31:71]
  assign _GEN_819 = 11'h333 == WADDR ? 11'h333 : _GEN_818; // @[RAM_ST.scala 31:71]
  assign _GEN_820 = 11'h334 == WADDR ? 11'h334 : _GEN_819; // @[RAM_ST.scala 31:71]
  assign _GEN_821 = 11'h335 == WADDR ? 11'h335 : _GEN_820; // @[RAM_ST.scala 31:71]
  assign _GEN_822 = 11'h336 == WADDR ? 11'h336 : _GEN_821; // @[RAM_ST.scala 31:71]
  assign _GEN_823 = 11'h337 == WADDR ? 11'h337 : _GEN_822; // @[RAM_ST.scala 31:71]
  assign _GEN_824 = 11'h338 == WADDR ? 11'h338 : _GEN_823; // @[RAM_ST.scala 31:71]
  assign _GEN_825 = 11'h339 == WADDR ? 11'h339 : _GEN_824; // @[RAM_ST.scala 31:71]
  assign _GEN_826 = 11'h33a == WADDR ? 11'h33a : _GEN_825; // @[RAM_ST.scala 31:71]
  assign _GEN_827 = 11'h33b == WADDR ? 11'h33b : _GEN_826; // @[RAM_ST.scala 31:71]
  assign _GEN_828 = 11'h33c == WADDR ? 11'h33c : _GEN_827; // @[RAM_ST.scala 31:71]
  assign _GEN_829 = 11'h33d == WADDR ? 11'h33d : _GEN_828; // @[RAM_ST.scala 31:71]
  assign _GEN_830 = 11'h33e == WADDR ? 11'h33e : _GEN_829; // @[RAM_ST.scala 31:71]
  assign _GEN_831 = 11'h33f == WADDR ? 11'h33f : _GEN_830; // @[RAM_ST.scala 31:71]
  assign _GEN_832 = 11'h340 == WADDR ? 11'h340 : _GEN_831; // @[RAM_ST.scala 31:71]
  assign _GEN_833 = 11'h341 == WADDR ? 11'h341 : _GEN_832; // @[RAM_ST.scala 31:71]
  assign _GEN_834 = 11'h342 == WADDR ? 11'h342 : _GEN_833; // @[RAM_ST.scala 31:71]
  assign _GEN_835 = 11'h343 == WADDR ? 11'h343 : _GEN_834; // @[RAM_ST.scala 31:71]
  assign _GEN_836 = 11'h344 == WADDR ? 11'h344 : _GEN_835; // @[RAM_ST.scala 31:71]
  assign _GEN_837 = 11'h345 == WADDR ? 11'h345 : _GEN_836; // @[RAM_ST.scala 31:71]
  assign _GEN_838 = 11'h346 == WADDR ? 11'h346 : _GEN_837; // @[RAM_ST.scala 31:71]
  assign _GEN_839 = 11'h347 == WADDR ? 11'h347 : _GEN_838; // @[RAM_ST.scala 31:71]
  assign _GEN_840 = 11'h348 == WADDR ? 11'h348 : _GEN_839; // @[RAM_ST.scala 31:71]
  assign _GEN_841 = 11'h349 == WADDR ? 11'h349 : _GEN_840; // @[RAM_ST.scala 31:71]
  assign _GEN_842 = 11'h34a == WADDR ? 11'h34a : _GEN_841; // @[RAM_ST.scala 31:71]
  assign _GEN_843 = 11'h34b == WADDR ? 11'h34b : _GEN_842; // @[RAM_ST.scala 31:71]
  assign _GEN_844 = 11'h34c == WADDR ? 11'h34c : _GEN_843; // @[RAM_ST.scala 31:71]
  assign _GEN_845 = 11'h34d == WADDR ? 11'h34d : _GEN_844; // @[RAM_ST.scala 31:71]
  assign _GEN_846 = 11'h34e == WADDR ? 11'h34e : _GEN_845; // @[RAM_ST.scala 31:71]
  assign _GEN_847 = 11'h34f == WADDR ? 11'h34f : _GEN_846; // @[RAM_ST.scala 31:71]
  assign _GEN_848 = 11'h350 == WADDR ? 11'h350 : _GEN_847; // @[RAM_ST.scala 31:71]
  assign _GEN_849 = 11'h351 == WADDR ? 11'h351 : _GEN_848; // @[RAM_ST.scala 31:71]
  assign _GEN_850 = 11'h352 == WADDR ? 11'h352 : _GEN_849; // @[RAM_ST.scala 31:71]
  assign _GEN_851 = 11'h353 == WADDR ? 11'h353 : _GEN_850; // @[RAM_ST.scala 31:71]
  assign _GEN_852 = 11'h354 == WADDR ? 11'h354 : _GEN_851; // @[RAM_ST.scala 31:71]
  assign _GEN_853 = 11'h355 == WADDR ? 11'h355 : _GEN_852; // @[RAM_ST.scala 31:71]
  assign _GEN_854 = 11'h356 == WADDR ? 11'h356 : _GEN_853; // @[RAM_ST.scala 31:71]
  assign _GEN_855 = 11'h357 == WADDR ? 11'h357 : _GEN_854; // @[RAM_ST.scala 31:71]
  assign _GEN_856 = 11'h358 == WADDR ? 11'h358 : _GEN_855; // @[RAM_ST.scala 31:71]
  assign _GEN_857 = 11'h359 == WADDR ? 11'h359 : _GEN_856; // @[RAM_ST.scala 31:71]
  assign _GEN_858 = 11'h35a == WADDR ? 11'h35a : _GEN_857; // @[RAM_ST.scala 31:71]
  assign _GEN_859 = 11'h35b == WADDR ? 11'h35b : _GEN_858; // @[RAM_ST.scala 31:71]
  assign _GEN_860 = 11'h35c == WADDR ? 11'h35c : _GEN_859; // @[RAM_ST.scala 31:71]
  assign _GEN_861 = 11'h35d == WADDR ? 11'h35d : _GEN_860; // @[RAM_ST.scala 31:71]
  assign _GEN_862 = 11'h35e == WADDR ? 11'h35e : _GEN_861; // @[RAM_ST.scala 31:71]
  assign _GEN_863 = 11'h35f == WADDR ? 11'h35f : _GEN_862; // @[RAM_ST.scala 31:71]
  assign _GEN_864 = 11'h360 == WADDR ? 11'h360 : _GEN_863; // @[RAM_ST.scala 31:71]
  assign _GEN_865 = 11'h361 == WADDR ? 11'h361 : _GEN_864; // @[RAM_ST.scala 31:71]
  assign _GEN_866 = 11'h362 == WADDR ? 11'h362 : _GEN_865; // @[RAM_ST.scala 31:71]
  assign _GEN_867 = 11'h363 == WADDR ? 11'h363 : _GEN_866; // @[RAM_ST.scala 31:71]
  assign _GEN_868 = 11'h364 == WADDR ? 11'h364 : _GEN_867; // @[RAM_ST.scala 31:71]
  assign _GEN_869 = 11'h365 == WADDR ? 11'h365 : _GEN_868; // @[RAM_ST.scala 31:71]
  assign _GEN_870 = 11'h366 == WADDR ? 11'h366 : _GEN_869; // @[RAM_ST.scala 31:71]
  assign _GEN_871 = 11'h367 == WADDR ? 11'h367 : _GEN_870; // @[RAM_ST.scala 31:71]
  assign _GEN_872 = 11'h368 == WADDR ? 11'h368 : _GEN_871; // @[RAM_ST.scala 31:71]
  assign _GEN_873 = 11'h369 == WADDR ? 11'h369 : _GEN_872; // @[RAM_ST.scala 31:71]
  assign _GEN_874 = 11'h36a == WADDR ? 11'h36a : _GEN_873; // @[RAM_ST.scala 31:71]
  assign _GEN_875 = 11'h36b == WADDR ? 11'h36b : _GEN_874; // @[RAM_ST.scala 31:71]
  assign _GEN_876 = 11'h36c == WADDR ? 11'h36c : _GEN_875; // @[RAM_ST.scala 31:71]
  assign _GEN_877 = 11'h36d == WADDR ? 11'h36d : _GEN_876; // @[RAM_ST.scala 31:71]
  assign _GEN_878 = 11'h36e == WADDR ? 11'h36e : _GEN_877; // @[RAM_ST.scala 31:71]
  assign _GEN_879 = 11'h36f == WADDR ? 11'h36f : _GEN_878; // @[RAM_ST.scala 31:71]
  assign _GEN_880 = 11'h370 == WADDR ? 11'h370 : _GEN_879; // @[RAM_ST.scala 31:71]
  assign _GEN_881 = 11'h371 == WADDR ? 11'h371 : _GEN_880; // @[RAM_ST.scala 31:71]
  assign _GEN_882 = 11'h372 == WADDR ? 11'h372 : _GEN_881; // @[RAM_ST.scala 31:71]
  assign _GEN_883 = 11'h373 == WADDR ? 11'h373 : _GEN_882; // @[RAM_ST.scala 31:71]
  assign _GEN_884 = 11'h374 == WADDR ? 11'h374 : _GEN_883; // @[RAM_ST.scala 31:71]
  assign _GEN_885 = 11'h375 == WADDR ? 11'h375 : _GEN_884; // @[RAM_ST.scala 31:71]
  assign _GEN_886 = 11'h376 == WADDR ? 11'h376 : _GEN_885; // @[RAM_ST.scala 31:71]
  assign _GEN_887 = 11'h377 == WADDR ? 11'h377 : _GEN_886; // @[RAM_ST.scala 31:71]
  assign _GEN_888 = 11'h378 == WADDR ? 11'h378 : _GEN_887; // @[RAM_ST.scala 31:71]
  assign _GEN_889 = 11'h379 == WADDR ? 11'h379 : _GEN_888; // @[RAM_ST.scala 31:71]
  assign _GEN_890 = 11'h37a == WADDR ? 11'h37a : _GEN_889; // @[RAM_ST.scala 31:71]
  assign _GEN_891 = 11'h37b == WADDR ? 11'h37b : _GEN_890; // @[RAM_ST.scala 31:71]
  assign _GEN_892 = 11'h37c == WADDR ? 11'h37c : _GEN_891; // @[RAM_ST.scala 31:71]
  assign _GEN_893 = 11'h37d == WADDR ? 11'h37d : _GEN_892; // @[RAM_ST.scala 31:71]
  assign _GEN_894 = 11'h37e == WADDR ? 11'h37e : _GEN_893; // @[RAM_ST.scala 31:71]
  assign _GEN_895 = 11'h37f == WADDR ? 11'h37f : _GEN_894; // @[RAM_ST.scala 31:71]
  assign _GEN_896 = 11'h380 == WADDR ? 11'h380 : _GEN_895; // @[RAM_ST.scala 31:71]
  assign _GEN_897 = 11'h381 == WADDR ? 11'h381 : _GEN_896; // @[RAM_ST.scala 31:71]
  assign _GEN_898 = 11'h382 == WADDR ? 11'h382 : _GEN_897; // @[RAM_ST.scala 31:71]
  assign _GEN_899 = 11'h383 == WADDR ? 11'h383 : _GEN_898; // @[RAM_ST.scala 31:71]
  assign _GEN_900 = 11'h384 == WADDR ? 11'h384 : _GEN_899; // @[RAM_ST.scala 31:71]
  assign _GEN_901 = 11'h385 == WADDR ? 11'h385 : _GEN_900; // @[RAM_ST.scala 31:71]
  assign _GEN_902 = 11'h386 == WADDR ? 11'h386 : _GEN_901; // @[RAM_ST.scala 31:71]
  assign _GEN_903 = 11'h387 == WADDR ? 11'h387 : _GEN_902; // @[RAM_ST.scala 31:71]
  assign _GEN_904 = 11'h388 == WADDR ? 11'h388 : _GEN_903; // @[RAM_ST.scala 31:71]
  assign _GEN_905 = 11'h389 == WADDR ? 11'h389 : _GEN_904; // @[RAM_ST.scala 31:71]
  assign _GEN_906 = 11'h38a == WADDR ? 11'h38a : _GEN_905; // @[RAM_ST.scala 31:71]
  assign _GEN_907 = 11'h38b == WADDR ? 11'h38b : _GEN_906; // @[RAM_ST.scala 31:71]
  assign _GEN_908 = 11'h38c == WADDR ? 11'h38c : _GEN_907; // @[RAM_ST.scala 31:71]
  assign _GEN_909 = 11'h38d == WADDR ? 11'h38d : _GEN_908; // @[RAM_ST.scala 31:71]
  assign _GEN_910 = 11'h38e == WADDR ? 11'h38e : _GEN_909; // @[RAM_ST.scala 31:71]
  assign _GEN_911 = 11'h38f == WADDR ? 11'h38f : _GEN_910; // @[RAM_ST.scala 31:71]
  assign _GEN_912 = 11'h390 == WADDR ? 11'h390 : _GEN_911; // @[RAM_ST.scala 31:71]
  assign _GEN_913 = 11'h391 == WADDR ? 11'h391 : _GEN_912; // @[RAM_ST.scala 31:71]
  assign _GEN_914 = 11'h392 == WADDR ? 11'h392 : _GEN_913; // @[RAM_ST.scala 31:71]
  assign _GEN_915 = 11'h393 == WADDR ? 11'h393 : _GEN_914; // @[RAM_ST.scala 31:71]
  assign _GEN_916 = 11'h394 == WADDR ? 11'h394 : _GEN_915; // @[RAM_ST.scala 31:71]
  assign _GEN_917 = 11'h395 == WADDR ? 11'h395 : _GEN_916; // @[RAM_ST.scala 31:71]
  assign _GEN_918 = 11'h396 == WADDR ? 11'h396 : _GEN_917; // @[RAM_ST.scala 31:71]
  assign _GEN_919 = 11'h397 == WADDR ? 11'h397 : _GEN_918; // @[RAM_ST.scala 31:71]
  assign _GEN_920 = 11'h398 == WADDR ? 11'h398 : _GEN_919; // @[RAM_ST.scala 31:71]
  assign _GEN_921 = 11'h399 == WADDR ? 11'h399 : _GEN_920; // @[RAM_ST.scala 31:71]
  assign _GEN_922 = 11'h39a == WADDR ? 11'h39a : _GEN_921; // @[RAM_ST.scala 31:71]
  assign _GEN_923 = 11'h39b == WADDR ? 11'h39b : _GEN_922; // @[RAM_ST.scala 31:71]
  assign _GEN_924 = 11'h39c == WADDR ? 11'h39c : _GEN_923; // @[RAM_ST.scala 31:71]
  assign _GEN_925 = 11'h39d == WADDR ? 11'h39d : _GEN_924; // @[RAM_ST.scala 31:71]
  assign _GEN_926 = 11'h39e == WADDR ? 11'h39e : _GEN_925; // @[RAM_ST.scala 31:71]
  assign _GEN_927 = 11'h39f == WADDR ? 11'h39f : _GEN_926; // @[RAM_ST.scala 31:71]
  assign _GEN_928 = 11'h3a0 == WADDR ? 11'h3a0 : _GEN_927; // @[RAM_ST.scala 31:71]
  assign _GEN_929 = 11'h3a1 == WADDR ? 11'h3a1 : _GEN_928; // @[RAM_ST.scala 31:71]
  assign _GEN_930 = 11'h3a2 == WADDR ? 11'h3a2 : _GEN_929; // @[RAM_ST.scala 31:71]
  assign _GEN_931 = 11'h3a3 == WADDR ? 11'h3a3 : _GEN_930; // @[RAM_ST.scala 31:71]
  assign _GEN_932 = 11'h3a4 == WADDR ? 11'h3a4 : _GEN_931; // @[RAM_ST.scala 31:71]
  assign _GEN_933 = 11'h3a5 == WADDR ? 11'h3a5 : _GEN_932; // @[RAM_ST.scala 31:71]
  assign _GEN_934 = 11'h3a6 == WADDR ? 11'h3a6 : _GEN_933; // @[RAM_ST.scala 31:71]
  assign _GEN_935 = 11'h3a7 == WADDR ? 11'h3a7 : _GEN_934; // @[RAM_ST.scala 31:71]
  assign _GEN_936 = 11'h3a8 == WADDR ? 11'h3a8 : _GEN_935; // @[RAM_ST.scala 31:71]
  assign _GEN_937 = 11'h3a9 == WADDR ? 11'h3a9 : _GEN_936; // @[RAM_ST.scala 31:71]
  assign _GEN_938 = 11'h3aa == WADDR ? 11'h3aa : _GEN_937; // @[RAM_ST.scala 31:71]
  assign _GEN_939 = 11'h3ab == WADDR ? 11'h3ab : _GEN_938; // @[RAM_ST.scala 31:71]
  assign _GEN_940 = 11'h3ac == WADDR ? 11'h3ac : _GEN_939; // @[RAM_ST.scala 31:71]
  assign _GEN_941 = 11'h3ad == WADDR ? 11'h3ad : _GEN_940; // @[RAM_ST.scala 31:71]
  assign _GEN_942 = 11'h3ae == WADDR ? 11'h3ae : _GEN_941; // @[RAM_ST.scala 31:71]
  assign _GEN_943 = 11'h3af == WADDR ? 11'h3af : _GEN_942; // @[RAM_ST.scala 31:71]
  assign _GEN_944 = 11'h3b0 == WADDR ? 11'h3b0 : _GEN_943; // @[RAM_ST.scala 31:71]
  assign _GEN_945 = 11'h3b1 == WADDR ? 11'h3b1 : _GEN_944; // @[RAM_ST.scala 31:71]
  assign _GEN_946 = 11'h3b2 == WADDR ? 11'h3b2 : _GEN_945; // @[RAM_ST.scala 31:71]
  assign _GEN_947 = 11'h3b3 == WADDR ? 11'h3b3 : _GEN_946; // @[RAM_ST.scala 31:71]
  assign _GEN_948 = 11'h3b4 == WADDR ? 11'h3b4 : _GEN_947; // @[RAM_ST.scala 31:71]
  assign _GEN_949 = 11'h3b5 == WADDR ? 11'h3b5 : _GEN_948; // @[RAM_ST.scala 31:71]
  assign _GEN_950 = 11'h3b6 == WADDR ? 11'h3b6 : _GEN_949; // @[RAM_ST.scala 31:71]
  assign _GEN_951 = 11'h3b7 == WADDR ? 11'h3b7 : _GEN_950; // @[RAM_ST.scala 31:71]
  assign _GEN_952 = 11'h3b8 == WADDR ? 11'h3b8 : _GEN_951; // @[RAM_ST.scala 31:71]
  assign _GEN_953 = 11'h3b9 == WADDR ? 11'h3b9 : _GEN_952; // @[RAM_ST.scala 31:71]
  assign _GEN_954 = 11'h3ba == WADDR ? 11'h3ba : _GEN_953; // @[RAM_ST.scala 31:71]
  assign _GEN_955 = 11'h3bb == WADDR ? 11'h3bb : _GEN_954; // @[RAM_ST.scala 31:71]
  assign _GEN_956 = 11'h3bc == WADDR ? 11'h3bc : _GEN_955; // @[RAM_ST.scala 31:71]
  assign _GEN_957 = 11'h3bd == WADDR ? 11'h3bd : _GEN_956; // @[RAM_ST.scala 31:71]
  assign _GEN_958 = 11'h3be == WADDR ? 11'h3be : _GEN_957; // @[RAM_ST.scala 31:71]
  assign _GEN_959 = 11'h3bf == WADDR ? 11'h3bf : _GEN_958; // @[RAM_ST.scala 31:71]
  assign _GEN_960 = 11'h3c0 == WADDR ? 11'h3c0 : _GEN_959; // @[RAM_ST.scala 31:71]
  assign _GEN_961 = 11'h3c1 == WADDR ? 11'h3c1 : _GEN_960; // @[RAM_ST.scala 31:71]
  assign _GEN_962 = 11'h3c2 == WADDR ? 11'h3c2 : _GEN_961; // @[RAM_ST.scala 31:71]
  assign _GEN_963 = 11'h3c3 == WADDR ? 11'h3c3 : _GEN_962; // @[RAM_ST.scala 31:71]
  assign _GEN_964 = 11'h3c4 == WADDR ? 11'h3c4 : _GEN_963; // @[RAM_ST.scala 31:71]
  assign _GEN_965 = 11'h3c5 == WADDR ? 11'h3c5 : _GEN_964; // @[RAM_ST.scala 31:71]
  assign _GEN_966 = 11'h3c6 == WADDR ? 11'h3c6 : _GEN_965; // @[RAM_ST.scala 31:71]
  assign _GEN_967 = 11'h3c7 == WADDR ? 11'h3c7 : _GEN_966; // @[RAM_ST.scala 31:71]
  assign _GEN_968 = 11'h3c8 == WADDR ? 11'h3c8 : _GEN_967; // @[RAM_ST.scala 31:71]
  assign _GEN_969 = 11'h3c9 == WADDR ? 11'h3c9 : _GEN_968; // @[RAM_ST.scala 31:71]
  assign _GEN_970 = 11'h3ca == WADDR ? 11'h3ca : _GEN_969; // @[RAM_ST.scala 31:71]
  assign _GEN_971 = 11'h3cb == WADDR ? 11'h3cb : _GEN_970; // @[RAM_ST.scala 31:71]
  assign _GEN_972 = 11'h3cc == WADDR ? 11'h3cc : _GEN_971; // @[RAM_ST.scala 31:71]
  assign _GEN_973 = 11'h3cd == WADDR ? 11'h3cd : _GEN_972; // @[RAM_ST.scala 31:71]
  assign _GEN_974 = 11'h3ce == WADDR ? 11'h3ce : _GEN_973; // @[RAM_ST.scala 31:71]
  assign _GEN_975 = 11'h3cf == WADDR ? 11'h3cf : _GEN_974; // @[RAM_ST.scala 31:71]
  assign _GEN_976 = 11'h3d0 == WADDR ? 11'h3d0 : _GEN_975; // @[RAM_ST.scala 31:71]
  assign _GEN_977 = 11'h3d1 == WADDR ? 11'h3d1 : _GEN_976; // @[RAM_ST.scala 31:71]
  assign _GEN_978 = 11'h3d2 == WADDR ? 11'h3d2 : _GEN_977; // @[RAM_ST.scala 31:71]
  assign _GEN_979 = 11'h3d3 == WADDR ? 11'h3d3 : _GEN_978; // @[RAM_ST.scala 31:71]
  assign _GEN_980 = 11'h3d4 == WADDR ? 11'h3d4 : _GEN_979; // @[RAM_ST.scala 31:71]
  assign _GEN_981 = 11'h3d5 == WADDR ? 11'h3d5 : _GEN_980; // @[RAM_ST.scala 31:71]
  assign _GEN_982 = 11'h3d6 == WADDR ? 11'h3d6 : _GEN_981; // @[RAM_ST.scala 31:71]
  assign _GEN_983 = 11'h3d7 == WADDR ? 11'h3d7 : _GEN_982; // @[RAM_ST.scala 31:71]
  assign _GEN_984 = 11'h3d8 == WADDR ? 11'h3d8 : _GEN_983; // @[RAM_ST.scala 31:71]
  assign _GEN_985 = 11'h3d9 == WADDR ? 11'h3d9 : _GEN_984; // @[RAM_ST.scala 31:71]
  assign _GEN_986 = 11'h3da == WADDR ? 11'h3da : _GEN_985; // @[RAM_ST.scala 31:71]
  assign _GEN_987 = 11'h3db == WADDR ? 11'h3db : _GEN_986; // @[RAM_ST.scala 31:71]
  assign _GEN_988 = 11'h3dc == WADDR ? 11'h3dc : _GEN_987; // @[RAM_ST.scala 31:71]
  assign _GEN_989 = 11'h3dd == WADDR ? 11'h3dd : _GEN_988; // @[RAM_ST.scala 31:71]
  assign _GEN_990 = 11'h3de == WADDR ? 11'h3de : _GEN_989; // @[RAM_ST.scala 31:71]
  assign _GEN_991 = 11'h3df == WADDR ? 11'h3df : _GEN_990; // @[RAM_ST.scala 31:71]
  assign _GEN_992 = 11'h3e0 == WADDR ? 11'h3e0 : _GEN_991; // @[RAM_ST.scala 31:71]
  assign _GEN_993 = 11'h3e1 == WADDR ? 11'h3e1 : _GEN_992; // @[RAM_ST.scala 31:71]
  assign _GEN_994 = 11'h3e2 == WADDR ? 11'h3e2 : _GEN_993; // @[RAM_ST.scala 31:71]
  assign _GEN_995 = 11'h3e3 == WADDR ? 11'h3e3 : _GEN_994; // @[RAM_ST.scala 31:71]
  assign _GEN_996 = 11'h3e4 == WADDR ? 11'h3e4 : _GEN_995; // @[RAM_ST.scala 31:71]
  assign _GEN_997 = 11'h3e5 == WADDR ? 11'h3e5 : _GEN_996; // @[RAM_ST.scala 31:71]
  assign _GEN_998 = 11'h3e6 == WADDR ? 11'h3e6 : _GEN_997; // @[RAM_ST.scala 31:71]
  assign _GEN_999 = 11'h3e7 == WADDR ? 11'h3e7 : _GEN_998; // @[RAM_ST.scala 31:71]
  assign _GEN_1000 = 11'h3e8 == WADDR ? 11'h3e8 : _GEN_999; // @[RAM_ST.scala 31:71]
  assign _GEN_1001 = 11'h3e9 == WADDR ? 11'h3e9 : _GEN_1000; // @[RAM_ST.scala 31:71]
  assign _GEN_1002 = 11'h3ea == WADDR ? 11'h3ea : _GEN_1001; // @[RAM_ST.scala 31:71]
  assign _GEN_1003 = 11'h3eb == WADDR ? 11'h3eb : _GEN_1002; // @[RAM_ST.scala 31:71]
  assign _GEN_1004 = 11'h3ec == WADDR ? 11'h3ec : _GEN_1003; // @[RAM_ST.scala 31:71]
  assign _GEN_1005 = 11'h3ed == WADDR ? 11'h3ed : _GEN_1004; // @[RAM_ST.scala 31:71]
  assign _GEN_1006 = 11'h3ee == WADDR ? 11'h3ee : _GEN_1005; // @[RAM_ST.scala 31:71]
  assign _GEN_1007 = 11'h3ef == WADDR ? 11'h3ef : _GEN_1006; // @[RAM_ST.scala 31:71]
  assign _GEN_1008 = 11'h3f0 == WADDR ? 11'h3f0 : _GEN_1007; // @[RAM_ST.scala 31:71]
  assign _GEN_1009 = 11'h3f1 == WADDR ? 11'h3f1 : _GEN_1008; // @[RAM_ST.scala 31:71]
  assign _GEN_1010 = 11'h3f2 == WADDR ? 11'h3f2 : _GEN_1009; // @[RAM_ST.scala 31:71]
  assign _GEN_1011 = 11'h3f3 == WADDR ? 11'h3f3 : _GEN_1010; // @[RAM_ST.scala 31:71]
  assign _GEN_1012 = 11'h3f4 == WADDR ? 11'h3f4 : _GEN_1011; // @[RAM_ST.scala 31:71]
  assign _GEN_1013 = 11'h3f5 == WADDR ? 11'h3f5 : _GEN_1012; // @[RAM_ST.scala 31:71]
  assign _GEN_1014 = 11'h3f6 == WADDR ? 11'h3f6 : _GEN_1013; // @[RAM_ST.scala 31:71]
  assign _GEN_1015 = 11'h3f7 == WADDR ? 11'h3f7 : _GEN_1014; // @[RAM_ST.scala 31:71]
  assign _GEN_1016 = 11'h3f8 == WADDR ? 11'h3f8 : _GEN_1015; // @[RAM_ST.scala 31:71]
  assign _GEN_1017 = 11'h3f9 == WADDR ? 11'h3f9 : _GEN_1016; // @[RAM_ST.scala 31:71]
  assign _GEN_1018 = 11'h3fa == WADDR ? 11'h3fa : _GEN_1017; // @[RAM_ST.scala 31:71]
  assign _GEN_1019 = 11'h3fb == WADDR ? 11'h3fb : _GEN_1018; // @[RAM_ST.scala 31:71]
  assign _GEN_1020 = 11'h3fc == WADDR ? 11'h3fc : _GEN_1019; // @[RAM_ST.scala 31:71]
  assign _GEN_1021 = 11'h3fd == WADDR ? 11'h3fd : _GEN_1020; // @[RAM_ST.scala 31:71]
  assign _GEN_1022 = 11'h3fe == WADDR ? 11'h3fe : _GEN_1021; // @[RAM_ST.scala 31:71]
  assign _GEN_1023 = 11'h3ff == WADDR ? 11'h3ff : _GEN_1022; // @[RAM_ST.scala 31:71]
  assign _GEN_1024 = 11'h400 == WADDR ? 11'h400 : _GEN_1023; // @[RAM_ST.scala 31:71]
  assign _GEN_1025 = 11'h401 == WADDR ? 11'h401 : _GEN_1024; // @[RAM_ST.scala 31:71]
  assign _GEN_1026 = 11'h402 == WADDR ? 11'h402 : _GEN_1025; // @[RAM_ST.scala 31:71]
  assign _GEN_1027 = 11'h403 == WADDR ? 11'h403 : _GEN_1026; // @[RAM_ST.scala 31:71]
  assign _GEN_1028 = 11'h404 == WADDR ? 11'h404 : _GEN_1027; // @[RAM_ST.scala 31:71]
  assign _GEN_1029 = 11'h405 == WADDR ? 11'h405 : _GEN_1028; // @[RAM_ST.scala 31:71]
  assign _GEN_1030 = 11'h406 == WADDR ? 11'h406 : _GEN_1029; // @[RAM_ST.scala 31:71]
  assign _GEN_1031 = 11'h407 == WADDR ? 11'h407 : _GEN_1030; // @[RAM_ST.scala 31:71]
  assign _GEN_1032 = 11'h408 == WADDR ? 11'h408 : _GEN_1031; // @[RAM_ST.scala 31:71]
  assign _GEN_1033 = 11'h409 == WADDR ? 11'h409 : _GEN_1032; // @[RAM_ST.scala 31:71]
  assign _GEN_1034 = 11'h40a == WADDR ? 11'h40a : _GEN_1033; // @[RAM_ST.scala 31:71]
  assign _GEN_1035 = 11'h40b == WADDR ? 11'h40b : _GEN_1034; // @[RAM_ST.scala 31:71]
  assign _GEN_1036 = 11'h40c == WADDR ? 11'h40c : _GEN_1035; // @[RAM_ST.scala 31:71]
  assign _GEN_1037 = 11'h40d == WADDR ? 11'h40d : _GEN_1036; // @[RAM_ST.scala 31:71]
  assign _GEN_1038 = 11'h40e == WADDR ? 11'h40e : _GEN_1037; // @[RAM_ST.scala 31:71]
  assign _GEN_1039 = 11'h40f == WADDR ? 11'h40f : _GEN_1038; // @[RAM_ST.scala 31:71]
  assign _GEN_1040 = 11'h410 == WADDR ? 11'h410 : _GEN_1039; // @[RAM_ST.scala 31:71]
  assign _GEN_1041 = 11'h411 == WADDR ? 11'h411 : _GEN_1040; // @[RAM_ST.scala 31:71]
  assign _GEN_1042 = 11'h412 == WADDR ? 11'h412 : _GEN_1041; // @[RAM_ST.scala 31:71]
  assign _GEN_1043 = 11'h413 == WADDR ? 11'h413 : _GEN_1042; // @[RAM_ST.scala 31:71]
  assign _GEN_1044 = 11'h414 == WADDR ? 11'h414 : _GEN_1043; // @[RAM_ST.scala 31:71]
  assign _GEN_1045 = 11'h415 == WADDR ? 11'h415 : _GEN_1044; // @[RAM_ST.scala 31:71]
  assign _GEN_1046 = 11'h416 == WADDR ? 11'h416 : _GEN_1045; // @[RAM_ST.scala 31:71]
  assign _GEN_1047 = 11'h417 == WADDR ? 11'h417 : _GEN_1046; // @[RAM_ST.scala 31:71]
  assign _GEN_1048 = 11'h418 == WADDR ? 11'h418 : _GEN_1047; // @[RAM_ST.scala 31:71]
  assign _GEN_1049 = 11'h419 == WADDR ? 11'h419 : _GEN_1048; // @[RAM_ST.scala 31:71]
  assign _GEN_1050 = 11'h41a == WADDR ? 11'h41a : _GEN_1049; // @[RAM_ST.scala 31:71]
  assign _GEN_1051 = 11'h41b == WADDR ? 11'h41b : _GEN_1050; // @[RAM_ST.scala 31:71]
  assign _GEN_1052 = 11'h41c == WADDR ? 11'h41c : _GEN_1051; // @[RAM_ST.scala 31:71]
  assign _GEN_1053 = 11'h41d == WADDR ? 11'h41d : _GEN_1052; // @[RAM_ST.scala 31:71]
  assign _GEN_1054 = 11'h41e == WADDR ? 11'h41e : _GEN_1053; // @[RAM_ST.scala 31:71]
  assign _GEN_1055 = 11'h41f == WADDR ? 11'h41f : _GEN_1054; // @[RAM_ST.scala 31:71]
  assign _GEN_1056 = 11'h420 == WADDR ? 11'h420 : _GEN_1055; // @[RAM_ST.scala 31:71]
  assign _GEN_1057 = 11'h421 == WADDR ? 11'h421 : _GEN_1056; // @[RAM_ST.scala 31:71]
  assign _GEN_1058 = 11'h422 == WADDR ? 11'h422 : _GEN_1057; // @[RAM_ST.scala 31:71]
  assign _GEN_1059 = 11'h423 == WADDR ? 11'h423 : _GEN_1058; // @[RAM_ST.scala 31:71]
  assign _GEN_1060 = 11'h424 == WADDR ? 11'h424 : _GEN_1059; // @[RAM_ST.scala 31:71]
  assign _GEN_1061 = 11'h425 == WADDR ? 11'h425 : _GEN_1060; // @[RAM_ST.scala 31:71]
  assign _GEN_1062 = 11'h426 == WADDR ? 11'h426 : _GEN_1061; // @[RAM_ST.scala 31:71]
  assign _GEN_1063 = 11'h427 == WADDR ? 11'h427 : _GEN_1062; // @[RAM_ST.scala 31:71]
  assign _GEN_1064 = 11'h428 == WADDR ? 11'h428 : _GEN_1063; // @[RAM_ST.scala 31:71]
  assign _GEN_1065 = 11'h429 == WADDR ? 11'h429 : _GEN_1064; // @[RAM_ST.scala 31:71]
  assign _GEN_1066 = 11'h42a == WADDR ? 11'h42a : _GEN_1065; // @[RAM_ST.scala 31:71]
  assign _GEN_1067 = 11'h42b == WADDR ? 11'h42b : _GEN_1066; // @[RAM_ST.scala 31:71]
  assign _GEN_1068 = 11'h42c == WADDR ? 11'h42c : _GEN_1067; // @[RAM_ST.scala 31:71]
  assign _GEN_1069 = 11'h42d == WADDR ? 11'h42d : _GEN_1068; // @[RAM_ST.scala 31:71]
  assign _GEN_1070 = 11'h42e == WADDR ? 11'h42e : _GEN_1069; // @[RAM_ST.scala 31:71]
  assign _GEN_1071 = 11'h42f == WADDR ? 11'h42f : _GEN_1070; // @[RAM_ST.scala 31:71]
  assign _GEN_1072 = 11'h430 == WADDR ? 11'h430 : _GEN_1071; // @[RAM_ST.scala 31:71]
  assign _GEN_1073 = 11'h431 == WADDR ? 11'h431 : _GEN_1072; // @[RAM_ST.scala 31:71]
  assign _GEN_1074 = 11'h432 == WADDR ? 11'h432 : _GEN_1073; // @[RAM_ST.scala 31:71]
  assign _GEN_1075 = 11'h433 == WADDR ? 11'h433 : _GEN_1074; // @[RAM_ST.scala 31:71]
  assign _GEN_1076 = 11'h434 == WADDR ? 11'h434 : _GEN_1075; // @[RAM_ST.scala 31:71]
  assign _GEN_1077 = 11'h435 == WADDR ? 11'h435 : _GEN_1076; // @[RAM_ST.scala 31:71]
  assign _GEN_1078 = 11'h436 == WADDR ? 11'h436 : _GEN_1077; // @[RAM_ST.scala 31:71]
  assign _GEN_1079 = 11'h437 == WADDR ? 11'h437 : _GEN_1078; // @[RAM_ST.scala 31:71]
  assign _GEN_1080 = 11'h438 == WADDR ? 11'h438 : _GEN_1079; // @[RAM_ST.scala 31:71]
  assign _GEN_1081 = 11'h439 == WADDR ? 11'h439 : _GEN_1080; // @[RAM_ST.scala 31:71]
  assign _GEN_1082 = 11'h43a == WADDR ? 11'h43a : _GEN_1081; // @[RAM_ST.scala 31:71]
  assign _GEN_1083 = 11'h43b == WADDR ? 11'h43b : _GEN_1082; // @[RAM_ST.scala 31:71]
  assign _GEN_1084 = 11'h43c == WADDR ? 11'h43c : _GEN_1083; // @[RAM_ST.scala 31:71]
  assign _GEN_1085 = 11'h43d == WADDR ? 11'h43d : _GEN_1084; // @[RAM_ST.scala 31:71]
  assign _GEN_1086 = 11'h43e == WADDR ? 11'h43e : _GEN_1085; // @[RAM_ST.scala 31:71]
  assign _GEN_1087 = 11'h43f == WADDR ? 11'h43f : _GEN_1086; // @[RAM_ST.scala 31:71]
  assign _GEN_1088 = 11'h440 == WADDR ? 11'h440 : _GEN_1087; // @[RAM_ST.scala 31:71]
  assign _GEN_1089 = 11'h441 == WADDR ? 11'h441 : _GEN_1088; // @[RAM_ST.scala 31:71]
  assign _GEN_1090 = 11'h442 == WADDR ? 11'h442 : _GEN_1089; // @[RAM_ST.scala 31:71]
  assign _GEN_1091 = 11'h443 == WADDR ? 11'h443 : _GEN_1090; // @[RAM_ST.scala 31:71]
  assign _GEN_1092 = 11'h444 == WADDR ? 11'h444 : _GEN_1091; // @[RAM_ST.scala 31:71]
  assign _GEN_1093 = 11'h445 == WADDR ? 11'h445 : _GEN_1092; // @[RAM_ST.scala 31:71]
  assign _GEN_1094 = 11'h446 == WADDR ? 11'h446 : _GEN_1093; // @[RAM_ST.scala 31:71]
  assign _GEN_1095 = 11'h447 == WADDR ? 11'h447 : _GEN_1094; // @[RAM_ST.scala 31:71]
  assign _GEN_1096 = 11'h448 == WADDR ? 11'h448 : _GEN_1095; // @[RAM_ST.scala 31:71]
  assign _GEN_1097 = 11'h449 == WADDR ? 11'h449 : _GEN_1096; // @[RAM_ST.scala 31:71]
  assign _GEN_1098 = 11'h44a == WADDR ? 11'h44a : _GEN_1097; // @[RAM_ST.scala 31:71]
  assign _GEN_1099 = 11'h44b == WADDR ? 11'h44b : _GEN_1098; // @[RAM_ST.scala 31:71]
  assign _GEN_1100 = 11'h44c == WADDR ? 11'h44c : _GEN_1099; // @[RAM_ST.scala 31:71]
  assign _GEN_1101 = 11'h44d == WADDR ? 11'h44d : _GEN_1100; // @[RAM_ST.scala 31:71]
  assign _GEN_1102 = 11'h44e == WADDR ? 11'h44e : _GEN_1101; // @[RAM_ST.scala 31:71]
  assign _GEN_1103 = 11'h44f == WADDR ? 11'h44f : _GEN_1102; // @[RAM_ST.scala 31:71]
  assign _GEN_1104 = 11'h450 == WADDR ? 11'h450 : _GEN_1103; // @[RAM_ST.scala 31:71]
  assign _GEN_1105 = 11'h451 == WADDR ? 11'h451 : _GEN_1104; // @[RAM_ST.scala 31:71]
  assign _GEN_1106 = 11'h452 == WADDR ? 11'h452 : _GEN_1105; // @[RAM_ST.scala 31:71]
  assign _GEN_1107 = 11'h453 == WADDR ? 11'h453 : _GEN_1106; // @[RAM_ST.scala 31:71]
  assign _GEN_1108 = 11'h454 == WADDR ? 11'h454 : _GEN_1107; // @[RAM_ST.scala 31:71]
  assign _GEN_1109 = 11'h455 == WADDR ? 11'h455 : _GEN_1108; // @[RAM_ST.scala 31:71]
  assign _GEN_1110 = 11'h456 == WADDR ? 11'h456 : _GEN_1109; // @[RAM_ST.scala 31:71]
  assign _GEN_1111 = 11'h457 == WADDR ? 11'h457 : _GEN_1110; // @[RAM_ST.scala 31:71]
  assign _GEN_1112 = 11'h458 == WADDR ? 11'h458 : _GEN_1111; // @[RAM_ST.scala 31:71]
  assign _GEN_1113 = 11'h459 == WADDR ? 11'h459 : _GEN_1112; // @[RAM_ST.scala 31:71]
  assign _GEN_1114 = 11'h45a == WADDR ? 11'h45a : _GEN_1113; // @[RAM_ST.scala 31:71]
  assign _GEN_1115 = 11'h45b == WADDR ? 11'h45b : _GEN_1114; // @[RAM_ST.scala 31:71]
  assign _GEN_1116 = 11'h45c == WADDR ? 11'h45c : _GEN_1115; // @[RAM_ST.scala 31:71]
  assign _GEN_1117 = 11'h45d == WADDR ? 11'h45d : _GEN_1116; // @[RAM_ST.scala 31:71]
  assign _GEN_1118 = 11'h45e == WADDR ? 11'h45e : _GEN_1117; // @[RAM_ST.scala 31:71]
  assign _GEN_1119 = 11'h45f == WADDR ? 11'h45f : _GEN_1118; // @[RAM_ST.scala 31:71]
  assign _GEN_1120 = 11'h460 == WADDR ? 11'h460 : _GEN_1119; // @[RAM_ST.scala 31:71]
  assign _GEN_1121 = 11'h461 == WADDR ? 11'h461 : _GEN_1120; // @[RAM_ST.scala 31:71]
  assign _GEN_1122 = 11'h462 == WADDR ? 11'h462 : _GEN_1121; // @[RAM_ST.scala 31:71]
  assign _GEN_1123 = 11'h463 == WADDR ? 11'h463 : _GEN_1122; // @[RAM_ST.scala 31:71]
  assign _GEN_1124 = 11'h464 == WADDR ? 11'h464 : _GEN_1123; // @[RAM_ST.scala 31:71]
  assign _GEN_1125 = 11'h465 == WADDR ? 11'h465 : _GEN_1124; // @[RAM_ST.scala 31:71]
  assign _GEN_1126 = 11'h466 == WADDR ? 11'h466 : _GEN_1125; // @[RAM_ST.scala 31:71]
  assign _GEN_1127 = 11'h467 == WADDR ? 11'h467 : _GEN_1126; // @[RAM_ST.scala 31:71]
  assign _GEN_1128 = 11'h468 == WADDR ? 11'h468 : _GEN_1127; // @[RAM_ST.scala 31:71]
  assign _GEN_1129 = 11'h469 == WADDR ? 11'h469 : _GEN_1128; // @[RAM_ST.scala 31:71]
  assign _GEN_1130 = 11'h46a == WADDR ? 11'h46a : _GEN_1129; // @[RAM_ST.scala 31:71]
  assign _GEN_1131 = 11'h46b == WADDR ? 11'h46b : _GEN_1130; // @[RAM_ST.scala 31:71]
  assign _GEN_1132 = 11'h46c == WADDR ? 11'h46c : _GEN_1131; // @[RAM_ST.scala 31:71]
  assign _GEN_1133 = 11'h46d == WADDR ? 11'h46d : _GEN_1132; // @[RAM_ST.scala 31:71]
  assign _GEN_1134 = 11'h46e == WADDR ? 11'h46e : _GEN_1133; // @[RAM_ST.scala 31:71]
  assign _GEN_1135 = 11'h46f == WADDR ? 11'h46f : _GEN_1134; // @[RAM_ST.scala 31:71]
  assign _GEN_1136 = 11'h470 == WADDR ? 11'h470 : _GEN_1135; // @[RAM_ST.scala 31:71]
  assign _GEN_1137 = 11'h471 == WADDR ? 11'h471 : _GEN_1136; // @[RAM_ST.scala 31:71]
  assign _GEN_1138 = 11'h472 == WADDR ? 11'h472 : _GEN_1137; // @[RAM_ST.scala 31:71]
  assign _GEN_1139 = 11'h473 == WADDR ? 11'h473 : _GEN_1138; // @[RAM_ST.scala 31:71]
  assign _GEN_1140 = 11'h474 == WADDR ? 11'h474 : _GEN_1139; // @[RAM_ST.scala 31:71]
  assign _GEN_1141 = 11'h475 == WADDR ? 11'h475 : _GEN_1140; // @[RAM_ST.scala 31:71]
  assign _GEN_1142 = 11'h476 == WADDR ? 11'h476 : _GEN_1141; // @[RAM_ST.scala 31:71]
  assign _GEN_1143 = 11'h477 == WADDR ? 11'h477 : _GEN_1142; // @[RAM_ST.scala 31:71]
  assign _GEN_1144 = 11'h478 == WADDR ? 11'h478 : _GEN_1143; // @[RAM_ST.scala 31:71]
  assign _GEN_1145 = 11'h479 == WADDR ? 11'h479 : _GEN_1144; // @[RAM_ST.scala 31:71]
  assign _GEN_1146 = 11'h47a == WADDR ? 11'h47a : _GEN_1145; // @[RAM_ST.scala 31:71]
  assign _GEN_1147 = 11'h47b == WADDR ? 11'h47b : _GEN_1146; // @[RAM_ST.scala 31:71]
  assign _GEN_1148 = 11'h47c == WADDR ? 11'h47c : _GEN_1147; // @[RAM_ST.scala 31:71]
  assign _GEN_1149 = 11'h47d == WADDR ? 11'h47d : _GEN_1148; // @[RAM_ST.scala 31:71]
  assign _GEN_1150 = 11'h47e == WADDR ? 11'h47e : _GEN_1149; // @[RAM_ST.scala 31:71]
  assign _GEN_1151 = 11'h47f == WADDR ? 11'h47f : _GEN_1150; // @[RAM_ST.scala 31:71]
  assign _GEN_1152 = 11'h480 == WADDR ? 11'h480 : _GEN_1151; // @[RAM_ST.scala 31:71]
  assign _GEN_1153 = 11'h481 == WADDR ? 11'h481 : _GEN_1152; // @[RAM_ST.scala 31:71]
  assign _GEN_1154 = 11'h482 == WADDR ? 11'h482 : _GEN_1153; // @[RAM_ST.scala 31:71]
  assign _GEN_1155 = 11'h483 == WADDR ? 11'h483 : _GEN_1154; // @[RAM_ST.scala 31:71]
  assign _GEN_1156 = 11'h484 == WADDR ? 11'h484 : _GEN_1155; // @[RAM_ST.scala 31:71]
  assign _GEN_1157 = 11'h485 == WADDR ? 11'h485 : _GEN_1156; // @[RAM_ST.scala 31:71]
  assign _GEN_1158 = 11'h486 == WADDR ? 11'h486 : _GEN_1157; // @[RAM_ST.scala 31:71]
  assign _GEN_1159 = 11'h487 == WADDR ? 11'h487 : _GEN_1158; // @[RAM_ST.scala 31:71]
  assign _GEN_1160 = 11'h488 == WADDR ? 11'h488 : _GEN_1159; // @[RAM_ST.scala 31:71]
  assign _GEN_1161 = 11'h489 == WADDR ? 11'h489 : _GEN_1160; // @[RAM_ST.scala 31:71]
  assign _GEN_1162 = 11'h48a == WADDR ? 11'h48a : _GEN_1161; // @[RAM_ST.scala 31:71]
  assign _GEN_1163 = 11'h48b == WADDR ? 11'h48b : _GEN_1162; // @[RAM_ST.scala 31:71]
  assign _GEN_1164 = 11'h48c == WADDR ? 11'h48c : _GEN_1163; // @[RAM_ST.scala 31:71]
  assign _GEN_1165 = 11'h48d == WADDR ? 11'h48d : _GEN_1164; // @[RAM_ST.scala 31:71]
  assign _GEN_1166 = 11'h48e == WADDR ? 11'h48e : _GEN_1165; // @[RAM_ST.scala 31:71]
  assign _GEN_1167 = 11'h48f == WADDR ? 11'h48f : _GEN_1166; // @[RAM_ST.scala 31:71]
  assign _GEN_1168 = 11'h490 == WADDR ? 11'h490 : _GEN_1167; // @[RAM_ST.scala 31:71]
  assign _GEN_1169 = 11'h491 == WADDR ? 11'h491 : _GEN_1168; // @[RAM_ST.scala 31:71]
  assign _GEN_1170 = 11'h492 == WADDR ? 11'h492 : _GEN_1169; // @[RAM_ST.scala 31:71]
  assign _GEN_1171 = 11'h493 == WADDR ? 11'h493 : _GEN_1170; // @[RAM_ST.scala 31:71]
  assign _GEN_1172 = 11'h494 == WADDR ? 11'h494 : _GEN_1171; // @[RAM_ST.scala 31:71]
  assign _GEN_1173 = 11'h495 == WADDR ? 11'h495 : _GEN_1172; // @[RAM_ST.scala 31:71]
  assign _GEN_1174 = 11'h496 == WADDR ? 11'h496 : _GEN_1173; // @[RAM_ST.scala 31:71]
  assign _GEN_1175 = 11'h497 == WADDR ? 11'h497 : _GEN_1174; // @[RAM_ST.scala 31:71]
  assign _GEN_1176 = 11'h498 == WADDR ? 11'h498 : _GEN_1175; // @[RAM_ST.scala 31:71]
  assign _GEN_1177 = 11'h499 == WADDR ? 11'h499 : _GEN_1176; // @[RAM_ST.scala 31:71]
  assign _GEN_1178 = 11'h49a == WADDR ? 11'h49a : _GEN_1177; // @[RAM_ST.scala 31:71]
  assign _GEN_1179 = 11'h49b == WADDR ? 11'h49b : _GEN_1178; // @[RAM_ST.scala 31:71]
  assign _GEN_1180 = 11'h49c == WADDR ? 11'h49c : _GEN_1179; // @[RAM_ST.scala 31:71]
  assign _GEN_1181 = 11'h49d == WADDR ? 11'h49d : _GEN_1180; // @[RAM_ST.scala 31:71]
  assign _GEN_1182 = 11'h49e == WADDR ? 11'h49e : _GEN_1181; // @[RAM_ST.scala 31:71]
  assign _GEN_1183 = 11'h49f == WADDR ? 11'h49f : _GEN_1182; // @[RAM_ST.scala 31:71]
  assign _GEN_1184 = 11'h4a0 == WADDR ? 11'h4a0 : _GEN_1183; // @[RAM_ST.scala 31:71]
  assign _GEN_1185 = 11'h4a1 == WADDR ? 11'h4a1 : _GEN_1184; // @[RAM_ST.scala 31:71]
  assign _GEN_1186 = 11'h4a2 == WADDR ? 11'h4a2 : _GEN_1185; // @[RAM_ST.scala 31:71]
  assign _GEN_1187 = 11'h4a3 == WADDR ? 11'h4a3 : _GEN_1186; // @[RAM_ST.scala 31:71]
  assign _GEN_1188 = 11'h4a4 == WADDR ? 11'h4a4 : _GEN_1187; // @[RAM_ST.scala 31:71]
  assign _GEN_1189 = 11'h4a5 == WADDR ? 11'h4a5 : _GEN_1188; // @[RAM_ST.scala 31:71]
  assign _GEN_1190 = 11'h4a6 == WADDR ? 11'h4a6 : _GEN_1189; // @[RAM_ST.scala 31:71]
  assign _GEN_1191 = 11'h4a7 == WADDR ? 11'h4a7 : _GEN_1190; // @[RAM_ST.scala 31:71]
  assign _GEN_1192 = 11'h4a8 == WADDR ? 11'h4a8 : _GEN_1191; // @[RAM_ST.scala 31:71]
  assign _GEN_1193 = 11'h4a9 == WADDR ? 11'h4a9 : _GEN_1192; // @[RAM_ST.scala 31:71]
  assign _GEN_1194 = 11'h4aa == WADDR ? 11'h4aa : _GEN_1193; // @[RAM_ST.scala 31:71]
  assign _GEN_1195 = 11'h4ab == WADDR ? 11'h4ab : _GEN_1194; // @[RAM_ST.scala 31:71]
  assign _GEN_1196 = 11'h4ac == WADDR ? 11'h4ac : _GEN_1195; // @[RAM_ST.scala 31:71]
  assign _GEN_1197 = 11'h4ad == WADDR ? 11'h4ad : _GEN_1196; // @[RAM_ST.scala 31:71]
  assign _GEN_1198 = 11'h4ae == WADDR ? 11'h4ae : _GEN_1197; // @[RAM_ST.scala 31:71]
  assign _GEN_1199 = 11'h4af == WADDR ? 11'h4af : _GEN_1198; // @[RAM_ST.scala 31:71]
  assign _GEN_1200 = 11'h4b0 == WADDR ? 11'h4b0 : _GEN_1199; // @[RAM_ST.scala 31:71]
  assign _GEN_1201 = 11'h4b1 == WADDR ? 11'h4b1 : _GEN_1200; // @[RAM_ST.scala 31:71]
  assign _GEN_1202 = 11'h4b2 == WADDR ? 11'h4b2 : _GEN_1201; // @[RAM_ST.scala 31:71]
  assign _GEN_1203 = 11'h4b3 == WADDR ? 11'h4b3 : _GEN_1202; // @[RAM_ST.scala 31:71]
  assign _GEN_1204 = 11'h4b4 == WADDR ? 11'h4b4 : _GEN_1203; // @[RAM_ST.scala 31:71]
  assign _GEN_1205 = 11'h4b5 == WADDR ? 11'h4b5 : _GEN_1204; // @[RAM_ST.scala 31:71]
  assign _GEN_1206 = 11'h4b6 == WADDR ? 11'h4b6 : _GEN_1205; // @[RAM_ST.scala 31:71]
  assign _GEN_1207 = 11'h4b7 == WADDR ? 11'h4b7 : _GEN_1206; // @[RAM_ST.scala 31:71]
  assign _GEN_1208 = 11'h4b8 == WADDR ? 11'h4b8 : _GEN_1207; // @[RAM_ST.scala 31:71]
  assign _GEN_1209 = 11'h4b9 == WADDR ? 11'h4b9 : _GEN_1208; // @[RAM_ST.scala 31:71]
  assign _GEN_1210 = 11'h4ba == WADDR ? 11'h4ba : _GEN_1209; // @[RAM_ST.scala 31:71]
  assign _GEN_1211 = 11'h4bb == WADDR ? 11'h4bb : _GEN_1210; // @[RAM_ST.scala 31:71]
  assign _GEN_1212 = 11'h4bc == WADDR ? 11'h4bc : _GEN_1211; // @[RAM_ST.scala 31:71]
  assign _GEN_1213 = 11'h4bd == WADDR ? 11'h4bd : _GEN_1212; // @[RAM_ST.scala 31:71]
  assign _GEN_1214 = 11'h4be == WADDR ? 11'h4be : _GEN_1213; // @[RAM_ST.scala 31:71]
  assign _GEN_1215 = 11'h4bf == WADDR ? 11'h4bf : _GEN_1214; // @[RAM_ST.scala 31:71]
  assign _GEN_1216 = 11'h4c0 == WADDR ? 11'h4c0 : _GEN_1215; // @[RAM_ST.scala 31:71]
  assign _GEN_1217 = 11'h4c1 == WADDR ? 11'h4c1 : _GEN_1216; // @[RAM_ST.scala 31:71]
  assign _GEN_1218 = 11'h4c2 == WADDR ? 11'h4c2 : _GEN_1217; // @[RAM_ST.scala 31:71]
  assign _GEN_1219 = 11'h4c3 == WADDR ? 11'h4c3 : _GEN_1218; // @[RAM_ST.scala 31:71]
  assign _GEN_1220 = 11'h4c4 == WADDR ? 11'h4c4 : _GEN_1219; // @[RAM_ST.scala 31:71]
  assign _GEN_1221 = 11'h4c5 == WADDR ? 11'h4c5 : _GEN_1220; // @[RAM_ST.scala 31:71]
  assign _GEN_1222 = 11'h4c6 == WADDR ? 11'h4c6 : _GEN_1221; // @[RAM_ST.scala 31:71]
  assign _GEN_1223 = 11'h4c7 == WADDR ? 11'h4c7 : _GEN_1222; // @[RAM_ST.scala 31:71]
  assign _GEN_1224 = 11'h4c8 == WADDR ? 11'h4c8 : _GEN_1223; // @[RAM_ST.scala 31:71]
  assign _GEN_1225 = 11'h4c9 == WADDR ? 11'h4c9 : _GEN_1224; // @[RAM_ST.scala 31:71]
  assign _GEN_1226 = 11'h4ca == WADDR ? 11'h4ca : _GEN_1225; // @[RAM_ST.scala 31:71]
  assign _GEN_1227 = 11'h4cb == WADDR ? 11'h4cb : _GEN_1226; // @[RAM_ST.scala 31:71]
  assign _GEN_1228 = 11'h4cc == WADDR ? 11'h4cc : _GEN_1227; // @[RAM_ST.scala 31:71]
  assign _GEN_1229 = 11'h4cd == WADDR ? 11'h4cd : _GEN_1228; // @[RAM_ST.scala 31:71]
  assign _GEN_1230 = 11'h4ce == WADDR ? 11'h4ce : _GEN_1229; // @[RAM_ST.scala 31:71]
  assign _GEN_1231 = 11'h4cf == WADDR ? 11'h4cf : _GEN_1230; // @[RAM_ST.scala 31:71]
  assign _GEN_1232 = 11'h4d0 == WADDR ? 11'h4d0 : _GEN_1231; // @[RAM_ST.scala 31:71]
  assign _GEN_1233 = 11'h4d1 == WADDR ? 11'h4d1 : _GEN_1232; // @[RAM_ST.scala 31:71]
  assign _GEN_1234 = 11'h4d2 == WADDR ? 11'h4d2 : _GEN_1233; // @[RAM_ST.scala 31:71]
  assign _GEN_1235 = 11'h4d3 == WADDR ? 11'h4d3 : _GEN_1234; // @[RAM_ST.scala 31:71]
  assign _GEN_1236 = 11'h4d4 == WADDR ? 11'h4d4 : _GEN_1235; // @[RAM_ST.scala 31:71]
  assign _GEN_1237 = 11'h4d5 == WADDR ? 11'h4d5 : _GEN_1236; // @[RAM_ST.scala 31:71]
  assign _GEN_1238 = 11'h4d6 == WADDR ? 11'h4d6 : _GEN_1237; // @[RAM_ST.scala 31:71]
  assign _GEN_1239 = 11'h4d7 == WADDR ? 11'h4d7 : _GEN_1238; // @[RAM_ST.scala 31:71]
  assign _GEN_1240 = 11'h4d8 == WADDR ? 11'h4d8 : _GEN_1239; // @[RAM_ST.scala 31:71]
  assign _GEN_1241 = 11'h4d9 == WADDR ? 11'h4d9 : _GEN_1240; // @[RAM_ST.scala 31:71]
  assign _GEN_1242 = 11'h4da == WADDR ? 11'h4da : _GEN_1241; // @[RAM_ST.scala 31:71]
  assign _GEN_1243 = 11'h4db == WADDR ? 11'h4db : _GEN_1242; // @[RAM_ST.scala 31:71]
  assign _GEN_1244 = 11'h4dc == WADDR ? 11'h4dc : _GEN_1243; // @[RAM_ST.scala 31:71]
  assign _GEN_1245 = 11'h4dd == WADDR ? 11'h4dd : _GEN_1244; // @[RAM_ST.scala 31:71]
  assign _GEN_1246 = 11'h4de == WADDR ? 11'h4de : _GEN_1245; // @[RAM_ST.scala 31:71]
  assign _GEN_1247 = 11'h4df == WADDR ? 11'h4df : _GEN_1246; // @[RAM_ST.scala 31:71]
  assign _GEN_1248 = 11'h4e0 == WADDR ? 11'h4e0 : _GEN_1247; // @[RAM_ST.scala 31:71]
  assign _GEN_1249 = 11'h4e1 == WADDR ? 11'h4e1 : _GEN_1248; // @[RAM_ST.scala 31:71]
  assign _GEN_1250 = 11'h4e2 == WADDR ? 11'h4e2 : _GEN_1249; // @[RAM_ST.scala 31:71]
  assign _GEN_1251 = 11'h4e3 == WADDR ? 11'h4e3 : _GEN_1250; // @[RAM_ST.scala 31:71]
  assign _GEN_1252 = 11'h4e4 == WADDR ? 11'h4e4 : _GEN_1251; // @[RAM_ST.scala 31:71]
  assign _GEN_1253 = 11'h4e5 == WADDR ? 11'h4e5 : _GEN_1252; // @[RAM_ST.scala 31:71]
  assign _GEN_1254 = 11'h4e6 == WADDR ? 11'h4e6 : _GEN_1253; // @[RAM_ST.scala 31:71]
  assign _GEN_1255 = 11'h4e7 == WADDR ? 11'h4e7 : _GEN_1254; // @[RAM_ST.scala 31:71]
  assign _GEN_1256 = 11'h4e8 == WADDR ? 11'h4e8 : _GEN_1255; // @[RAM_ST.scala 31:71]
  assign _GEN_1257 = 11'h4e9 == WADDR ? 11'h4e9 : _GEN_1256; // @[RAM_ST.scala 31:71]
  assign _GEN_1258 = 11'h4ea == WADDR ? 11'h4ea : _GEN_1257; // @[RAM_ST.scala 31:71]
  assign _GEN_1259 = 11'h4eb == WADDR ? 11'h4eb : _GEN_1258; // @[RAM_ST.scala 31:71]
  assign _GEN_1260 = 11'h4ec == WADDR ? 11'h4ec : _GEN_1259; // @[RAM_ST.scala 31:71]
  assign _GEN_1261 = 11'h4ed == WADDR ? 11'h4ed : _GEN_1260; // @[RAM_ST.scala 31:71]
  assign _GEN_1262 = 11'h4ee == WADDR ? 11'h4ee : _GEN_1261; // @[RAM_ST.scala 31:71]
  assign _GEN_1263 = 11'h4ef == WADDR ? 11'h4ef : _GEN_1262; // @[RAM_ST.scala 31:71]
  assign _GEN_1264 = 11'h4f0 == WADDR ? 11'h4f0 : _GEN_1263; // @[RAM_ST.scala 31:71]
  assign _GEN_1265 = 11'h4f1 == WADDR ? 11'h4f1 : _GEN_1264; // @[RAM_ST.scala 31:71]
  assign _GEN_1266 = 11'h4f2 == WADDR ? 11'h4f2 : _GEN_1265; // @[RAM_ST.scala 31:71]
  assign _GEN_1267 = 11'h4f3 == WADDR ? 11'h4f3 : _GEN_1266; // @[RAM_ST.scala 31:71]
  assign _GEN_1268 = 11'h4f4 == WADDR ? 11'h4f4 : _GEN_1267; // @[RAM_ST.scala 31:71]
  assign _GEN_1269 = 11'h4f5 == WADDR ? 11'h4f5 : _GEN_1268; // @[RAM_ST.scala 31:71]
  assign _GEN_1270 = 11'h4f6 == WADDR ? 11'h4f6 : _GEN_1269; // @[RAM_ST.scala 31:71]
  assign _GEN_1271 = 11'h4f7 == WADDR ? 11'h4f7 : _GEN_1270; // @[RAM_ST.scala 31:71]
  assign _GEN_1272 = 11'h4f8 == WADDR ? 11'h4f8 : _GEN_1271; // @[RAM_ST.scala 31:71]
  assign _GEN_1273 = 11'h4f9 == WADDR ? 11'h4f9 : _GEN_1272; // @[RAM_ST.scala 31:71]
  assign _GEN_1274 = 11'h4fa == WADDR ? 11'h4fa : _GEN_1273; // @[RAM_ST.scala 31:71]
  assign _GEN_1275 = 11'h4fb == WADDR ? 11'h4fb : _GEN_1274; // @[RAM_ST.scala 31:71]
  assign _GEN_1276 = 11'h4fc == WADDR ? 11'h4fc : _GEN_1275; // @[RAM_ST.scala 31:71]
  assign _GEN_1277 = 11'h4fd == WADDR ? 11'h4fd : _GEN_1276; // @[RAM_ST.scala 31:71]
  assign _GEN_1278 = 11'h4fe == WADDR ? 11'h4fe : _GEN_1277; // @[RAM_ST.scala 31:71]
  assign _GEN_1279 = 11'h4ff == WADDR ? 11'h4ff : _GEN_1278; // @[RAM_ST.scala 31:71]
  assign _GEN_1280 = 11'h500 == WADDR ? 11'h500 : _GEN_1279; // @[RAM_ST.scala 31:71]
  assign _GEN_1281 = 11'h501 == WADDR ? 11'h501 : _GEN_1280; // @[RAM_ST.scala 31:71]
  assign _GEN_1282 = 11'h502 == WADDR ? 11'h502 : _GEN_1281; // @[RAM_ST.scala 31:71]
  assign _GEN_1283 = 11'h503 == WADDR ? 11'h503 : _GEN_1282; // @[RAM_ST.scala 31:71]
  assign _GEN_1284 = 11'h504 == WADDR ? 11'h504 : _GEN_1283; // @[RAM_ST.scala 31:71]
  assign _GEN_1285 = 11'h505 == WADDR ? 11'h505 : _GEN_1284; // @[RAM_ST.scala 31:71]
  assign _GEN_1286 = 11'h506 == WADDR ? 11'h506 : _GEN_1285; // @[RAM_ST.scala 31:71]
  assign _GEN_1287 = 11'h507 == WADDR ? 11'h507 : _GEN_1286; // @[RAM_ST.scala 31:71]
  assign _GEN_1288 = 11'h508 == WADDR ? 11'h508 : _GEN_1287; // @[RAM_ST.scala 31:71]
  assign _GEN_1289 = 11'h509 == WADDR ? 11'h509 : _GEN_1288; // @[RAM_ST.scala 31:71]
  assign _GEN_1290 = 11'h50a == WADDR ? 11'h50a : _GEN_1289; // @[RAM_ST.scala 31:71]
  assign _GEN_1291 = 11'h50b == WADDR ? 11'h50b : _GEN_1290; // @[RAM_ST.scala 31:71]
  assign _GEN_1292 = 11'h50c == WADDR ? 11'h50c : _GEN_1291; // @[RAM_ST.scala 31:71]
  assign _GEN_1293 = 11'h50d == WADDR ? 11'h50d : _GEN_1292; // @[RAM_ST.scala 31:71]
  assign _GEN_1294 = 11'h50e == WADDR ? 11'h50e : _GEN_1293; // @[RAM_ST.scala 31:71]
  assign _GEN_1295 = 11'h50f == WADDR ? 11'h50f : _GEN_1294; // @[RAM_ST.scala 31:71]
  assign _GEN_1296 = 11'h510 == WADDR ? 11'h510 : _GEN_1295; // @[RAM_ST.scala 31:71]
  assign _GEN_1297 = 11'h511 == WADDR ? 11'h511 : _GEN_1296; // @[RAM_ST.scala 31:71]
  assign _GEN_1298 = 11'h512 == WADDR ? 11'h512 : _GEN_1297; // @[RAM_ST.scala 31:71]
  assign _GEN_1299 = 11'h513 == WADDR ? 11'h513 : _GEN_1298; // @[RAM_ST.scala 31:71]
  assign _GEN_1300 = 11'h514 == WADDR ? 11'h514 : _GEN_1299; // @[RAM_ST.scala 31:71]
  assign _GEN_1301 = 11'h515 == WADDR ? 11'h515 : _GEN_1300; // @[RAM_ST.scala 31:71]
  assign _GEN_1302 = 11'h516 == WADDR ? 11'h516 : _GEN_1301; // @[RAM_ST.scala 31:71]
  assign _GEN_1303 = 11'h517 == WADDR ? 11'h517 : _GEN_1302; // @[RAM_ST.scala 31:71]
  assign _GEN_1304 = 11'h518 == WADDR ? 11'h518 : _GEN_1303; // @[RAM_ST.scala 31:71]
  assign _GEN_1305 = 11'h519 == WADDR ? 11'h519 : _GEN_1304; // @[RAM_ST.scala 31:71]
  assign _GEN_1306 = 11'h51a == WADDR ? 11'h51a : _GEN_1305; // @[RAM_ST.scala 31:71]
  assign _GEN_1307 = 11'h51b == WADDR ? 11'h51b : _GEN_1306; // @[RAM_ST.scala 31:71]
  assign _GEN_1308 = 11'h51c == WADDR ? 11'h51c : _GEN_1307; // @[RAM_ST.scala 31:71]
  assign _GEN_1309 = 11'h51d == WADDR ? 11'h51d : _GEN_1308; // @[RAM_ST.scala 31:71]
  assign _GEN_1310 = 11'h51e == WADDR ? 11'h51e : _GEN_1309; // @[RAM_ST.scala 31:71]
  assign _GEN_1311 = 11'h51f == WADDR ? 11'h51f : _GEN_1310; // @[RAM_ST.scala 31:71]
  assign _GEN_1312 = 11'h520 == WADDR ? 11'h520 : _GEN_1311; // @[RAM_ST.scala 31:71]
  assign _GEN_1313 = 11'h521 == WADDR ? 11'h521 : _GEN_1312; // @[RAM_ST.scala 31:71]
  assign _GEN_1314 = 11'h522 == WADDR ? 11'h522 : _GEN_1313; // @[RAM_ST.scala 31:71]
  assign _GEN_1315 = 11'h523 == WADDR ? 11'h523 : _GEN_1314; // @[RAM_ST.scala 31:71]
  assign _GEN_1316 = 11'h524 == WADDR ? 11'h524 : _GEN_1315; // @[RAM_ST.scala 31:71]
  assign _GEN_1317 = 11'h525 == WADDR ? 11'h525 : _GEN_1316; // @[RAM_ST.scala 31:71]
  assign _GEN_1318 = 11'h526 == WADDR ? 11'h526 : _GEN_1317; // @[RAM_ST.scala 31:71]
  assign _GEN_1319 = 11'h527 == WADDR ? 11'h527 : _GEN_1318; // @[RAM_ST.scala 31:71]
  assign _GEN_1320 = 11'h528 == WADDR ? 11'h528 : _GEN_1319; // @[RAM_ST.scala 31:71]
  assign _GEN_1321 = 11'h529 == WADDR ? 11'h529 : _GEN_1320; // @[RAM_ST.scala 31:71]
  assign _GEN_1322 = 11'h52a == WADDR ? 11'h52a : _GEN_1321; // @[RAM_ST.scala 31:71]
  assign _GEN_1323 = 11'h52b == WADDR ? 11'h52b : _GEN_1322; // @[RAM_ST.scala 31:71]
  assign _GEN_1324 = 11'h52c == WADDR ? 11'h52c : _GEN_1323; // @[RAM_ST.scala 31:71]
  assign _GEN_1325 = 11'h52d == WADDR ? 11'h52d : _GEN_1324; // @[RAM_ST.scala 31:71]
  assign _GEN_1326 = 11'h52e == WADDR ? 11'h52e : _GEN_1325; // @[RAM_ST.scala 31:71]
  assign _GEN_1327 = 11'h52f == WADDR ? 11'h52f : _GEN_1326; // @[RAM_ST.scala 31:71]
  assign _GEN_1328 = 11'h530 == WADDR ? 11'h530 : _GEN_1327; // @[RAM_ST.scala 31:71]
  assign _GEN_1329 = 11'h531 == WADDR ? 11'h531 : _GEN_1328; // @[RAM_ST.scala 31:71]
  assign _GEN_1330 = 11'h532 == WADDR ? 11'h532 : _GEN_1329; // @[RAM_ST.scala 31:71]
  assign _GEN_1331 = 11'h533 == WADDR ? 11'h533 : _GEN_1330; // @[RAM_ST.scala 31:71]
  assign _GEN_1332 = 11'h534 == WADDR ? 11'h534 : _GEN_1331; // @[RAM_ST.scala 31:71]
  assign _GEN_1333 = 11'h535 == WADDR ? 11'h535 : _GEN_1332; // @[RAM_ST.scala 31:71]
  assign _GEN_1334 = 11'h536 == WADDR ? 11'h536 : _GEN_1333; // @[RAM_ST.scala 31:71]
  assign _GEN_1335 = 11'h537 == WADDR ? 11'h537 : _GEN_1334; // @[RAM_ST.scala 31:71]
  assign _GEN_1336 = 11'h538 == WADDR ? 11'h538 : _GEN_1335; // @[RAM_ST.scala 31:71]
  assign _GEN_1337 = 11'h539 == WADDR ? 11'h539 : _GEN_1336; // @[RAM_ST.scala 31:71]
  assign _GEN_1338 = 11'h53a == WADDR ? 11'h53a : _GEN_1337; // @[RAM_ST.scala 31:71]
  assign _GEN_1339 = 11'h53b == WADDR ? 11'h53b : _GEN_1338; // @[RAM_ST.scala 31:71]
  assign _GEN_1340 = 11'h53c == WADDR ? 11'h53c : _GEN_1339; // @[RAM_ST.scala 31:71]
  assign _GEN_1341 = 11'h53d == WADDR ? 11'h53d : _GEN_1340; // @[RAM_ST.scala 31:71]
  assign _GEN_1342 = 11'h53e == WADDR ? 11'h53e : _GEN_1341; // @[RAM_ST.scala 31:71]
  assign _GEN_1343 = 11'h53f == WADDR ? 11'h53f : _GEN_1342; // @[RAM_ST.scala 31:71]
  assign _GEN_1344 = 11'h540 == WADDR ? 11'h540 : _GEN_1343; // @[RAM_ST.scala 31:71]
  assign _GEN_1345 = 11'h541 == WADDR ? 11'h541 : _GEN_1344; // @[RAM_ST.scala 31:71]
  assign _GEN_1346 = 11'h542 == WADDR ? 11'h542 : _GEN_1345; // @[RAM_ST.scala 31:71]
  assign _GEN_1347 = 11'h543 == WADDR ? 11'h543 : _GEN_1346; // @[RAM_ST.scala 31:71]
  assign _GEN_1348 = 11'h544 == WADDR ? 11'h544 : _GEN_1347; // @[RAM_ST.scala 31:71]
  assign _GEN_1349 = 11'h545 == WADDR ? 11'h545 : _GEN_1348; // @[RAM_ST.scala 31:71]
  assign _GEN_1350 = 11'h546 == WADDR ? 11'h546 : _GEN_1349; // @[RAM_ST.scala 31:71]
  assign _GEN_1351 = 11'h547 == WADDR ? 11'h547 : _GEN_1350; // @[RAM_ST.scala 31:71]
  assign _GEN_1352 = 11'h548 == WADDR ? 11'h548 : _GEN_1351; // @[RAM_ST.scala 31:71]
  assign _GEN_1353 = 11'h549 == WADDR ? 11'h549 : _GEN_1352; // @[RAM_ST.scala 31:71]
  assign _GEN_1354 = 11'h54a == WADDR ? 11'h54a : _GEN_1353; // @[RAM_ST.scala 31:71]
  assign _GEN_1355 = 11'h54b == WADDR ? 11'h54b : _GEN_1354; // @[RAM_ST.scala 31:71]
  assign _GEN_1356 = 11'h54c == WADDR ? 11'h54c : _GEN_1355; // @[RAM_ST.scala 31:71]
  assign _GEN_1357 = 11'h54d == WADDR ? 11'h54d : _GEN_1356; // @[RAM_ST.scala 31:71]
  assign _GEN_1358 = 11'h54e == WADDR ? 11'h54e : _GEN_1357; // @[RAM_ST.scala 31:71]
  assign _GEN_1359 = 11'h54f == WADDR ? 11'h54f : _GEN_1358; // @[RAM_ST.scala 31:71]
  assign _GEN_1360 = 11'h550 == WADDR ? 11'h550 : _GEN_1359; // @[RAM_ST.scala 31:71]
  assign _GEN_1361 = 11'h551 == WADDR ? 11'h551 : _GEN_1360; // @[RAM_ST.scala 31:71]
  assign _GEN_1362 = 11'h552 == WADDR ? 11'h552 : _GEN_1361; // @[RAM_ST.scala 31:71]
  assign _GEN_1363 = 11'h553 == WADDR ? 11'h553 : _GEN_1362; // @[RAM_ST.scala 31:71]
  assign _GEN_1364 = 11'h554 == WADDR ? 11'h554 : _GEN_1363; // @[RAM_ST.scala 31:71]
  assign _GEN_1365 = 11'h555 == WADDR ? 11'h555 : _GEN_1364; // @[RAM_ST.scala 31:71]
  assign _GEN_1366 = 11'h556 == WADDR ? 11'h556 : _GEN_1365; // @[RAM_ST.scala 31:71]
  assign _GEN_1367 = 11'h557 == WADDR ? 11'h557 : _GEN_1366; // @[RAM_ST.scala 31:71]
  assign _GEN_1368 = 11'h558 == WADDR ? 11'h558 : _GEN_1367; // @[RAM_ST.scala 31:71]
  assign _GEN_1369 = 11'h559 == WADDR ? 11'h559 : _GEN_1368; // @[RAM_ST.scala 31:71]
  assign _GEN_1370 = 11'h55a == WADDR ? 11'h55a : _GEN_1369; // @[RAM_ST.scala 31:71]
  assign _GEN_1371 = 11'h55b == WADDR ? 11'h55b : _GEN_1370; // @[RAM_ST.scala 31:71]
  assign _GEN_1372 = 11'h55c == WADDR ? 11'h55c : _GEN_1371; // @[RAM_ST.scala 31:71]
  assign _GEN_1373 = 11'h55d == WADDR ? 11'h55d : _GEN_1372; // @[RAM_ST.scala 31:71]
  assign _GEN_1374 = 11'h55e == WADDR ? 11'h55e : _GEN_1373; // @[RAM_ST.scala 31:71]
  assign _GEN_1375 = 11'h55f == WADDR ? 11'h55f : _GEN_1374; // @[RAM_ST.scala 31:71]
  assign _GEN_1376 = 11'h560 == WADDR ? 11'h560 : _GEN_1375; // @[RAM_ST.scala 31:71]
  assign _GEN_1377 = 11'h561 == WADDR ? 11'h561 : _GEN_1376; // @[RAM_ST.scala 31:71]
  assign _GEN_1378 = 11'h562 == WADDR ? 11'h562 : _GEN_1377; // @[RAM_ST.scala 31:71]
  assign _GEN_1379 = 11'h563 == WADDR ? 11'h563 : _GEN_1378; // @[RAM_ST.scala 31:71]
  assign _GEN_1380 = 11'h564 == WADDR ? 11'h564 : _GEN_1379; // @[RAM_ST.scala 31:71]
  assign _GEN_1381 = 11'h565 == WADDR ? 11'h565 : _GEN_1380; // @[RAM_ST.scala 31:71]
  assign _GEN_1382 = 11'h566 == WADDR ? 11'h566 : _GEN_1381; // @[RAM_ST.scala 31:71]
  assign _GEN_1383 = 11'h567 == WADDR ? 11'h567 : _GEN_1382; // @[RAM_ST.scala 31:71]
  assign _GEN_1384 = 11'h568 == WADDR ? 11'h568 : _GEN_1383; // @[RAM_ST.scala 31:71]
  assign _GEN_1385 = 11'h569 == WADDR ? 11'h569 : _GEN_1384; // @[RAM_ST.scala 31:71]
  assign _GEN_1386 = 11'h56a == WADDR ? 11'h56a : _GEN_1385; // @[RAM_ST.scala 31:71]
  assign _GEN_1387 = 11'h56b == WADDR ? 11'h56b : _GEN_1386; // @[RAM_ST.scala 31:71]
  assign _GEN_1388 = 11'h56c == WADDR ? 11'h56c : _GEN_1387; // @[RAM_ST.scala 31:71]
  assign _GEN_1389 = 11'h56d == WADDR ? 11'h56d : _GEN_1388; // @[RAM_ST.scala 31:71]
  assign _GEN_1390 = 11'h56e == WADDR ? 11'h56e : _GEN_1389; // @[RAM_ST.scala 31:71]
  assign _GEN_1391 = 11'h56f == WADDR ? 11'h56f : _GEN_1390; // @[RAM_ST.scala 31:71]
  assign _GEN_1392 = 11'h570 == WADDR ? 11'h570 : _GEN_1391; // @[RAM_ST.scala 31:71]
  assign _GEN_1393 = 11'h571 == WADDR ? 11'h571 : _GEN_1392; // @[RAM_ST.scala 31:71]
  assign _GEN_1394 = 11'h572 == WADDR ? 11'h572 : _GEN_1393; // @[RAM_ST.scala 31:71]
  assign _GEN_1395 = 11'h573 == WADDR ? 11'h573 : _GEN_1394; // @[RAM_ST.scala 31:71]
  assign _GEN_1396 = 11'h574 == WADDR ? 11'h574 : _GEN_1395; // @[RAM_ST.scala 31:71]
  assign _GEN_1397 = 11'h575 == WADDR ? 11'h575 : _GEN_1396; // @[RAM_ST.scala 31:71]
  assign _GEN_1398 = 11'h576 == WADDR ? 11'h576 : _GEN_1397; // @[RAM_ST.scala 31:71]
  assign _GEN_1399 = 11'h577 == WADDR ? 11'h577 : _GEN_1398; // @[RAM_ST.scala 31:71]
  assign _GEN_1400 = 11'h578 == WADDR ? 11'h578 : _GEN_1399; // @[RAM_ST.scala 31:71]
  assign _GEN_1401 = 11'h579 == WADDR ? 11'h579 : _GEN_1400; // @[RAM_ST.scala 31:71]
  assign _GEN_1402 = 11'h57a == WADDR ? 11'h57a : _GEN_1401; // @[RAM_ST.scala 31:71]
  assign _GEN_1403 = 11'h57b == WADDR ? 11'h57b : _GEN_1402; // @[RAM_ST.scala 31:71]
  assign _GEN_1404 = 11'h57c == WADDR ? 11'h57c : _GEN_1403; // @[RAM_ST.scala 31:71]
  assign _GEN_1405 = 11'h57d == WADDR ? 11'h57d : _GEN_1404; // @[RAM_ST.scala 31:71]
  assign _GEN_1406 = 11'h57e == WADDR ? 11'h57e : _GEN_1405; // @[RAM_ST.scala 31:71]
  assign _GEN_1407 = 11'h57f == WADDR ? 11'h57f : _GEN_1406; // @[RAM_ST.scala 31:71]
  assign _GEN_1408 = 11'h580 == WADDR ? 11'h580 : _GEN_1407; // @[RAM_ST.scala 31:71]
  assign _GEN_1409 = 11'h581 == WADDR ? 11'h581 : _GEN_1408; // @[RAM_ST.scala 31:71]
  assign _GEN_1410 = 11'h582 == WADDR ? 11'h582 : _GEN_1409; // @[RAM_ST.scala 31:71]
  assign _GEN_1411 = 11'h583 == WADDR ? 11'h583 : _GEN_1410; // @[RAM_ST.scala 31:71]
  assign _GEN_1412 = 11'h584 == WADDR ? 11'h584 : _GEN_1411; // @[RAM_ST.scala 31:71]
  assign _GEN_1413 = 11'h585 == WADDR ? 11'h585 : _GEN_1412; // @[RAM_ST.scala 31:71]
  assign _GEN_1414 = 11'h586 == WADDR ? 11'h586 : _GEN_1413; // @[RAM_ST.scala 31:71]
  assign _GEN_1415 = 11'h587 == WADDR ? 11'h587 : _GEN_1414; // @[RAM_ST.scala 31:71]
  assign _GEN_1416 = 11'h588 == WADDR ? 11'h588 : _GEN_1415; // @[RAM_ST.scala 31:71]
  assign _GEN_1417 = 11'h589 == WADDR ? 11'h589 : _GEN_1416; // @[RAM_ST.scala 31:71]
  assign _GEN_1418 = 11'h58a == WADDR ? 11'h58a : _GEN_1417; // @[RAM_ST.scala 31:71]
  assign _GEN_1419 = 11'h58b == WADDR ? 11'h58b : _GEN_1418; // @[RAM_ST.scala 31:71]
  assign _GEN_1420 = 11'h58c == WADDR ? 11'h58c : _GEN_1419; // @[RAM_ST.scala 31:71]
  assign _GEN_1421 = 11'h58d == WADDR ? 11'h58d : _GEN_1420; // @[RAM_ST.scala 31:71]
  assign _GEN_1422 = 11'h58e == WADDR ? 11'h58e : _GEN_1421; // @[RAM_ST.scala 31:71]
  assign _GEN_1423 = 11'h58f == WADDR ? 11'h58f : _GEN_1422; // @[RAM_ST.scala 31:71]
  assign _GEN_1424 = 11'h590 == WADDR ? 11'h590 : _GEN_1423; // @[RAM_ST.scala 31:71]
  assign _GEN_1425 = 11'h591 == WADDR ? 11'h591 : _GEN_1424; // @[RAM_ST.scala 31:71]
  assign _GEN_1426 = 11'h592 == WADDR ? 11'h592 : _GEN_1425; // @[RAM_ST.scala 31:71]
  assign _GEN_1427 = 11'h593 == WADDR ? 11'h593 : _GEN_1426; // @[RAM_ST.scala 31:71]
  assign _GEN_1428 = 11'h594 == WADDR ? 11'h594 : _GEN_1427; // @[RAM_ST.scala 31:71]
  assign _GEN_1429 = 11'h595 == WADDR ? 11'h595 : _GEN_1428; // @[RAM_ST.scala 31:71]
  assign _GEN_1430 = 11'h596 == WADDR ? 11'h596 : _GEN_1429; // @[RAM_ST.scala 31:71]
  assign _GEN_1431 = 11'h597 == WADDR ? 11'h597 : _GEN_1430; // @[RAM_ST.scala 31:71]
  assign _GEN_1432 = 11'h598 == WADDR ? 11'h598 : _GEN_1431; // @[RAM_ST.scala 31:71]
  assign _GEN_1433 = 11'h599 == WADDR ? 11'h599 : _GEN_1432; // @[RAM_ST.scala 31:71]
  assign _GEN_1434 = 11'h59a == WADDR ? 11'h59a : _GEN_1433; // @[RAM_ST.scala 31:71]
  assign _GEN_1435 = 11'h59b == WADDR ? 11'h59b : _GEN_1434; // @[RAM_ST.scala 31:71]
  assign _GEN_1436 = 11'h59c == WADDR ? 11'h59c : _GEN_1435; // @[RAM_ST.scala 31:71]
  assign _GEN_1437 = 11'h59d == WADDR ? 11'h59d : _GEN_1436; // @[RAM_ST.scala 31:71]
  assign _GEN_1438 = 11'h59e == WADDR ? 11'h59e : _GEN_1437; // @[RAM_ST.scala 31:71]
  assign _GEN_1439 = 11'h59f == WADDR ? 11'h59f : _GEN_1438; // @[RAM_ST.scala 31:71]
  assign _GEN_1440 = 11'h5a0 == WADDR ? 11'h5a0 : _GEN_1439; // @[RAM_ST.scala 31:71]
  assign _GEN_1441 = 11'h5a1 == WADDR ? 11'h5a1 : _GEN_1440; // @[RAM_ST.scala 31:71]
  assign _GEN_1442 = 11'h5a2 == WADDR ? 11'h5a2 : _GEN_1441; // @[RAM_ST.scala 31:71]
  assign _GEN_1443 = 11'h5a3 == WADDR ? 11'h5a3 : _GEN_1442; // @[RAM_ST.scala 31:71]
  assign _GEN_1444 = 11'h5a4 == WADDR ? 11'h5a4 : _GEN_1443; // @[RAM_ST.scala 31:71]
  assign _GEN_1445 = 11'h5a5 == WADDR ? 11'h5a5 : _GEN_1444; // @[RAM_ST.scala 31:71]
  assign _GEN_1446 = 11'h5a6 == WADDR ? 11'h5a6 : _GEN_1445; // @[RAM_ST.scala 31:71]
  assign _GEN_1447 = 11'h5a7 == WADDR ? 11'h5a7 : _GEN_1446; // @[RAM_ST.scala 31:71]
  assign _GEN_1448 = 11'h5a8 == WADDR ? 11'h5a8 : _GEN_1447; // @[RAM_ST.scala 31:71]
  assign _GEN_1449 = 11'h5a9 == WADDR ? 11'h5a9 : _GEN_1448; // @[RAM_ST.scala 31:71]
  assign _GEN_1450 = 11'h5aa == WADDR ? 11'h5aa : _GEN_1449; // @[RAM_ST.scala 31:71]
  assign _GEN_1451 = 11'h5ab == WADDR ? 11'h5ab : _GEN_1450; // @[RAM_ST.scala 31:71]
  assign _GEN_1452 = 11'h5ac == WADDR ? 11'h5ac : _GEN_1451; // @[RAM_ST.scala 31:71]
  assign _GEN_1453 = 11'h5ad == WADDR ? 11'h5ad : _GEN_1452; // @[RAM_ST.scala 31:71]
  assign _GEN_1454 = 11'h5ae == WADDR ? 11'h5ae : _GEN_1453; // @[RAM_ST.scala 31:71]
  assign _GEN_1455 = 11'h5af == WADDR ? 11'h5af : _GEN_1454; // @[RAM_ST.scala 31:71]
  assign _GEN_1456 = 11'h5b0 == WADDR ? 11'h5b0 : _GEN_1455; // @[RAM_ST.scala 31:71]
  assign _GEN_1457 = 11'h5b1 == WADDR ? 11'h5b1 : _GEN_1456; // @[RAM_ST.scala 31:71]
  assign _GEN_1458 = 11'h5b2 == WADDR ? 11'h5b2 : _GEN_1457; // @[RAM_ST.scala 31:71]
  assign _GEN_1459 = 11'h5b3 == WADDR ? 11'h5b3 : _GEN_1458; // @[RAM_ST.scala 31:71]
  assign _GEN_1460 = 11'h5b4 == WADDR ? 11'h5b4 : _GEN_1459; // @[RAM_ST.scala 31:71]
  assign _GEN_1461 = 11'h5b5 == WADDR ? 11'h5b5 : _GEN_1460; // @[RAM_ST.scala 31:71]
  assign _GEN_1462 = 11'h5b6 == WADDR ? 11'h5b6 : _GEN_1461; // @[RAM_ST.scala 31:71]
  assign _GEN_1463 = 11'h5b7 == WADDR ? 11'h5b7 : _GEN_1462; // @[RAM_ST.scala 31:71]
  assign _GEN_1464 = 11'h5b8 == WADDR ? 11'h5b8 : _GEN_1463; // @[RAM_ST.scala 31:71]
  assign _GEN_1465 = 11'h5b9 == WADDR ? 11'h5b9 : _GEN_1464; // @[RAM_ST.scala 31:71]
  assign _GEN_1466 = 11'h5ba == WADDR ? 11'h5ba : _GEN_1465; // @[RAM_ST.scala 31:71]
  assign _GEN_1467 = 11'h5bb == WADDR ? 11'h5bb : _GEN_1466; // @[RAM_ST.scala 31:71]
  assign _GEN_1468 = 11'h5bc == WADDR ? 11'h5bc : _GEN_1467; // @[RAM_ST.scala 31:71]
  assign _GEN_1469 = 11'h5bd == WADDR ? 11'h5bd : _GEN_1468; // @[RAM_ST.scala 31:71]
  assign _GEN_1470 = 11'h5be == WADDR ? 11'h5be : _GEN_1469; // @[RAM_ST.scala 31:71]
  assign _GEN_1471 = 11'h5bf == WADDR ? 11'h5bf : _GEN_1470; // @[RAM_ST.scala 31:71]
  assign _GEN_1472 = 11'h5c0 == WADDR ? 11'h5c0 : _GEN_1471; // @[RAM_ST.scala 31:71]
  assign _GEN_1473 = 11'h5c1 == WADDR ? 11'h5c1 : _GEN_1472; // @[RAM_ST.scala 31:71]
  assign _GEN_1474 = 11'h5c2 == WADDR ? 11'h5c2 : _GEN_1473; // @[RAM_ST.scala 31:71]
  assign _GEN_1475 = 11'h5c3 == WADDR ? 11'h5c3 : _GEN_1474; // @[RAM_ST.scala 31:71]
  assign _GEN_1476 = 11'h5c4 == WADDR ? 11'h5c4 : _GEN_1475; // @[RAM_ST.scala 31:71]
  assign _GEN_1477 = 11'h5c5 == WADDR ? 11'h5c5 : _GEN_1476; // @[RAM_ST.scala 31:71]
  assign _GEN_1478 = 11'h5c6 == WADDR ? 11'h5c6 : _GEN_1477; // @[RAM_ST.scala 31:71]
  assign _GEN_1479 = 11'h5c7 == WADDR ? 11'h5c7 : _GEN_1478; // @[RAM_ST.scala 31:71]
  assign _GEN_1480 = 11'h5c8 == WADDR ? 11'h5c8 : _GEN_1479; // @[RAM_ST.scala 31:71]
  assign _GEN_1481 = 11'h5c9 == WADDR ? 11'h5c9 : _GEN_1480; // @[RAM_ST.scala 31:71]
  assign _GEN_1482 = 11'h5ca == WADDR ? 11'h5ca : _GEN_1481; // @[RAM_ST.scala 31:71]
  assign _GEN_1483 = 11'h5cb == WADDR ? 11'h5cb : _GEN_1482; // @[RAM_ST.scala 31:71]
  assign _GEN_1484 = 11'h5cc == WADDR ? 11'h5cc : _GEN_1483; // @[RAM_ST.scala 31:71]
  assign _GEN_1485 = 11'h5cd == WADDR ? 11'h5cd : _GEN_1484; // @[RAM_ST.scala 31:71]
  assign _GEN_1486 = 11'h5ce == WADDR ? 11'h5ce : _GEN_1485; // @[RAM_ST.scala 31:71]
  assign _GEN_1487 = 11'h5cf == WADDR ? 11'h5cf : _GEN_1486; // @[RAM_ST.scala 31:71]
  assign _GEN_1488 = 11'h5d0 == WADDR ? 11'h5d0 : _GEN_1487; // @[RAM_ST.scala 31:71]
  assign _GEN_1489 = 11'h5d1 == WADDR ? 11'h5d1 : _GEN_1488; // @[RAM_ST.scala 31:71]
  assign _GEN_1490 = 11'h5d2 == WADDR ? 11'h5d2 : _GEN_1489; // @[RAM_ST.scala 31:71]
  assign _GEN_1491 = 11'h5d3 == WADDR ? 11'h5d3 : _GEN_1490; // @[RAM_ST.scala 31:71]
  assign _GEN_1492 = 11'h5d4 == WADDR ? 11'h5d4 : _GEN_1491; // @[RAM_ST.scala 31:71]
  assign _GEN_1493 = 11'h5d5 == WADDR ? 11'h5d5 : _GEN_1492; // @[RAM_ST.scala 31:71]
  assign _GEN_1494 = 11'h5d6 == WADDR ? 11'h5d6 : _GEN_1493; // @[RAM_ST.scala 31:71]
  assign _GEN_1495 = 11'h5d7 == WADDR ? 11'h5d7 : _GEN_1494; // @[RAM_ST.scala 31:71]
  assign _GEN_1496 = 11'h5d8 == WADDR ? 11'h5d8 : _GEN_1495; // @[RAM_ST.scala 31:71]
  assign _GEN_1497 = 11'h5d9 == WADDR ? 11'h5d9 : _GEN_1496; // @[RAM_ST.scala 31:71]
  assign _GEN_1498 = 11'h5da == WADDR ? 11'h5da : _GEN_1497; // @[RAM_ST.scala 31:71]
  assign _GEN_1499 = 11'h5db == WADDR ? 11'h5db : _GEN_1498; // @[RAM_ST.scala 31:71]
  assign _GEN_1500 = 11'h5dc == WADDR ? 11'h5dc : _GEN_1499; // @[RAM_ST.scala 31:71]
  assign _GEN_1501 = 11'h5dd == WADDR ? 11'h5dd : _GEN_1500; // @[RAM_ST.scala 31:71]
  assign _GEN_1502 = 11'h5de == WADDR ? 11'h5de : _GEN_1501; // @[RAM_ST.scala 31:71]
  assign _GEN_1503 = 11'h5df == WADDR ? 11'h5df : _GEN_1502; // @[RAM_ST.scala 31:71]
  assign _GEN_1504 = 11'h5e0 == WADDR ? 11'h5e0 : _GEN_1503; // @[RAM_ST.scala 31:71]
  assign _GEN_1505 = 11'h5e1 == WADDR ? 11'h5e1 : _GEN_1504; // @[RAM_ST.scala 31:71]
  assign _GEN_1506 = 11'h5e2 == WADDR ? 11'h5e2 : _GEN_1505; // @[RAM_ST.scala 31:71]
  assign _GEN_1507 = 11'h5e3 == WADDR ? 11'h5e3 : _GEN_1506; // @[RAM_ST.scala 31:71]
  assign _GEN_1508 = 11'h5e4 == WADDR ? 11'h5e4 : _GEN_1507; // @[RAM_ST.scala 31:71]
  assign _GEN_1509 = 11'h5e5 == WADDR ? 11'h5e5 : _GEN_1508; // @[RAM_ST.scala 31:71]
  assign _GEN_1510 = 11'h5e6 == WADDR ? 11'h5e6 : _GEN_1509; // @[RAM_ST.scala 31:71]
  assign _GEN_1511 = 11'h5e7 == WADDR ? 11'h5e7 : _GEN_1510; // @[RAM_ST.scala 31:71]
  assign _GEN_1512 = 11'h5e8 == WADDR ? 11'h5e8 : _GEN_1511; // @[RAM_ST.scala 31:71]
  assign _GEN_1513 = 11'h5e9 == WADDR ? 11'h5e9 : _GEN_1512; // @[RAM_ST.scala 31:71]
  assign _GEN_1514 = 11'h5ea == WADDR ? 11'h5ea : _GEN_1513; // @[RAM_ST.scala 31:71]
  assign _GEN_1515 = 11'h5eb == WADDR ? 11'h5eb : _GEN_1514; // @[RAM_ST.scala 31:71]
  assign _GEN_1516 = 11'h5ec == WADDR ? 11'h5ec : _GEN_1515; // @[RAM_ST.scala 31:71]
  assign _GEN_1517 = 11'h5ed == WADDR ? 11'h5ed : _GEN_1516; // @[RAM_ST.scala 31:71]
  assign _GEN_1518 = 11'h5ee == WADDR ? 11'h5ee : _GEN_1517; // @[RAM_ST.scala 31:71]
  assign _GEN_1519 = 11'h5ef == WADDR ? 11'h5ef : _GEN_1518; // @[RAM_ST.scala 31:71]
  assign _GEN_1520 = 11'h5f0 == WADDR ? 11'h5f0 : _GEN_1519; // @[RAM_ST.scala 31:71]
  assign _GEN_1521 = 11'h5f1 == WADDR ? 11'h5f1 : _GEN_1520; // @[RAM_ST.scala 31:71]
  assign _GEN_1522 = 11'h5f2 == WADDR ? 11'h5f2 : _GEN_1521; // @[RAM_ST.scala 31:71]
  assign _GEN_1523 = 11'h5f3 == WADDR ? 11'h5f3 : _GEN_1522; // @[RAM_ST.scala 31:71]
  assign _GEN_1524 = 11'h5f4 == WADDR ? 11'h5f4 : _GEN_1523; // @[RAM_ST.scala 31:71]
  assign _GEN_1525 = 11'h5f5 == WADDR ? 11'h5f5 : _GEN_1524; // @[RAM_ST.scala 31:71]
  assign _GEN_1526 = 11'h5f6 == WADDR ? 11'h5f6 : _GEN_1525; // @[RAM_ST.scala 31:71]
  assign _GEN_1527 = 11'h5f7 == WADDR ? 11'h5f7 : _GEN_1526; // @[RAM_ST.scala 31:71]
  assign _GEN_1528 = 11'h5f8 == WADDR ? 11'h5f8 : _GEN_1527; // @[RAM_ST.scala 31:71]
  assign _GEN_1529 = 11'h5f9 == WADDR ? 11'h5f9 : _GEN_1528; // @[RAM_ST.scala 31:71]
  assign _GEN_1530 = 11'h5fa == WADDR ? 11'h5fa : _GEN_1529; // @[RAM_ST.scala 31:71]
  assign _GEN_1531 = 11'h5fb == WADDR ? 11'h5fb : _GEN_1530; // @[RAM_ST.scala 31:71]
  assign _GEN_1532 = 11'h5fc == WADDR ? 11'h5fc : _GEN_1531; // @[RAM_ST.scala 31:71]
  assign _GEN_1533 = 11'h5fd == WADDR ? 11'h5fd : _GEN_1532; // @[RAM_ST.scala 31:71]
  assign _GEN_1534 = 11'h5fe == WADDR ? 11'h5fe : _GEN_1533; // @[RAM_ST.scala 31:71]
  assign _GEN_1535 = 11'h5ff == WADDR ? 11'h5ff : _GEN_1534; // @[RAM_ST.scala 31:71]
  assign _GEN_1536 = 11'h600 == WADDR ? 11'h600 : _GEN_1535; // @[RAM_ST.scala 31:71]
  assign _GEN_1537 = 11'h601 == WADDR ? 11'h601 : _GEN_1536; // @[RAM_ST.scala 31:71]
  assign _GEN_1538 = 11'h602 == WADDR ? 11'h602 : _GEN_1537; // @[RAM_ST.scala 31:71]
  assign _GEN_1539 = 11'h603 == WADDR ? 11'h603 : _GEN_1538; // @[RAM_ST.scala 31:71]
  assign _GEN_1540 = 11'h604 == WADDR ? 11'h604 : _GEN_1539; // @[RAM_ST.scala 31:71]
  assign _GEN_1541 = 11'h605 == WADDR ? 11'h605 : _GEN_1540; // @[RAM_ST.scala 31:71]
  assign _GEN_1542 = 11'h606 == WADDR ? 11'h606 : _GEN_1541; // @[RAM_ST.scala 31:71]
  assign _GEN_1543 = 11'h607 == WADDR ? 11'h607 : _GEN_1542; // @[RAM_ST.scala 31:71]
  assign _GEN_1544 = 11'h608 == WADDR ? 11'h608 : _GEN_1543; // @[RAM_ST.scala 31:71]
  assign _GEN_1545 = 11'h609 == WADDR ? 11'h609 : _GEN_1544; // @[RAM_ST.scala 31:71]
  assign _GEN_1546 = 11'h60a == WADDR ? 11'h60a : _GEN_1545; // @[RAM_ST.scala 31:71]
  assign _GEN_1547 = 11'h60b == WADDR ? 11'h60b : _GEN_1546; // @[RAM_ST.scala 31:71]
  assign _GEN_1548 = 11'h60c == WADDR ? 11'h60c : _GEN_1547; // @[RAM_ST.scala 31:71]
  assign _GEN_1549 = 11'h60d == WADDR ? 11'h60d : _GEN_1548; // @[RAM_ST.scala 31:71]
  assign _GEN_1550 = 11'h60e == WADDR ? 11'h60e : _GEN_1549; // @[RAM_ST.scala 31:71]
  assign _GEN_1551 = 11'h60f == WADDR ? 11'h60f : _GEN_1550; // @[RAM_ST.scala 31:71]
  assign _GEN_1552 = 11'h610 == WADDR ? 11'h610 : _GEN_1551; // @[RAM_ST.scala 31:71]
  assign _GEN_1553 = 11'h611 == WADDR ? 11'h611 : _GEN_1552; // @[RAM_ST.scala 31:71]
  assign _GEN_1554 = 11'h612 == WADDR ? 11'h612 : _GEN_1553; // @[RAM_ST.scala 31:71]
  assign _GEN_1555 = 11'h613 == WADDR ? 11'h613 : _GEN_1554; // @[RAM_ST.scala 31:71]
  assign _GEN_1556 = 11'h614 == WADDR ? 11'h614 : _GEN_1555; // @[RAM_ST.scala 31:71]
  assign _GEN_1557 = 11'h615 == WADDR ? 11'h615 : _GEN_1556; // @[RAM_ST.scala 31:71]
  assign _GEN_1558 = 11'h616 == WADDR ? 11'h616 : _GEN_1557; // @[RAM_ST.scala 31:71]
  assign _GEN_1559 = 11'h617 == WADDR ? 11'h617 : _GEN_1558; // @[RAM_ST.scala 31:71]
  assign _GEN_1560 = 11'h618 == WADDR ? 11'h618 : _GEN_1559; // @[RAM_ST.scala 31:71]
  assign _GEN_1561 = 11'h619 == WADDR ? 11'h619 : _GEN_1560; // @[RAM_ST.scala 31:71]
  assign _GEN_1562 = 11'h61a == WADDR ? 11'h61a : _GEN_1561; // @[RAM_ST.scala 31:71]
  assign _GEN_1563 = 11'h61b == WADDR ? 11'h61b : _GEN_1562; // @[RAM_ST.scala 31:71]
  assign _GEN_1564 = 11'h61c == WADDR ? 11'h61c : _GEN_1563; // @[RAM_ST.scala 31:71]
  assign _GEN_1565 = 11'h61d == WADDR ? 11'h61d : _GEN_1564; // @[RAM_ST.scala 31:71]
  assign _GEN_1566 = 11'h61e == WADDR ? 11'h61e : _GEN_1565; // @[RAM_ST.scala 31:71]
  assign _GEN_1567 = 11'h61f == WADDR ? 11'h61f : _GEN_1566; // @[RAM_ST.scala 31:71]
  assign _GEN_1568 = 11'h620 == WADDR ? 11'h620 : _GEN_1567; // @[RAM_ST.scala 31:71]
  assign _GEN_1569 = 11'h621 == WADDR ? 11'h621 : _GEN_1568; // @[RAM_ST.scala 31:71]
  assign _GEN_1570 = 11'h622 == WADDR ? 11'h622 : _GEN_1569; // @[RAM_ST.scala 31:71]
  assign _GEN_1571 = 11'h623 == WADDR ? 11'h623 : _GEN_1570; // @[RAM_ST.scala 31:71]
  assign _GEN_1572 = 11'h624 == WADDR ? 11'h624 : _GEN_1571; // @[RAM_ST.scala 31:71]
  assign _GEN_1573 = 11'h625 == WADDR ? 11'h625 : _GEN_1572; // @[RAM_ST.scala 31:71]
  assign _GEN_1574 = 11'h626 == WADDR ? 11'h626 : _GEN_1573; // @[RAM_ST.scala 31:71]
  assign _GEN_1575 = 11'h627 == WADDR ? 11'h627 : _GEN_1574; // @[RAM_ST.scala 31:71]
  assign _GEN_1576 = 11'h628 == WADDR ? 11'h628 : _GEN_1575; // @[RAM_ST.scala 31:71]
  assign _GEN_1577 = 11'h629 == WADDR ? 11'h629 : _GEN_1576; // @[RAM_ST.scala 31:71]
  assign _GEN_1578 = 11'h62a == WADDR ? 11'h62a : _GEN_1577; // @[RAM_ST.scala 31:71]
  assign _GEN_1579 = 11'h62b == WADDR ? 11'h62b : _GEN_1578; // @[RAM_ST.scala 31:71]
  assign _GEN_1580 = 11'h62c == WADDR ? 11'h62c : _GEN_1579; // @[RAM_ST.scala 31:71]
  assign _GEN_1581 = 11'h62d == WADDR ? 11'h62d : _GEN_1580; // @[RAM_ST.scala 31:71]
  assign _GEN_1582 = 11'h62e == WADDR ? 11'h62e : _GEN_1581; // @[RAM_ST.scala 31:71]
  assign _GEN_1583 = 11'h62f == WADDR ? 11'h62f : _GEN_1582; // @[RAM_ST.scala 31:71]
  assign _GEN_1584 = 11'h630 == WADDR ? 11'h630 : _GEN_1583; // @[RAM_ST.scala 31:71]
  assign _GEN_1585 = 11'h631 == WADDR ? 11'h631 : _GEN_1584; // @[RAM_ST.scala 31:71]
  assign _GEN_1586 = 11'h632 == WADDR ? 11'h632 : _GEN_1585; // @[RAM_ST.scala 31:71]
  assign _GEN_1587 = 11'h633 == WADDR ? 11'h633 : _GEN_1586; // @[RAM_ST.scala 31:71]
  assign _GEN_1588 = 11'h634 == WADDR ? 11'h634 : _GEN_1587; // @[RAM_ST.scala 31:71]
  assign _GEN_1589 = 11'h635 == WADDR ? 11'h635 : _GEN_1588; // @[RAM_ST.scala 31:71]
  assign _GEN_1590 = 11'h636 == WADDR ? 11'h636 : _GEN_1589; // @[RAM_ST.scala 31:71]
  assign _GEN_1591 = 11'h637 == WADDR ? 11'h637 : _GEN_1590; // @[RAM_ST.scala 31:71]
  assign _GEN_1592 = 11'h638 == WADDR ? 11'h638 : _GEN_1591; // @[RAM_ST.scala 31:71]
  assign _GEN_1593 = 11'h639 == WADDR ? 11'h639 : _GEN_1592; // @[RAM_ST.scala 31:71]
  assign _GEN_1594 = 11'h63a == WADDR ? 11'h63a : _GEN_1593; // @[RAM_ST.scala 31:71]
  assign _GEN_1595 = 11'h63b == WADDR ? 11'h63b : _GEN_1594; // @[RAM_ST.scala 31:71]
  assign _GEN_1596 = 11'h63c == WADDR ? 11'h63c : _GEN_1595; // @[RAM_ST.scala 31:71]
  assign _GEN_1597 = 11'h63d == WADDR ? 11'h63d : _GEN_1596; // @[RAM_ST.scala 31:71]
  assign _GEN_1598 = 11'h63e == WADDR ? 11'h63e : _GEN_1597; // @[RAM_ST.scala 31:71]
  assign _GEN_1599 = 11'h63f == WADDR ? 11'h63f : _GEN_1598; // @[RAM_ST.scala 31:71]
  assign _GEN_1600 = 11'h640 == WADDR ? 11'h640 : _GEN_1599; // @[RAM_ST.scala 31:71]
  assign _GEN_1601 = 11'h641 == WADDR ? 11'h641 : _GEN_1600; // @[RAM_ST.scala 31:71]
  assign _GEN_1602 = 11'h642 == WADDR ? 11'h642 : _GEN_1601; // @[RAM_ST.scala 31:71]
  assign _GEN_1603 = 11'h643 == WADDR ? 11'h643 : _GEN_1602; // @[RAM_ST.scala 31:71]
  assign _GEN_1604 = 11'h644 == WADDR ? 11'h644 : _GEN_1603; // @[RAM_ST.scala 31:71]
  assign _GEN_1605 = 11'h645 == WADDR ? 11'h645 : _GEN_1604; // @[RAM_ST.scala 31:71]
  assign _GEN_1606 = 11'h646 == WADDR ? 11'h646 : _GEN_1605; // @[RAM_ST.scala 31:71]
  assign _GEN_1607 = 11'h647 == WADDR ? 11'h647 : _GEN_1606; // @[RAM_ST.scala 31:71]
  assign _GEN_1608 = 11'h648 == WADDR ? 11'h648 : _GEN_1607; // @[RAM_ST.scala 31:71]
  assign _GEN_1609 = 11'h649 == WADDR ? 11'h649 : _GEN_1608; // @[RAM_ST.scala 31:71]
  assign _GEN_1610 = 11'h64a == WADDR ? 11'h64a : _GEN_1609; // @[RAM_ST.scala 31:71]
  assign _GEN_1611 = 11'h64b == WADDR ? 11'h64b : _GEN_1610; // @[RAM_ST.scala 31:71]
  assign _GEN_1612 = 11'h64c == WADDR ? 11'h64c : _GEN_1611; // @[RAM_ST.scala 31:71]
  assign _GEN_1613 = 11'h64d == WADDR ? 11'h64d : _GEN_1612; // @[RAM_ST.scala 31:71]
  assign _GEN_1614 = 11'h64e == WADDR ? 11'h64e : _GEN_1613; // @[RAM_ST.scala 31:71]
  assign _GEN_1615 = 11'h64f == WADDR ? 11'h64f : _GEN_1614; // @[RAM_ST.scala 31:71]
  assign _GEN_1616 = 11'h650 == WADDR ? 11'h650 : _GEN_1615; // @[RAM_ST.scala 31:71]
  assign _GEN_1617 = 11'h651 == WADDR ? 11'h651 : _GEN_1616; // @[RAM_ST.scala 31:71]
  assign _GEN_1618 = 11'h652 == WADDR ? 11'h652 : _GEN_1617; // @[RAM_ST.scala 31:71]
  assign _GEN_1619 = 11'h653 == WADDR ? 11'h653 : _GEN_1618; // @[RAM_ST.scala 31:71]
  assign _GEN_1620 = 11'h654 == WADDR ? 11'h654 : _GEN_1619; // @[RAM_ST.scala 31:71]
  assign _GEN_1621 = 11'h655 == WADDR ? 11'h655 : _GEN_1620; // @[RAM_ST.scala 31:71]
  assign _GEN_1622 = 11'h656 == WADDR ? 11'h656 : _GEN_1621; // @[RAM_ST.scala 31:71]
  assign _GEN_1623 = 11'h657 == WADDR ? 11'h657 : _GEN_1622; // @[RAM_ST.scala 31:71]
  assign _GEN_1624 = 11'h658 == WADDR ? 11'h658 : _GEN_1623; // @[RAM_ST.scala 31:71]
  assign _GEN_1625 = 11'h659 == WADDR ? 11'h659 : _GEN_1624; // @[RAM_ST.scala 31:71]
  assign _GEN_1626 = 11'h65a == WADDR ? 11'h65a : _GEN_1625; // @[RAM_ST.scala 31:71]
  assign _GEN_1627 = 11'h65b == WADDR ? 11'h65b : _GEN_1626; // @[RAM_ST.scala 31:71]
  assign _GEN_1628 = 11'h65c == WADDR ? 11'h65c : _GEN_1627; // @[RAM_ST.scala 31:71]
  assign _GEN_1629 = 11'h65d == WADDR ? 11'h65d : _GEN_1628; // @[RAM_ST.scala 31:71]
  assign _GEN_1630 = 11'h65e == WADDR ? 11'h65e : _GEN_1629; // @[RAM_ST.scala 31:71]
  assign _GEN_1631 = 11'h65f == WADDR ? 11'h65f : _GEN_1630; // @[RAM_ST.scala 31:71]
  assign _GEN_1632 = 11'h660 == WADDR ? 11'h660 : _GEN_1631; // @[RAM_ST.scala 31:71]
  assign _GEN_1633 = 11'h661 == WADDR ? 11'h661 : _GEN_1632; // @[RAM_ST.scala 31:71]
  assign _GEN_1634 = 11'h662 == WADDR ? 11'h662 : _GEN_1633; // @[RAM_ST.scala 31:71]
  assign _GEN_1635 = 11'h663 == WADDR ? 11'h663 : _GEN_1634; // @[RAM_ST.scala 31:71]
  assign _GEN_1636 = 11'h664 == WADDR ? 11'h664 : _GEN_1635; // @[RAM_ST.scala 31:71]
  assign _GEN_1637 = 11'h665 == WADDR ? 11'h665 : _GEN_1636; // @[RAM_ST.scala 31:71]
  assign _GEN_1638 = 11'h666 == WADDR ? 11'h666 : _GEN_1637; // @[RAM_ST.scala 31:71]
  assign _GEN_1639 = 11'h667 == WADDR ? 11'h667 : _GEN_1638; // @[RAM_ST.scala 31:71]
  assign _GEN_1640 = 11'h668 == WADDR ? 11'h668 : _GEN_1639; // @[RAM_ST.scala 31:71]
  assign _GEN_1641 = 11'h669 == WADDR ? 11'h669 : _GEN_1640; // @[RAM_ST.scala 31:71]
  assign _GEN_1642 = 11'h66a == WADDR ? 11'h66a : _GEN_1641; // @[RAM_ST.scala 31:71]
  assign _GEN_1643 = 11'h66b == WADDR ? 11'h66b : _GEN_1642; // @[RAM_ST.scala 31:71]
  assign _GEN_1644 = 11'h66c == WADDR ? 11'h66c : _GEN_1643; // @[RAM_ST.scala 31:71]
  assign _GEN_1645 = 11'h66d == WADDR ? 11'h66d : _GEN_1644; // @[RAM_ST.scala 31:71]
  assign _GEN_1646 = 11'h66e == WADDR ? 11'h66e : _GEN_1645; // @[RAM_ST.scala 31:71]
  assign _GEN_1647 = 11'h66f == WADDR ? 11'h66f : _GEN_1646; // @[RAM_ST.scala 31:71]
  assign _GEN_1648 = 11'h670 == WADDR ? 11'h670 : _GEN_1647; // @[RAM_ST.scala 31:71]
  assign _GEN_1649 = 11'h671 == WADDR ? 11'h671 : _GEN_1648; // @[RAM_ST.scala 31:71]
  assign _GEN_1650 = 11'h672 == WADDR ? 11'h672 : _GEN_1649; // @[RAM_ST.scala 31:71]
  assign _GEN_1651 = 11'h673 == WADDR ? 11'h673 : _GEN_1650; // @[RAM_ST.scala 31:71]
  assign _GEN_1652 = 11'h674 == WADDR ? 11'h674 : _GEN_1651; // @[RAM_ST.scala 31:71]
  assign _GEN_1653 = 11'h675 == WADDR ? 11'h675 : _GEN_1652; // @[RAM_ST.scala 31:71]
  assign _GEN_1654 = 11'h676 == WADDR ? 11'h676 : _GEN_1653; // @[RAM_ST.scala 31:71]
  assign _GEN_1655 = 11'h677 == WADDR ? 11'h677 : _GEN_1654; // @[RAM_ST.scala 31:71]
  assign _GEN_1656 = 11'h678 == WADDR ? 11'h678 : _GEN_1655; // @[RAM_ST.scala 31:71]
  assign _GEN_1657 = 11'h679 == WADDR ? 11'h679 : _GEN_1656; // @[RAM_ST.scala 31:71]
  assign _GEN_1658 = 11'h67a == WADDR ? 11'h67a : _GEN_1657; // @[RAM_ST.scala 31:71]
  assign _GEN_1659 = 11'h67b == WADDR ? 11'h67b : _GEN_1658; // @[RAM_ST.scala 31:71]
  assign _GEN_1660 = 11'h67c == WADDR ? 11'h67c : _GEN_1659; // @[RAM_ST.scala 31:71]
  assign _GEN_1661 = 11'h67d == WADDR ? 11'h67d : _GEN_1660; // @[RAM_ST.scala 31:71]
  assign _GEN_1662 = 11'h67e == WADDR ? 11'h67e : _GEN_1661; // @[RAM_ST.scala 31:71]
  assign _GEN_1663 = 11'h67f == WADDR ? 11'h67f : _GEN_1662; // @[RAM_ST.scala 31:71]
  assign _GEN_1664 = 11'h680 == WADDR ? 11'h680 : _GEN_1663; // @[RAM_ST.scala 31:71]
  assign _GEN_1665 = 11'h681 == WADDR ? 11'h681 : _GEN_1664; // @[RAM_ST.scala 31:71]
  assign _GEN_1666 = 11'h682 == WADDR ? 11'h682 : _GEN_1665; // @[RAM_ST.scala 31:71]
  assign _GEN_1667 = 11'h683 == WADDR ? 11'h683 : _GEN_1666; // @[RAM_ST.scala 31:71]
  assign _GEN_1668 = 11'h684 == WADDR ? 11'h684 : _GEN_1667; // @[RAM_ST.scala 31:71]
  assign _GEN_1669 = 11'h685 == WADDR ? 11'h685 : _GEN_1668; // @[RAM_ST.scala 31:71]
  assign _GEN_1670 = 11'h686 == WADDR ? 11'h686 : _GEN_1669; // @[RAM_ST.scala 31:71]
  assign _GEN_1671 = 11'h687 == WADDR ? 11'h687 : _GEN_1670; // @[RAM_ST.scala 31:71]
  assign _GEN_1672 = 11'h688 == WADDR ? 11'h688 : _GEN_1671; // @[RAM_ST.scala 31:71]
  assign _GEN_1673 = 11'h689 == WADDR ? 11'h689 : _GEN_1672; // @[RAM_ST.scala 31:71]
  assign _GEN_1674 = 11'h68a == WADDR ? 11'h68a : _GEN_1673; // @[RAM_ST.scala 31:71]
  assign _GEN_1675 = 11'h68b == WADDR ? 11'h68b : _GEN_1674; // @[RAM_ST.scala 31:71]
  assign _GEN_1676 = 11'h68c == WADDR ? 11'h68c : _GEN_1675; // @[RAM_ST.scala 31:71]
  assign _GEN_1677 = 11'h68d == WADDR ? 11'h68d : _GEN_1676; // @[RAM_ST.scala 31:71]
  assign _GEN_1678 = 11'h68e == WADDR ? 11'h68e : _GEN_1677; // @[RAM_ST.scala 31:71]
  assign _GEN_1679 = 11'h68f == WADDR ? 11'h68f : _GEN_1678; // @[RAM_ST.scala 31:71]
  assign _GEN_1680 = 11'h690 == WADDR ? 11'h690 : _GEN_1679; // @[RAM_ST.scala 31:71]
  assign _GEN_1681 = 11'h691 == WADDR ? 11'h691 : _GEN_1680; // @[RAM_ST.scala 31:71]
  assign _GEN_1682 = 11'h692 == WADDR ? 11'h692 : _GEN_1681; // @[RAM_ST.scala 31:71]
  assign _GEN_1683 = 11'h693 == WADDR ? 11'h693 : _GEN_1682; // @[RAM_ST.scala 31:71]
  assign _GEN_1684 = 11'h694 == WADDR ? 11'h694 : _GEN_1683; // @[RAM_ST.scala 31:71]
  assign _GEN_1685 = 11'h695 == WADDR ? 11'h695 : _GEN_1684; // @[RAM_ST.scala 31:71]
  assign _GEN_1686 = 11'h696 == WADDR ? 11'h696 : _GEN_1685; // @[RAM_ST.scala 31:71]
  assign _GEN_1687 = 11'h697 == WADDR ? 11'h697 : _GEN_1686; // @[RAM_ST.scala 31:71]
  assign _GEN_1688 = 11'h698 == WADDR ? 11'h698 : _GEN_1687; // @[RAM_ST.scala 31:71]
  assign _GEN_1689 = 11'h699 == WADDR ? 11'h699 : _GEN_1688; // @[RAM_ST.scala 31:71]
  assign _GEN_1690 = 11'h69a == WADDR ? 11'h69a : _GEN_1689; // @[RAM_ST.scala 31:71]
  assign _GEN_1691 = 11'h69b == WADDR ? 11'h69b : _GEN_1690; // @[RAM_ST.scala 31:71]
  assign _GEN_1692 = 11'h69c == WADDR ? 11'h69c : _GEN_1691; // @[RAM_ST.scala 31:71]
  assign _GEN_1693 = 11'h69d == WADDR ? 11'h69d : _GEN_1692; // @[RAM_ST.scala 31:71]
  assign _GEN_1694 = 11'h69e == WADDR ? 11'h69e : _GEN_1693; // @[RAM_ST.scala 31:71]
  assign _GEN_1695 = 11'h69f == WADDR ? 11'h69f : _GEN_1694; // @[RAM_ST.scala 31:71]
  assign _GEN_1696 = 11'h6a0 == WADDR ? 11'h6a0 : _GEN_1695; // @[RAM_ST.scala 31:71]
  assign _GEN_1697 = 11'h6a1 == WADDR ? 11'h6a1 : _GEN_1696; // @[RAM_ST.scala 31:71]
  assign _GEN_1698 = 11'h6a2 == WADDR ? 11'h6a2 : _GEN_1697; // @[RAM_ST.scala 31:71]
  assign _GEN_1699 = 11'h6a3 == WADDR ? 11'h6a3 : _GEN_1698; // @[RAM_ST.scala 31:71]
  assign _GEN_1700 = 11'h6a4 == WADDR ? 11'h6a4 : _GEN_1699; // @[RAM_ST.scala 31:71]
  assign _GEN_1701 = 11'h6a5 == WADDR ? 11'h6a5 : _GEN_1700; // @[RAM_ST.scala 31:71]
  assign _GEN_1702 = 11'h6a6 == WADDR ? 11'h6a6 : _GEN_1701; // @[RAM_ST.scala 31:71]
  assign _GEN_1703 = 11'h6a7 == WADDR ? 11'h6a7 : _GEN_1702; // @[RAM_ST.scala 31:71]
  assign _GEN_1704 = 11'h6a8 == WADDR ? 11'h6a8 : _GEN_1703; // @[RAM_ST.scala 31:71]
  assign _GEN_1705 = 11'h6a9 == WADDR ? 11'h6a9 : _GEN_1704; // @[RAM_ST.scala 31:71]
  assign _GEN_1706 = 11'h6aa == WADDR ? 11'h6aa : _GEN_1705; // @[RAM_ST.scala 31:71]
  assign _GEN_1707 = 11'h6ab == WADDR ? 11'h6ab : _GEN_1706; // @[RAM_ST.scala 31:71]
  assign _GEN_1708 = 11'h6ac == WADDR ? 11'h6ac : _GEN_1707; // @[RAM_ST.scala 31:71]
  assign _GEN_1709 = 11'h6ad == WADDR ? 11'h6ad : _GEN_1708; // @[RAM_ST.scala 31:71]
  assign _GEN_1710 = 11'h6ae == WADDR ? 11'h6ae : _GEN_1709; // @[RAM_ST.scala 31:71]
  assign _GEN_1711 = 11'h6af == WADDR ? 11'h6af : _GEN_1710; // @[RAM_ST.scala 31:71]
  assign _GEN_1712 = 11'h6b0 == WADDR ? 11'h6b0 : _GEN_1711; // @[RAM_ST.scala 31:71]
  assign _GEN_1713 = 11'h6b1 == WADDR ? 11'h6b1 : _GEN_1712; // @[RAM_ST.scala 31:71]
  assign _GEN_1714 = 11'h6b2 == WADDR ? 11'h6b2 : _GEN_1713; // @[RAM_ST.scala 31:71]
  assign _GEN_1715 = 11'h6b3 == WADDR ? 11'h6b3 : _GEN_1714; // @[RAM_ST.scala 31:71]
  assign _GEN_1716 = 11'h6b4 == WADDR ? 11'h6b4 : _GEN_1715; // @[RAM_ST.scala 31:71]
  assign _GEN_1717 = 11'h6b5 == WADDR ? 11'h6b5 : _GEN_1716; // @[RAM_ST.scala 31:71]
  assign _GEN_1718 = 11'h6b6 == WADDR ? 11'h6b6 : _GEN_1717; // @[RAM_ST.scala 31:71]
  assign _GEN_1719 = 11'h6b7 == WADDR ? 11'h6b7 : _GEN_1718; // @[RAM_ST.scala 31:71]
  assign _GEN_1720 = 11'h6b8 == WADDR ? 11'h6b8 : _GEN_1719; // @[RAM_ST.scala 31:71]
  assign _GEN_1721 = 11'h6b9 == WADDR ? 11'h6b9 : _GEN_1720; // @[RAM_ST.scala 31:71]
  assign _GEN_1722 = 11'h6ba == WADDR ? 11'h6ba : _GEN_1721; // @[RAM_ST.scala 31:71]
  assign _GEN_1723 = 11'h6bb == WADDR ? 11'h6bb : _GEN_1722; // @[RAM_ST.scala 31:71]
  assign _GEN_1724 = 11'h6bc == WADDR ? 11'h6bc : _GEN_1723; // @[RAM_ST.scala 31:71]
  assign _GEN_1725 = 11'h6bd == WADDR ? 11'h6bd : _GEN_1724; // @[RAM_ST.scala 31:71]
  assign _GEN_1726 = 11'h6be == WADDR ? 11'h6be : _GEN_1725; // @[RAM_ST.scala 31:71]
  assign _GEN_1727 = 11'h6bf == WADDR ? 11'h6bf : _GEN_1726; // @[RAM_ST.scala 31:71]
  assign _GEN_1728 = 11'h6c0 == WADDR ? 11'h6c0 : _GEN_1727; // @[RAM_ST.scala 31:71]
  assign _GEN_1729 = 11'h6c1 == WADDR ? 11'h6c1 : _GEN_1728; // @[RAM_ST.scala 31:71]
  assign _GEN_1730 = 11'h6c2 == WADDR ? 11'h6c2 : _GEN_1729; // @[RAM_ST.scala 31:71]
  assign _GEN_1731 = 11'h6c3 == WADDR ? 11'h6c3 : _GEN_1730; // @[RAM_ST.scala 31:71]
  assign _GEN_1732 = 11'h6c4 == WADDR ? 11'h6c4 : _GEN_1731; // @[RAM_ST.scala 31:71]
  assign _GEN_1733 = 11'h6c5 == WADDR ? 11'h6c5 : _GEN_1732; // @[RAM_ST.scala 31:71]
  assign _GEN_1734 = 11'h6c6 == WADDR ? 11'h6c6 : _GEN_1733; // @[RAM_ST.scala 31:71]
  assign _GEN_1735 = 11'h6c7 == WADDR ? 11'h6c7 : _GEN_1734; // @[RAM_ST.scala 31:71]
  assign _GEN_1736 = 11'h6c8 == WADDR ? 11'h6c8 : _GEN_1735; // @[RAM_ST.scala 31:71]
  assign _GEN_1737 = 11'h6c9 == WADDR ? 11'h6c9 : _GEN_1736; // @[RAM_ST.scala 31:71]
  assign _GEN_1738 = 11'h6ca == WADDR ? 11'h6ca : _GEN_1737; // @[RAM_ST.scala 31:71]
  assign _GEN_1739 = 11'h6cb == WADDR ? 11'h6cb : _GEN_1738; // @[RAM_ST.scala 31:71]
  assign _GEN_1740 = 11'h6cc == WADDR ? 11'h6cc : _GEN_1739; // @[RAM_ST.scala 31:71]
  assign _GEN_1741 = 11'h6cd == WADDR ? 11'h6cd : _GEN_1740; // @[RAM_ST.scala 31:71]
  assign _GEN_1742 = 11'h6ce == WADDR ? 11'h6ce : _GEN_1741; // @[RAM_ST.scala 31:71]
  assign _GEN_1743 = 11'h6cf == WADDR ? 11'h6cf : _GEN_1742; // @[RAM_ST.scala 31:71]
  assign _GEN_1744 = 11'h6d0 == WADDR ? 11'h6d0 : _GEN_1743; // @[RAM_ST.scala 31:71]
  assign _GEN_1745 = 11'h6d1 == WADDR ? 11'h6d1 : _GEN_1744; // @[RAM_ST.scala 31:71]
  assign _GEN_1746 = 11'h6d2 == WADDR ? 11'h6d2 : _GEN_1745; // @[RAM_ST.scala 31:71]
  assign _GEN_1747 = 11'h6d3 == WADDR ? 11'h6d3 : _GEN_1746; // @[RAM_ST.scala 31:71]
  assign _GEN_1748 = 11'h6d4 == WADDR ? 11'h6d4 : _GEN_1747; // @[RAM_ST.scala 31:71]
  assign _GEN_1749 = 11'h6d5 == WADDR ? 11'h6d5 : _GEN_1748; // @[RAM_ST.scala 31:71]
  assign _GEN_1750 = 11'h6d6 == WADDR ? 11'h6d6 : _GEN_1749; // @[RAM_ST.scala 31:71]
  assign _GEN_1751 = 11'h6d7 == WADDR ? 11'h6d7 : _GEN_1750; // @[RAM_ST.scala 31:71]
  assign _GEN_1752 = 11'h6d8 == WADDR ? 11'h6d8 : _GEN_1751; // @[RAM_ST.scala 31:71]
  assign _GEN_1753 = 11'h6d9 == WADDR ? 11'h6d9 : _GEN_1752; // @[RAM_ST.scala 31:71]
  assign _GEN_1754 = 11'h6da == WADDR ? 11'h6da : _GEN_1753; // @[RAM_ST.scala 31:71]
  assign _GEN_1755 = 11'h6db == WADDR ? 11'h6db : _GEN_1754; // @[RAM_ST.scala 31:71]
  assign _GEN_1756 = 11'h6dc == WADDR ? 11'h6dc : _GEN_1755; // @[RAM_ST.scala 31:71]
  assign _GEN_1757 = 11'h6dd == WADDR ? 11'h6dd : _GEN_1756; // @[RAM_ST.scala 31:71]
  assign _GEN_1758 = 11'h6de == WADDR ? 11'h6de : _GEN_1757; // @[RAM_ST.scala 31:71]
  assign _GEN_1759 = 11'h6df == WADDR ? 11'h6df : _GEN_1758; // @[RAM_ST.scala 31:71]
  assign _GEN_1760 = 11'h6e0 == WADDR ? 11'h6e0 : _GEN_1759; // @[RAM_ST.scala 31:71]
  assign _GEN_1761 = 11'h6e1 == WADDR ? 11'h6e1 : _GEN_1760; // @[RAM_ST.scala 31:71]
  assign _GEN_1762 = 11'h6e2 == WADDR ? 11'h6e2 : _GEN_1761; // @[RAM_ST.scala 31:71]
  assign _GEN_1763 = 11'h6e3 == WADDR ? 11'h6e3 : _GEN_1762; // @[RAM_ST.scala 31:71]
  assign _GEN_1764 = 11'h6e4 == WADDR ? 11'h6e4 : _GEN_1763; // @[RAM_ST.scala 31:71]
  assign _GEN_1765 = 11'h6e5 == WADDR ? 11'h6e5 : _GEN_1764; // @[RAM_ST.scala 31:71]
  assign _GEN_1766 = 11'h6e6 == WADDR ? 11'h6e6 : _GEN_1765; // @[RAM_ST.scala 31:71]
  assign _GEN_1767 = 11'h6e7 == WADDR ? 11'h6e7 : _GEN_1766; // @[RAM_ST.scala 31:71]
  assign _GEN_1768 = 11'h6e8 == WADDR ? 11'h6e8 : _GEN_1767; // @[RAM_ST.scala 31:71]
  assign _GEN_1769 = 11'h6e9 == WADDR ? 11'h6e9 : _GEN_1768; // @[RAM_ST.scala 31:71]
  assign _GEN_1770 = 11'h6ea == WADDR ? 11'h6ea : _GEN_1769; // @[RAM_ST.scala 31:71]
  assign _GEN_1771 = 11'h6eb == WADDR ? 11'h6eb : _GEN_1770; // @[RAM_ST.scala 31:71]
  assign _GEN_1772 = 11'h6ec == WADDR ? 11'h6ec : _GEN_1771; // @[RAM_ST.scala 31:71]
  assign _GEN_1773 = 11'h6ed == WADDR ? 11'h6ed : _GEN_1772; // @[RAM_ST.scala 31:71]
  assign _GEN_1774 = 11'h6ee == WADDR ? 11'h6ee : _GEN_1773; // @[RAM_ST.scala 31:71]
  assign _GEN_1775 = 11'h6ef == WADDR ? 11'h6ef : _GEN_1774; // @[RAM_ST.scala 31:71]
  assign _GEN_1776 = 11'h6f0 == WADDR ? 11'h6f0 : _GEN_1775; // @[RAM_ST.scala 31:71]
  assign _GEN_1777 = 11'h6f1 == WADDR ? 11'h6f1 : _GEN_1776; // @[RAM_ST.scala 31:71]
  assign _GEN_1778 = 11'h6f2 == WADDR ? 11'h6f2 : _GEN_1777; // @[RAM_ST.scala 31:71]
  assign _GEN_1779 = 11'h6f3 == WADDR ? 11'h6f3 : _GEN_1778; // @[RAM_ST.scala 31:71]
  assign _GEN_1780 = 11'h6f4 == WADDR ? 11'h6f4 : _GEN_1779; // @[RAM_ST.scala 31:71]
  assign _GEN_1781 = 11'h6f5 == WADDR ? 11'h6f5 : _GEN_1780; // @[RAM_ST.scala 31:71]
  assign _GEN_1782 = 11'h6f6 == WADDR ? 11'h6f6 : _GEN_1781; // @[RAM_ST.scala 31:71]
  assign _GEN_1783 = 11'h6f7 == WADDR ? 11'h6f7 : _GEN_1782; // @[RAM_ST.scala 31:71]
  assign _GEN_1784 = 11'h6f8 == WADDR ? 11'h6f8 : _GEN_1783; // @[RAM_ST.scala 31:71]
  assign _GEN_1785 = 11'h6f9 == WADDR ? 11'h6f9 : _GEN_1784; // @[RAM_ST.scala 31:71]
  assign _GEN_1786 = 11'h6fa == WADDR ? 11'h6fa : _GEN_1785; // @[RAM_ST.scala 31:71]
  assign _GEN_1787 = 11'h6fb == WADDR ? 11'h6fb : _GEN_1786; // @[RAM_ST.scala 31:71]
  assign _GEN_1788 = 11'h6fc == WADDR ? 11'h6fc : _GEN_1787; // @[RAM_ST.scala 31:71]
  assign _GEN_1789 = 11'h6fd == WADDR ? 11'h6fd : _GEN_1788; // @[RAM_ST.scala 31:71]
  assign _GEN_1790 = 11'h6fe == WADDR ? 11'h6fe : _GEN_1789; // @[RAM_ST.scala 31:71]
  assign _GEN_1791 = 11'h6ff == WADDR ? 11'h6ff : _GEN_1790; // @[RAM_ST.scala 31:71]
  assign _GEN_1792 = 11'h700 == WADDR ? 11'h700 : _GEN_1791; // @[RAM_ST.scala 31:71]
  assign _GEN_1793 = 11'h701 == WADDR ? 11'h701 : _GEN_1792; // @[RAM_ST.scala 31:71]
  assign _GEN_1794 = 11'h702 == WADDR ? 11'h702 : _GEN_1793; // @[RAM_ST.scala 31:71]
  assign _GEN_1795 = 11'h703 == WADDR ? 11'h703 : _GEN_1794; // @[RAM_ST.scala 31:71]
  assign _GEN_1796 = 11'h704 == WADDR ? 11'h704 : _GEN_1795; // @[RAM_ST.scala 31:71]
  assign _GEN_1797 = 11'h705 == WADDR ? 11'h705 : _GEN_1796; // @[RAM_ST.scala 31:71]
  assign _GEN_1798 = 11'h706 == WADDR ? 11'h706 : _GEN_1797; // @[RAM_ST.scala 31:71]
  assign _GEN_1799 = 11'h707 == WADDR ? 11'h707 : _GEN_1798; // @[RAM_ST.scala 31:71]
  assign _GEN_1800 = 11'h708 == WADDR ? 11'h708 : _GEN_1799; // @[RAM_ST.scala 31:71]
  assign _GEN_1801 = 11'h709 == WADDR ? 11'h709 : _GEN_1800; // @[RAM_ST.scala 31:71]
  assign _GEN_1802 = 11'h70a == WADDR ? 11'h70a : _GEN_1801; // @[RAM_ST.scala 31:71]
  assign _GEN_1803 = 11'h70b == WADDR ? 11'h70b : _GEN_1802; // @[RAM_ST.scala 31:71]
  assign _GEN_1804 = 11'h70c == WADDR ? 11'h70c : _GEN_1803; // @[RAM_ST.scala 31:71]
  assign _GEN_1805 = 11'h70d == WADDR ? 11'h70d : _GEN_1804; // @[RAM_ST.scala 31:71]
  assign _GEN_1806 = 11'h70e == WADDR ? 11'h70e : _GEN_1805; // @[RAM_ST.scala 31:71]
  assign _GEN_1807 = 11'h70f == WADDR ? 11'h70f : _GEN_1806; // @[RAM_ST.scala 31:71]
  assign _GEN_1808 = 11'h710 == WADDR ? 11'h710 : _GEN_1807; // @[RAM_ST.scala 31:71]
  assign _GEN_1809 = 11'h711 == WADDR ? 11'h711 : _GEN_1808; // @[RAM_ST.scala 31:71]
  assign _GEN_1810 = 11'h712 == WADDR ? 11'h712 : _GEN_1809; // @[RAM_ST.scala 31:71]
  assign _GEN_1811 = 11'h713 == WADDR ? 11'h713 : _GEN_1810; // @[RAM_ST.scala 31:71]
  assign _GEN_1812 = 11'h714 == WADDR ? 11'h714 : _GEN_1811; // @[RAM_ST.scala 31:71]
  assign _GEN_1813 = 11'h715 == WADDR ? 11'h715 : _GEN_1812; // @[RAM_ST.scala 31:71]
  assign _GEN_1814 = 11'h716 == WADDR ? 11'h716 : _GEN_1813; // @[RAM_ST.scala 31:71]
  assign _GEN_1815 = 11'h717 == WADDR ? 11'h717 : _GEN_1814; // @[RAM_ST.scala 31:71]
  assign _GEN_1816 = 11'h718 == WADDR ? 11'h718 : _GEN_1815; // @[RAM_ST.scala 31:71]
  assign _GEN_1817 = 11'h719 == WADDR ? 11'h719 : _GEN_1816; // @[RAM_ST.scala 31:71]
  assign _GEN_1818 = 11'h71a == WADDR ? 11'h71a : _GEN_1817; // @[RAM_ST.scala 31:71]
  assign _GEN_1819 = 11'h71b == WADDR ? 11'h71b : _GEN_1818; // @[RAM_ST.scala 31:71]
  assign _GEN_1820 = 11'h71c == WADDR ? 11'h71c : _GEN_1819; // @[RAM_ST.scala 31:71]
  assign _GEN_1821 = 11'h71d == WADDR ? 11'h71d : _GEN_1820; // @[RAM_ST.scala 31:71]
  assign _GEN_1822 = 11'h71e == WADDR ? 11'h71e : _GEN_1821; // @[RAM_ST.scala 31:71]
  assign _GEN_1823 = 11'h71f == WADDR ? 11'h71f : _GEN_1822; // @[RAM_ST.scala 31:71]
  assign _GEN_1824 = 11'h720 == WADDR ? 11'h720 : _GEN_1823; // @[RAM_ST.scala 31:71]
  assign _GEN_1825 = 11'h721 == WADDR ? 11'h721 : _GEN_1824; // @[RAM_ST.scala 31:71]
  assign _GEN_1826 = 11'h722 == WADDR ? 11'h722 : _GEN_1825; // @[RAM_ST.scala 31:71]
  assign _GEN_1827 = 11'h723 == WADDR ? 11'h723 : _GEN_1826; // @[RAM_ST.scala 31:71]
  assign _GEN_1828 = 11'h724 == WADDR ? 11'h724 : _GEN_1827; // @[RAM_ST.scala 31:71]
  assign _GEN_1829 = 11'h725 == WADDR ? 11'h725 : _GEN_1828; // @[RAM_ST.scala 31:71]
  assign _GEN_1830 = 11'h726 == WADDR ? 11'h726 : _GEN_1829; // @[RAM_ST.scala 31:71]
  assign _GEN_1831 = 11'h727 == WADDR ? 11'h727 : _GEN_1830; // @[RAM_ST.scala 31:71]
  assign _GEN_1832 = 11'h728 == WADDR ? 11'h728 : _GEN_1831; // @[RAM_ST.scala 31:71]
  assign _GEN_1833 = 11'h729 == WADDR ? 11'h729 : _GEN_1832; // @[RAM_ST.scala 31:71]
  assign _GEN_1834 = 11'h72a == WADDR ? 11'h72a : _GEN_1833; // @[RAM_ST.scala 31:71]
  assign _GEN_1835 = 11'h72b == WADDR ? 11'h72b : _GEN_1834; // @[RAM_ST.scala 31:71]
  assign _GEN_1836 = 11'h72c == WADDR ? 11'h72c : _GEN_1835; // @[RAM_ST.scala 31:71]
  assign _GEN_1837 = 11'h72d == WADDR ? 11'h72d : _GEN_1836; // @[RAM_ST.scala 31:71]
  assign _GEN_1838 = 11'h72e == WADDR ? 11'h72e : _GEN_1837; // @[RAM_ST.scala 31:71]
  assign _GEN_1839 = 11'h72f == WADDR ? 11'h72f : _GEN_1838; // @[RAM_ST.scala 31:71]
  assign _GEN_1840 = 11'h730 == WADDR ? 11'h730 : _GEN_1839; // @[RAM_ST.scala 31:71]
  assign _GEN_1841 = 11'h731 == WADDR ? 11'h731 : _GEN_1840; // @[RAM_ST.scala 31:71]
  assign _GEN_1842 = 11'h732 == WADDR ? 11'h732 : _GEN_1841; // @[RAM_ST.scala 31:71]
  assign _GEN_1843 = 11'h733 == WADDR ? 11'h733 : _GEN_1842; // @[RAM_ST.scala 31:71]
  assign _GEN_1844 = 11'h734 == WADDR ? 11'h734 : _GEN_1843; // @[RAM_ST.scala 31:71]
  assign _GEN_1845 = 11'h735 == WADDR ? 11'h735 : _GEN_1844; // @[RAM_ST.scala 31:71]
  assign _GEN_1846 = 11'h736 == WADDR ? 11'h736 : _GEN_1845; // @[RAM_ST.scala 31:71]
  assign _GEN_1847 = 11'h737 == WADDR ? 11'h737 : _GEN_1846; // @[RAM_ST.scala 31:71]
  assign _GEN_1848 = 11'h738 == WADDR ? 11'h738 : _GEN_1847; // @[RAM_ST.scala 31:71]
  assign _GEN_1849 = 11'h739 == WADDR ? 11'h739 : _GEN_1848; // @[RAM_ST.scala 31:71]
  assign _GEN_1850 = 11'h73a == WADDR ? 11'h73a : _GEN_1849; // @[RAM_ST.scala 31:71]
  assign _GEN_1851 = 11'h73b == WADDR ? 11'h73b : _GEN_1850; // @[RAM_ST.scala 31:71]
  assign _GEN_1852 = 11'h73c == WADDR ? 11'h73c : _GEN_1851; // @[RAM_ST.scala 31:71]
  assign _GEN_1853 = 11'h73d == WADDR ? 11'h73d : _GEN_1852; // @[RAM_ST.scala 31:71]
  assign _GEN_1854 = 11'h73e == WADDR ? 11'h73e : _GEN_1853; // @[RAM_ST.scala 31:71]
  assign _GEN_1855 = 11'h73f == WADDR ? 11'h73f : _GEN_1854; // @[RAM_ST.scala 31:71]
  assign _GEN_1856 = 11'h740 == WADDR ? 11'h740 : _GEN_1855; // @[RAM_ST.scala 31:71]
  assign _GEN_1857 = 11'h741 == WADDR ? 11'h741 : _GEN_1856; // @[RAM_ST.scala 31:71]
  assign _GEN_1858 = 11'h742 == WADDR ? 11'h742 : _GEN_1857; // @[RAM_ST.scala 31:71]
  assign _GEN_1859 = 11'h743 == WADDR ? 11'h743 : _GEN_1858; // @[RAM_ST.scala 31:71]
  assign _GEN_1860 = 11'h744 == WADDR ? 11'h744 : _GEN_1859; // @[RAM_ST.scala 31:71]
  assign _GEN_1861 = 11'h745 == WADDR ? 11'h745 : _GEN_1860; // @[RAM_ST.scala 31:71]
  assign _GEN_1862 = 11'h746 == WADDR ? 11'h746 : _GEN_1861; // @[RAM_ST.scala 31:71]
  assign _GEN_1863 = 11'h747 == WADDR ? 11'h747 : _GEN_1862; // @[RAM_ST.scala 31:71]
  assign _GEN_1864 = 11'h748 == WADDR ? 11'h748 : _GEN_1863; // @[RAM_ST.scala 31:71]
  assign _GEN_1865 = 11'h749 == WADDR ? 11'h749 : _GEN_1864; // @[RAM_ST.scala 31:71]
  assign _GEN_1866 = 11'h74a == WADDR ? 11'h74a : _GEN_1865; // @[RAM_ST.scala 31:71]
  assign _GEN_1867 = 11'h74b == WADDR ? 11'h74b : _GEN_1866; // @[RAM_ST.scala 31:71]
  assign _GEN_1868 = 11'h74c == WADDR ? 11'h74c : _GEN_1867; // @[RAM_ST.scala 31:71]
  assign _GEN_1869 = 11'h74d == WADDR ? 11'h74d : _GEN_1868; // @[RAM_ST.scala 31:71]
  assign _GEN_1870 = 11'h74e == WADDR ? 11'h74e : _GEN_1869; // @[RAM_ST.scala 31:71]
  assign _GEN_1871 = 11'h74f == WADDR ? 11'h74f : _GEN_1870; // @[RAM_ST.scala 31:71]
  assign _GEN_1872 = 11'h750 == WADDR ? 11'h750 : _GEN_1871; // @[RAM_ST.scala 31:71]
  assign _GEN_1873 = 11'h751 == WADDR ? 11'h751 : _GEN_1872; // @[RAM_ST.scala 31:71]
  assign _GEN_1874 = 11'h752 == WADDR ? 11'h752 : _GEN_1873; // @[RAM_ST.scala 31:71]
  assign _GEN_1875 = 11'h753 == WADDR ? 11'h753 : _GEN_1874; // @[RAM_ST.scala 31:71]
  assign _GEN_1876 = 11'h754 == WADDR ? 11'h754 : _GEN_1875; // @[RAM_ST.scala 31:71]
  assign _GEN_1877 = 11'h755 == WADDR ? 11'h755 : _GEN_1876; // @[RAM_ST.scala 31:71]
  assign _GEN_1878 = 11'h756 == WADDR ? 11'h756 : _GEN_1877; // @[RAM_ST.scala 31:71]
  assign _GEN_1879 = 11'h757 == WADDR ? 11'h757 : _GEN_1878; // @[RAM_ST.scala 31:71]
  assign _GEN_1880 = 11'h758 == WADDR ? 11'h758 : _GEN_1879; // @[RAM_ST.scala 31:71]
  assign _GEN_1881 = 11'h759 == WADDR ? 11'h759 : _GEN_1880; // @[RAM_ST.scala 31:71]
  assign _GEN_1882 = 11'h75a == WADDR ? 11'h75a : _GEN_1881; // @[RAM_ST.scala 31:71]
  assign _GEN_1883 = 11'h75b == WADDR ? 11'h75b : _GEN_1882; // @[RAM_ST.scala 31:71]
  assign _GEN_1884 = 11'h75c == WADDR ? 11'h75c : _GEN_1883; // @[RAM_ST.scala 31:71]
  assign _GEN_1885 = 11'h75d == WADDR ? 11'h75d : _GEN_1884; // @[RAM_ST.scala 31:71]
  assign _GEN_1886 = 11'h75e == WADDR ? 11'h75e : _GEN_1885; // @[RAM_ST.scala 31:71]
  assign _GEN_1887 = 11'h75f == WADDR ? 11'h75f : _GEN_1886; // @[RAM_ST.scala 31:71]
  assign _GEN_1888 = 11'h760 == WADDR ? 11'h760 : _GEN_1887; // @[RAM_ST.scala 31:71]
  assign _GEN_1889 = 11'h761 == WADDR ? 11'h761 : _GEN_1888; // @[RAM_ST.scala 31:71]
  assign _GEN_1890 = 11'h762 == WADDR ? 11'h762 : _GEN_1889; // @[RAM_ST.scala 31:71]
  assign _GEN_1891 = 11'h763 == WADDR ? 11'h763 : _GEN_1890; // @[RAM_ST.scala 31:71]
  assign _GEN_1892 = 11'h764 == WADDR ? 11'h764 : _GEN_1891; // @[RAM_ST.scala 31:71]
  assign _GEN_1893 = 11'h765 == WADDR ? 11'h765 : _GEN_1892; // @[RAM_ST.scala 31:71]
  assign _GEN_1894 = 11'h766 == WADDR ? 11'h766 : _GEN_1893; // @[RAM_ST.scala 31:71]
  assign _GEN_1895 = 11'h767 == WADDR ? 11'h767 : _GEN_1894; // @[RAM_ST.scala 31:71]
  assign _GEN_1896 = 11'h768 == WADDR ? 11'h768 : _GEN_1895; // @[RAM_ST.scala 31:71]
  assign _GEN_1897 = 11'h769 == WADDR ? 11'h769 : _GEN_1896; // @[RAM_ST.scala 31:71]
  assign _GEN_1898 = 11'h76a == WADDR ? 11'h76a : _GEN_1897; // @[RAM_ST.scala 31:71]
  assign _GEN_1899 = 11'h76b == WADDR ? 11'h76b : _GEN_1898; // @[RAM_ST.scala 31:71]
  assign _GEN_1900 = 11'h76c == WADDR ? 11'h76c : _GEN_1899; // @[RAM_ST.scala 31:71]
  assign _GEN_1901 = 11'h76d == WADDR ? 11'h76d : _GEN_1900; // @[RAM_ST.scala 31:71]
  assign _GEN_1902 = 11'h76e == WADDR ? 11'h76e : _GEN_1901; // @[RAM_ST.scala 31:71]
  assign _GEN_1903 = 11'h76f == WADDR ? 11'h76f : _GEN_1902; // @[RAM_ST.scala 31:71]
  assign _GEN_1904 = 11'h770 == WADDR ? 11'h770 : _GEN_1903; // @[RAM_ST.scala 31:71]
  assign _GEN_1905 = 11'h771 == WADDR ? 11'h771 : _GEN_1904; // @[RAM_ST.scala 31:71]
  assign _GEN_1906 = 11'h772 == WADDR ? 11'h772 : _GEN_1905; // @[RAM_ST.scala 31:71]
  assign _GEN_1907 = 11'h773 == WADDR ? 11'h773 : _GEN_1906; // @[RAM_ST.scala 31:71]
  assign _GEN_1908 = 11'h774 == WADDR ? 11'h774 : _GEN_1907; // @[RAM_ST.scala 31:71]
  assign _GEN_1909 = 11'h775 == WADDR ? 11'h775 : _GEN_1908; // @[RAM_ST.scala 31:71]
  assign _GEN_1910 = 11'h776 == WADDR ? 11'h776 : _GEN_1909; // @[RAM_ST.scala 31:71]
  assign _GEN_1911 = 11'h777 == WADDR ? 11'h777 : _GEN_1910; // @[RAM_ST.scala 31:71]
  assign _GEN_1912 = 11'h778 == WADDR ? 11'h778 : _GEN_1911; // @[RAM_ST.scala 31:71]
  assign _GEN_1913 = 11'h779 == WADDR ? 11'h779 : _GEN_1912; // @[RAM_ST.scala 31:71]
  assign _GEN_1914 = 11'h77a == WADDR ? 11'h77a : _GEN_1913; // @[RAM_ST.scala 31:71]
  assign _GEN_1915 = 11'h77b == WADDR ? 11'h77b : _GEN_1914; // @[RAM_ST.scala 31:71]
  assign _GEN_1916 = 11'h77c == WADDR ? 11'h77c : _GEN_1915; // @[RAM_ST.scala 31:71]
  assign _GEN_1917 = 11'h77d == WADDR ? 11'h77d : _GEN_1916; // @[RAM_ST.scala 31:71]
  assign _GEN_1918 = 11'h77e == WADDR ? 11'h77e : _GEN_1917; // @[RAM_ST.scala 31:71]
  assign _GEN_1919 = 11'h77f == WADDR ? 11'h77f : _GEN_1918; // @[RAM_ST.scala 31:71]
  assign _T = {{1'd0}, _GEN_1919}; // @[RAM_ST.scala 31:71]
  assign _GEN_1926 = 11'h1 == RADDR ? 11'h1 : 11'h0; // @[RAM_ST.scala 32:46]
  assign _GEN_1927 = 11'h2 == RADDR ? 11'h2 : _GEN_1926; // @[RAM_ST.scala 32:46]
  assign _GEN_1928 = 11'h3 == RADDR ? 11'h3 : _GEN_1927; // @[RAM_ST.scala 32:46]
  assign _GEN_1929 = 11'h4 == RADDR ? 11'h4 : _GEN_1928; // @[RAM_ST.scala 32:46]
  assign _GEN_1930 = 11'h5 == RADDR ? 11'h5 : _GEN_1929; // @[RAM_ST.scala 32:46]
  assign _GEN_1931 = 11'h6 == RADDR ? 11'h6 : _GEN_1930; // @[RAM_ST.scala 32:46]
  assign _GEN_1932 = 11'h7 == RADDR ? 11'h7 : _GEN_1931; // @[RAM_ST.scala 32:46]
  assign _GEN_1933 = 11'h8 == RADDR ? 11'h8 : _GEN_1932; // @[RAM_ST.scala 32:46]
  assign _GEN_1934 = 11'h9 == RADDR ? 11'h9 : _GEN_1933; // @[RAM_ST.scala 32:46]
  assign _GEN_1935 = 11'ha == RADDR ? 11'ha : _GEN_1934; // @[RAM_ST.scala 32:46]
  assign _GEN_1936 = 11'hb == RADDR ? 11'hb : _GEN_1935; // @[RAM_ST.scala 32:46]
  assign _GEN_1937 = 11'hc == RADDR ? 11'hc : _GEN_1936; // @[RAM_ST.scala 32:46]
  assign _GEN_1938 = 11'hd == RADDR ? 11'hd : _GEN_1937; // @[RAM_ST.scala 32:46]
  assign _GEN_1939 = 11'he == RADDR ? 11'he : _GEN_1938; // @[RAM_ST.scala 32:46]
  assign _GEN_1940 = 11'hf == RADDR ? 11'hf : _GEN_1939; // @[RAM_ST.scala 32:46]
  assign _GEN_1941 = 11'h10 == RADDR ? 11'h10 : _GEN_1940; // @[RAM_ST.scala 32:46]
  assign _GEN_1942 = 11'h11 == RADDR ? 11'h11 : _GEN_1941; // @[RAM_ST.scala 32:46]
  assign _GEN_1943 = 11'h12 == RADDR ? 11'h12 : _GEN_1942; // @[RAM_ST.scala 32:46]
  assign _GEN_1944 = 11'h13 == RADDR ? 11'h13 : _GEN_1943; // @[RAM_ST.scala 32:46]
  assign _GEN_1945 = 11'h14 == RADDR ? 11'h14 : _GEN_1944; // @[RAM_ST.scala 32:46]
  assign _GEN_1946 = 11'h15 == RADDR ? 11'h15 : _GEN_1945; // @[RAM_ST.scala 32:46]
  assign _GEN_1947 = 11'h16 == RADDR ? 11'h16 : _GEN_1946; // @[RAM_ST.scala 32:46]
  assign _GEN_1948 = 11'h17 == RADDR ? 11'h17 : _GEN_1947; // @[RAM_ST.scala 32:46]
  assign _GEN_1949 = 11'h18 == RADDR ? 11'h18 : _GEN_1948; // @[RAM_ST.scala 32:46]
  assign _GEN_1950 = 11'h19 == RADDR ? 11'h19 : _GEN_1949; // @[RAM_ST.scala 32:46]
  assign _GEN_1951 = 11'h1a == RADDR ? 11'h1a : _GEN_1950; // @[RAM_ST.scala 32:46]
  assign _GEN_1952 = 11'h1b == RADDR ? 11'h1b : _GEN_1951; // @[RAM_ST.scala 32:46]
  assign _GEN_1953 = 11'h1c == RADDR ? 11'h1c : _GEN_1952; // @[RAM_ST.scala 32:46]
  assign _GEN_1954 = 11'h1d == RADDR ? 11'h1d : _GEN_1953; // @[RAM_ST.scala 32:46]
  assign _GEN_1955 = 11'h1e == RADDR ? 11'h1e : _GEN_1954; // @[RAM_ST.scala 32:46]
  assign _GEN_1956 = 11'h1f == RADDR ? 11'h1f : _GEN_1955; // @[RAM_ST.scala 32:46]
  assign _GEN_1957 = 11'h20 == RADDR ? 11'h20 : _GEN_1956; // @[RAM_ST.scala 32:46]
  assign _GEN_1958 = 11'h21 == RADDR ? 11'h21 : _GEN_1957; // @[RAM_ST.scala 32:46]
  assign _GEN_1959 = 11'h22 == RADDR ? 11'h22 : _GEN_1958; // @[RAM_ST.scala 32:46]
  assign _GEN_1960 = 11'h23 == RADDR ? 11'h23 : _GEN_1959; // @[RAM_ST.scala 32:46]
  assign _GEN_1961 = 11'h24 == RADDR ? 11'h24 : _GEN_1960; // @[RAM_ST.scala 32:46]
  assign _GEN_1962 = 11'h25 == RADDR ? 11'h25 : _GEN_1961; // @[RAM_ST.scala 32:46]
  assign _GEN_1963 = 11'h26 == RADDR ? 11'h26 : _GEN_1962; // @[RAM_ST.scala 32:46]
  assign _GEN_1964 = 11'h27 == RADDR ? 11'h27 : _GEN_1963; // @[RAM_ST.scala 32:46]
  assign _GEN_1965 = 11'h28 == RADDR ? 11'h28 : _GEN_1964; // @[RAM_ST.scala 32:46]
  assign _GEN_1966 = 11'h29 == RADDR ? 11'h29 : _GEN_1965; // @[RAM_ST.scala 32:46]
  assign _GEN_1967 = 11'h2a == RADDR ? 11'h2a : _GEN_1966; // @[RAM_ST.scala 32:46]
  assign _GEN_1968 = 11'h2b == RADDR ? 11'h2b : _GEN_1967; // @[RAM_ST.scala 32:46]
  assign _GEN_1969 = 11'h2c == RADDR ? 11'h2c : _GEN_1968; // @[RAM_ST.scala 32:46]
  assign _GEN_1970 = 11'h2d == RADDR ? 11'h2d : _GEN_1969; // @[RAM_ST.scala 32:46]
  assign _GEN_1971 = 11'h2e == RADDR ? 11'h2e : _GEN_1970; // @[RAM_ST.scala 32:46]
  assign _GEN_1972 = 11'h2f == RADDR ? 11'h2f : _GEN_1971; // @[RAM_ST.scala 32:46]
  assign _GEN_1973 = 11'h30 == RADDR ? 11'h30 : _GEN_1972; // @[RAM_ST.scala 32:46]
  assign _GEN_1974 = 11'h31 == RADDR ? 11'h31 : _GEN_1973; // @[RAM_ST.scala 32:46]
  assign _GEN_1975 = 11'h32 == RADDR ? 11'h32 : _GEN_1974; // @[RAM_ST.scala 32:46]
  assign _GEN_1976 = 11'h33 == RADDR ? 11'h33 : _GEN_1975; // @[RAM_ST.scala 32:46]
  assign _GEN_1977 = 11'h34 == RADDR ? 11'h34 : _GEN_1976; // @[RAM_ST.scala 32:46]
  assign _GEN_1978 = 11'h35 == RADDR ? 11'h35 : _GEN_1977; // @[RAM_ST.scala 32:46]
  assign _GEN_1979 = 11'h36 == RADDR ? 11'h36 : _GEN_1978; // @[RAM_ST.scala 32:46]
  assign _GEN_1980 = 11'h37 == RADDR ? 11'h37 : _GEN_1979; // @[RAM_ST.scala 32:46]
  assign _GEN_1981 = 11'h38 == RADDR ? 11'h38 : _GEN_1980; // @[RAM_ST.scala 32:46]
  assign _GEN_1982 = 11'h39 == RADDR ? 11'h39 : _GEN_1981; // @[RAM_ST.scala 32:46]
  assign _GEN_1983 = 11'h3a == RADDR ? 11'h3a : _GEN_1982; // @[RAM_ST.scala 32:46]
  assign _GEN_1984 = 11'h3b == RADDR ? 11'h3b : _GEN_1983; // @[RAM_ST.scala 32:46]
  assign _GEN_1985 = 11'h3c == RADDR ? 11'h3c : _GEN_1984; // @[RAM_ST.scala 32:46]
  assign _GEN_1986 = 11'h3d == RADDR ? 11'h3d : _GEN_1985; // @[RAM_ST.scala 32:46]
  assign _GEN_1987 = 11'h3e == RADDR ? 11'h3e : _GEN_1986; // @[RAM_ST.scala 32:46]
  assign _GEN_1988 = 11'h3f == RADDR ? 11'h3f : _GEN_1987; // @[RAM_ST.scala 32:46]
  assign _GEN_1989 = 11'h40 == RADDR ? 11'h40 : _GEN_1988; // @[RAM_ST.scala 32:46]
  assign _GEN_1990 = 11'h41 == RADDR ? 11'h41 : _GEN_1989; // @[RAM_ST.scala 32:46]
  assign _GEN_1991 = 11'h42 == RADDR ? 11'h42 : _GEN_1990; // @[RAM_ST.scala 32:46]
  assign _GEN_1992 = 11'h43 == RADDR ? 11'h43 : _GEN_1991; // @[RAM_ST.scala 32:46]
  assign _GEN_1993 = 11'h44 == RADDR ? 11'h44 : _GEN_1992; // @[RAM_ST.scala 32:46]
  assign _GEN_1994 = 11'h45 == RADDR ? 11'h45 : _GEN_1993; // @[RAM_ST.scala 32:46]
  assign _GEN_1995 = 11'h46 == RADDR ? 11'h46 : _GEN_1994; // @[RAM_ST.scala 32:46]
  assign _GEN_1996 = 11'h47 == RADDR ? 11'h47 : _GEN_1995; // @[RAM_ST.scala 32:46]
  assign _GEN_1997 = 11'h48 == RADDR ? 11'h48 : _GEN_1996; // @[RAM_ST.scala 32:46]
  assign _GEN_1998 = 11'h49 == RADDR ? 11'h49 : _GEN_1997; // @[RAM_ST.scala 32:46]
  assign _GEN_1999 = 11'h4a == RADDR ? 11'h4a : _GEN_1998; // @[RAM_ST.scala 32:46]
  assign _GEN_2000 = 11'h4b == RADDR ? 11'h4b : _GEN_1999; // @[RAM_ST.scala 32:46]
  assign _GEN_2001 = 11'h4c == RADDR ? 11'h4c : _GEN_2000; // @[RAM_ST.scala 32:46]
  assign _GEN_2002 = 11'h4d == RADDR ? 11'h4d : _GEN_2001; // @[RAM_ST.scala 32:46]
  assign _GEN_2003 = 11'h4e == RADDR ? 11'h4e : _GEN_2002; // @[RAM_ST.scala 32:46]
  assign _GEN_2004 = 11'h4f == RADDR ? 11'h4f : _GEN_2003; // @[RAM_ST.scala 32:46]
  assign _GEN_2005 = 11'h50 == RADDR ? 11'h50 : _GEN_2004; // @[RAM_ST.scala 32:46]
  assign _GEN_2006 = 11'h51 == RADDR ? 11'h51 : _GEN_2005; // @[RAM_ST.scala 32:46]
  assign _GEN_2007 = 11'h52 == RADDR ? 11'h52 : _GEN_2006; // @[RAM_ST.scala 32:46]
  assign _GEN_2008 = 11'h53 == RADDR ? 11'h53 : _GEN_2007; // @[RAM_ST.scala 32:46]
  assign _GEN_2009 = 11'h54 == RADDR ? 11'h54 : _GEN_2008; // @[RAM_ST.scala 32:46]
  assign _GEN_2010 = 11'h55 == RADDR ? 11'h55 : _GEN_2009; // @[RAM_ST.scala 32:46]
  assign _GEN_2011 = 11'h56 == RADDR ? 11'h56 : _GEN_2010; // @[RAM_ST.scala 32:46]
  assign _GEN_2012 = 11'h57 == RADDR ? 11'h57 : _GEN_2011; // @[RAM_ST.scala 32:46]
  assign _GEN_2013 = 11'h58 == RADDR ? 11'h58 : _GEN_2012; // @[RAM_ST.scala 32:46]
  assign _GEN_2014 = 11'h59 == RADDR ? 11'h59 : _GEN_2013; // @[RAM_ST.scala 32:46]
  assign _GEN_2015 = 11'h5a == RADDR ? 11'h5a : _GEN_2014; // @[RAM_ST.scala 32:46]
  assign _GEN_2016 = 11'h5b == RADDR ? 11'h5b : _GEN_2015; // @[RAM_ST.scala 32:46]
  assign _GEN_2017 = 11'h5c == RADDR ? 11'h5c : _GEN_2016; // @[RAM_ST.scala 32:46]
  assign _GEN_2018 = 11'h5d == RADDR ? 11'h5d : _GEN_2017; // @[RAM_ST.scala 32:46]
  assign _GEN_2019 = 11'h5e == RADDR ? 11'h5e : _GEN_2018; // @[RAM_ST.scala 32:46]
  assign _GEN_2020 = 11'h5f == RADDR ? 11'h5f : _GEN_2019; // @[RAM_ST.scala 32:46]
  assign _GEN_2021 = 11'h60 == RADDR ? 11'h60 : _GEN_2020; // @[RAM_ST.scala 32:46]
  assign _GEN_2022 = 11'h61 == RADDR ? 11'h61 : _GEN_2021; // @[RAM_ST.scala 32:46]
  assign _GEN_2023 = 11'h62 == RADDR ? 11'h62 : _GEN_2022; // @[RAM_ST.scala 32:46]
  assign _GEN_2024 = 11'h63 == RADDR ? 11'h63 : _GEN_2023; // @[RAM_ST.scala 32:46]
  assign _GEN_2025 = 11'h64 == RADDR ? 11'h64 : _GEN_2024; // @[RAM_ST.scala 32:46]
  assign _GEN_2026 = 11'h65 == RADDR ? 11'h65 : _GEN_2025; // @[RAM_ST.scala 32:46]
  assign _GEN_2027 = 11'h66 == RADDR ? 11'h66 : _GEN_2026; // @[RAM_ST.scala 32:46]
  assign _GEN_2028 = 11'h67 == RADDR ? 11'h67 : _GEN_2027; // @[RAM_ST.scala 32:46]
  assign _GEN_2029 = 11'h68 == RADDR ? 11'h68 : _GEN_2028; // @[RAM_ST.scala 32:46]
  assign _GEN_2030 = 11'h69 == RADDR ? 11'h69 : _GEN_2029; // @[RAM_ST.scala 32:46]
  assign _GEN_2031 = 11'h6a == RADDR ? 11'h6a : _GEN_2030; // @[RAM_ST.scala 32:46]
  assign _GEN_2032 = 11'h6b == RADDR ? 11'h6b : _GEN_2031; // @[RAM_ST.scala 32:46]
  assign _GEN_2033 = 11'h6c == RADDR ? 11'h6c : _GEN_2032; // @[RAM_ST.scala 32:46]
  assign _GEN_2034 = 11'h6d == RADDR ? 11'h6d : _GEN_2033; // @[RAM_ST.scala 32:46]
  assign _GEN_2035 = 11'h6e == RADDR ? 11'h6e : _GEN_2034; // @[RAM_ST.scala 32:46]
  assign _GEN_2036 = 11'h6f == RADDR ? 11'h6f : _GEN_2035; // @[RAM_ST.scala 32:46]
  assign _GEN_2037 = 11'h70 == RADDR ? 11'h70 : _GEN_2036; // @[RAM_ST.scala 32:46]
  assign _GEN_2038 = 11'h71 == RADDR ? 11'h71 : _GEN_2037; // @[RAM_ST.scala 32:46]
  assign _GEN_2039 = 11'h72 == RADDR ? 11'h72 : _GEN_2038; // @[RAM_ST.scala 32:46]
  assign _GEN_2040 = 11'h73 == RADDR ? 11'h73 : _GEN_2039; // @[RAM_ST.scala 32:46]
  assign _GEN_2041 = 11'h74 == RADDR ? 11'h74 : _GEN_2040; // @[RAM_ST.scala 32:46]
  assign _GEN_2042 = 11'h75 == RADDR ? 11'h75 : _GEN_2041; // @[RAM_ST.scala 32:46]
  assign _GEN_2043 = 11'h76 == RADDR ? 11'h76 : _GEN_2042; // @[RAM_ST.scala 32:46]
  assign _GEN_2044 = 11'h77 == RADDR ? 11'h77 : _GEN_2043; // @[RAM_ST.scala 32:46]
  assign _GEN_2045 = 11'h78 == RADDR ? 11'h78 : _GEN_2044; // @[RAM_ST.scala 32:46]
  assign _GEN_2046 = 11'h79 == RADDR ? 11'h79 : _GEN_2045; // @[RAM_ST.scala 32:46]
  assign _GEN_2047 = 11'h7a == RADDR ? 11'h7a : _GEN_2046; // @[RAM_ST.scala 32:46]
  assign _GEN_2048 = 11'h7b == RADDR ? 11'h7b : _GEN_2047; // @[RAM_ST.scala 32:46]
  assign _GEN_2049 = 11'h7c == RADDR ? 11'h7c : _GEN_2048; // @[RAM_ST.scala 32:46]
  assign _GEN_2050 = 11'h7d == RADDR ? 11'h7d : _GEN_2049; // @[RAM_ST.scala 32:46]
  assign _GEN_2051 = 11'h7e == RADDR ? 11'h7e : _GEN_2050; // @[RAM_ST.scala 32:46]
  assign _GEN_2052 = 11'h7f == RADDR ? 11'h7f : _GEN_2051; // @[RAM_ST.scala 32:46]
  assign _GEN_2053 = 11'h80 == RADDR ? 11'h80 : _GEN_2052; // @[RAM_ST.scala 32:46]
  assign _GEN_2054 = 11'h81 == RADDR ? 11'h81 : _GEN_2053; // @[RAM_ST.scala 32:46]
  assign _GEN_2055 = 11'h82 == RADDR ? 11'h82 : _GEN_2054; // @[RAM_ST.scala 32:46]
  assign _GEN_2056 = 11'h83 == RADDR ? 11'h83 : _GEN_2055; // @[RAM_ST.scala 32:46]
  assign _GEN_2057 = 11'h84 == RADDR ? 11'h84 : _GEN_2056; // @[RAM_ST.scala 32:46]
  assign _GEN_2058 = 11'h85 == RADDR ? 11'h85 : _GEN_2057; // @[RAM_ST.scala 32:46]
  assign _GEN_2059 = 11'h86 == RADDR ? 11'h86 : _GEN_2058; // @[RAM_ST.scala 32:46]
  assign _GEN_2060 = 11'h87 == RADDR ? 11'h87 : _GEN_2059; // @[RAM_ST.scala 32:46]
  assign _GEN_2061 = 11'h88 == RADDR ? 11'h88 : _GEN_2060; // @[RAM_ST.scala 32:46]
  assign _GEN_2062 = 11'h89 == RADDR ? 11'h89 : _GEN_2061; // @[RAM_ST.scala 32:46]
  assign _GEN_2063 = 11'h8a == RADDR ? 11'h8a : _GEN_2062; // @[RAM_ST.scala 32:46]
  assign _GEN_2064 = 11'h8b == RADDR ? 11'h8b : _GEN_2063; // @[RAM_ST.scala 32:46]
  assign _GEN_2065 = 11'h8c == RADDR ? 11'h8c : _GEN_2064; // @[RAM_ST.scala 32:46]
  assign _GEN_2066 = 11'h8d == RADDR ? 11'h8d : _GEN_2065; // @[RAM_ST.scala 32:46]
  assign _GEN_2067 = 11'h8e == RADDR ? 11'h8e : _GEN_2066; // @[RAM_ST.scala 32:46]
  assign _GEN_2068 = 11'h8f == RADDR ? 11'h8f : _GEN_2067; // @[RAM_ST.scala 32:46]
  assign _GEN_2069 = 11'h90 == RADDR ? 11'h90 : _GEN_2068; // @[RAM_ST.scala 32:46]
  assign _GEN_2070 = 11'h91 == RADDR ? 11'h91 : _GEN_2069; // @[RAM_ST.scala 32:46]
  assign _GEN_2071 = 11'h92 == RADDR ? 11'h92 : _GEN_2070; // @[RAM_ST.scala 32:46]
  assign _GEN_2072 = 11'h93 == RADDR ? 11'h93 : _GEN_2071; // @[RAM_ST.scala 32:46]
  assign _GEN_2073 = 11'h94 == RADDR ? 11'h94 : _GEN_2072; // @[RAM_ST.scala 32:46]
  assign _GEN_2074 = 11'h95 == RADDR ? 11'h95 : _GEN_2073; // @[RAM_ST.scala 32:46]
  assign _GEN_2075 = 11'h96 == RADDR ? 11'h96 : _GEN_2074; // @[RAM_ST.scala 32:46]
  assign _GEN_2076 = 11'h97 == RADDR ? 11'h97 : _GEN_2075; // @[RAM_ST.scala 32:46]
  assign _GEN_2077 = 11'h98 == RADDR ? 11'h98 : _GEN_2076; // @[RAM_ST.scala 32:46]
  assign _GEN_2078 = 11'h99 == RADDR ? 11'h99 : _GEN_2077; // @[RAM_ST.scala 32:46]
  assign _GEN_2079 = 11'h9a == RADDR ? 11'h9a : _GEN_2078; // @[RAM_ST.scala 32:46]
  assign _GEN_2080 = 11'h9b == RADDR ? 11'h9b : _GEN_2079; // @[RAM_ST.scala 32:46]
  assign _GEN_2081 = 11'h9c == RADDR ? 11'h9c : _GEN_2080; // @[RAM_ST.scala 32:46]
  assign _GEN_2082 = 11'h9d == RADDR ? 11'h9d : _GEN_2081; // @[RAM_ST.scala 32:46]
  assign _GEN_2083 = 11'h9e == RADDR ? 11'h9e : _GEN_2082; // @[RAM_ST.scala 32:46]
  assign _GEN_2084 = 11'h9f == RADDR ? 11'h9f : _GEN_2083; // @[RAM_ST.scala 32:46]
  assign _GEN_2085 = 11'ha0 == RADDR ? 11'ha0 : _GEN_2084; // @[RAM_ST.scala 32:46]
  assign _GEN_2086 = 11'ha1 == RADDR ? 11'ha1 : _GEN_2085; // @[RAM_ST.scala 32:46]
  assign _GEN_2087 = 11'ha2 == RADDR ? 11'ha2 : _GEN_2086; // @[RAM_ST.scala 32:46]
  assign _GEN_2088 = 11'ha3 == RADDR ? 11'ha3 : _GEN_2087; // @[RAM_ST.scala 32:46]
  assign _GEN_2089 = 11'ha4 == RADDR ? 11'ha4 : _GEN_2088; // @[RAM_ST.scala 32:46]
  assign _GEN_2090 = 11'ha5 == RADDR ? 11'ha5 : _GEN_2089; // @[RAM_ST.scala 32:46]
  assign _GEN_2091 = 11'ha6 == RADDR ? 11'ha6 : _GEN_2090; // @[RAM_ST.scala 32:46]
  assign _GEN_2092 = 11'ha7 == RADDR ? 11'ha7 : _GEN_2091; // @[RAM_ST.scala 32:46]
  assign _GEN_2093 = 11'ha8 == RADDR ? 11'ha8 : _GEN_2092; // @[RAM_ST.scala 32:46]
  assign _GEN_2094 = 11'ha9 == RADDR ? 11'ha9 : _GEN_2093; // @[RAM_ST.scala 32:46]
  assign _GEN_2095 = 11'haa == RADDR ? 11'haa : _GEN_2094; // @[RAM_ST.scala 32:46]
  assign _GEN_2096 = 11'hab == RADDR ? 11'hab : _GEN_2095; // @[RAM_ST.scala 32:46]
  assign _GEN_2097 = 11'hac == RADDR ? 11'hac : _GEN_2096; // @[RAM_ST.scala 32:46]
  assign _GEN_2098 = 11'had == RADDR ? 11'had : _GEN_2097; // @[RAM_ST.scala 32:46]
  assign _GEN_2099 = 11'hae == RADDR ? 11'hae : _GEN_2098; // @[RAM_ST.scala 32:46]
  assign _GEN_2100 = 11'haf == RADDR ? 11'haf : _GEN_2099; // @[RAM_ST.scala 32:46]
  assign _GEN_2101 = 11'hb0 == RADDR ? 11'hb0 : _GEN_2100; // @[RAM_ST.scala 32:46]
  assign _GEN_2102 = 11'hb1 == RADDR ? 11'hb1 : _GEN_2101; // @[RAM_ST.scala 32:46]
  assign _GEN_2103 = 11'hb2 == RADDR ? 11'hb2 : _GEN_2102; // @[RAM_ST.scala 32:46]
  assign _GEN_2104 = 11'hb3 == RADDR ? 11'hb3 : _GEN_2103; // @[RAM_ST.scala 32:46]
  assign _GEN_2105 = 11'hb4 == RADDR ? 11'hb4 : _GEN_2104; // @[RAM_ST.scala 32:46]
  assign _GEN_2106 = 11'hb5 == RADDR ? 11'hb5 : _GEN_2105; // @[RAM_ST.scala 32:46]
  assign _GEN_2107 = 11'hb6 == RADDR ? 11'hb6 : _GEN_2106; // @[RAM_ST.scala 32:46]
  assign _GEN_2108 = 11'hb7 == RADDR ? 11'hb7 : _GEN_2107; // @[RAM_ST.scala 32:46]
  assign _GEN_2109 = 11'hb8 == RADDR ? 11'hb8 : _GEN_2108; // @[RAM_ST.scala 32:46]
  assign _GEN_2110 = 11'hb9 == RADDR ? 11'hb9 : _GEN_2109; // @[RAM_ST.scala 32:46]
  assign _GEN_2111 = 11'hba == RADDR ? 11'hba : _GEN_2110; // @[RAM_ST.scala 32:46]
  assign _GEN_2112 = 11'hbb == RADDR ? 11'hbb : _GEN_2111; // @[RAM_ST.scala 32:46]
  assign _GEN_2113 = 11'hbc == RADDR ? 11'hbc : _GEN_2112; // @[RAM_ST.scala 32:46]
  assign _GEN_2114 = 11'hbd == RADDR ? 11'hbd : _GEN_2113; // @[RAM_ST.scala 32:46]
  assign _GEN_2115 = 11'hbe == RADDR ? 11'hbe : _GEN_2114; // @[RAM_ST.scala 32:46]
  assign _GEN_2116 = 11'hbf == RADDR ? 11'hbf : _GEN_2115; // @[RAM_ST.scala 32:46]
  assign _GEN_2117 = 11'hc0 == RADDR ? 11'hc0 : _GEN_2116; // @[RAM_ST.scala 32:46]
  assign _GEN_2118 = 11'hc1 == RADDR ? 11'hc1 : _GEN_2117; // @[RAM_ST.scala 32:46]
  assign _GEN_2119 = 11'hc2 == RADDR ? 11'hc2 : _GEN_2118; // @[RAM_ST.scala 32:46]
  assign _GEN_2120 = 11'hc3 == RADDR ? 11'hc3 : _GEN_2119; // @[RAM_ST.scala 32:46]
  assign _GEN_2121 = 11'hc4 == RADDR ? 11'hc4 : _GEN_2120; // @[RAM_ST.scala 32:46]
  assign _GEN_2122 = 11'hc5 == RADDR ? 11'hc5 : _GEN_2121; // @[RAM_ST.scala 32:46]
  assign _GEN_2123 = 11'hc6 == RADDR ? 11'hc6 : _GEN_2122; // @[RAM_ST.scala 32:46]
  assign _GEN_2124 = 11'hc7 == RADDR ? 11'hc7 : _GEN_2123; // @[RAM_ST.scala 32:46]
  assign _GEN_2125 = 11'hc8 == RADDR ? 11'hc8 : _GEN_2124; // @[RAM_ST.scala 32:46]
  assign _GEN_2126 = 11'hc9 == RADDR ? 11'hc9 : _GEN_2125; // @[RAM_ST.scala 32:46]
  assign _GEN_2127 = 11'hca == RADDR ? 11'hca : _GEN_2126; // @[RAM_ST.scala 32:46]
  assign _GEN_2128 = 11'hcb == RADDR ? 11'hcb : _GEN_2127; // @[RAM_ST.scala 32:46]
  assign _GEN_2129 = 11'hcc == RADDR ? 11'hcc : _GEN_2128; // @[RAM_ST.scala 32:46]
  assign _GEN_2130 = 11'hcd == RADDR ? 11'hcd : _GEN_2129; // @[RAM_ST.scala 32:46]
  assign _GEN_2131 = 11'hce == RADDR ? 11'hce : _GEN_2130; // @[RAM_ST.scala 32:46]
  assign _GEN_2132 = 11'hcf == RADDR ? 11'hcf : _GEN_2131; // @[RAM_ST.scala 32:46]
  assign _GEN_2133 = 11'hd0 == RADDR ? 11'hd0 : _GEN_2132; // @[RAM_ST.scala 32:46]
  assign _GEN_2134 = 11'hd1 == RADDR ? 11'hd1 : _GEN_2133; // @[RAM_ST.scala 32:46]
  assign _GEN_2135 = 11'hd2 == RADDR ? 11'hd2 : _GEN_2134; // @[RAM_ST.scala 32:46]
  assign _GEN_2136 = 11'hd3 == RADDR ? 11'hd3 : _GEN_2135; // @[RAM_ST.scala 32:46]
  assign _GEN_2137 = 11'hd4 == RADDR ? 11'hd4 : _GEN_2136; // @[RAM_ST.scala 32:46]
  assign _GEN_2138 = 11'hd5 == RADDR ? 11'hd5 : _GEN_2137; // @[RAM_ST.scala 32:46]
  assign _GEN_2139 = 11'hd6 == RADDR ? 11'hd6 : _GEN_2138; // @[RAM_ST.scala 32:46]
  assign _GEN_2140 = 11'hd7 == RADDR ? 11'hd7 : _GEN_2139; // @[RAM_ST.scala 32:46]
  assign _GEN_2141 = 11'hd8 == RADDR ? 11'hd8 : _GEN_2140; // @[RAM_ST.scala 32:46]
  assign _GEN_2142 = 11'hd9 == RADDR ? 11'hd9 : _GEN_2141; // @[RAM_ST.scala 32:46]
  assign _GEN_2143 = 11'hda == RADDR ? 11'hda : _GEN_2142; // @[RAM_ST.scala 32:46]
  assign _GEN_2144 = 11'hdb == RADDR ? 11'hdb : _GEN_2143; // @[RAM_ST.scala 32:46]
  assign _GEN_2145 = 11'hdc == RADDR ? 11'hdc : _GEN_2144; // @[RAM_ST.scala 32:46]
  assign _GEN_2146 = 11'hdd == RADDR ? 11'hdd : _GEN_2145; // @[RAM_ST.scala 32:46]
  assign _GEN_2147 = 11'hde == RADDR ? 11'hde : _GEN_2146; // @[RAM_ST.scala 32:46]
  assign _GEN_2148 = 11'hdf == RADDR ? 11'hdf : _GEN_2147; // @[RAM_ST.scala 32:46]
  assign _GEN_2149 = 11'he0 == RADDR ? 11'he0 : _GEN_2148; // @[RAM_ST.scala 32:46]
  assign _GEN_2150 = 11'he1 == RADDR ? 11'he1 : _GEN_2149; // @[RAM_ST.scala 32:46]
  assign _GEN_2151 = 11'he2 == RADDR ? 11'he2 : _GEN_2150; // @[RAM_ST.scala 32:46]
  assign _GEN_2152 = 11'he3 == RADDR ? 11'he3 : _GEN_2151; // @[RAM_ST.scala 32:46]
  assign _GEN_2153 = 11'he4 == RADDR ? 11'he4 : _GEN_2152; // @[RAM_ST.scala 32:46]
  assign _GEN_2154 = 11'he5 == RADDR ? 11'he5 : _GEN_2153; // @[RAM_ST.scala 32:46]
  assign _GEN_2155 = 11'he6 == RADDR ? 11'he6 : _GEN_2154; // @[RAM_ST.scala 32:46]
  assign _GEN_2156 = 11'he7 == RADDR ? 11'he7 : _GEN_2155; // @[RAM_ST.scala 32:46]
  assign _GEN_2157 = 11'he8 == RADDR ? 11'he8 : _GEN_2156; // @[RAM_ST.scala 32:46]
  assign _GEN_2158 = 11'he9 == RADDR ? 11'he9 : _GEN_2157; // @[RAM_ST.scala 32:46]
  assign _GEN_2159 = 11'hea == RADDR ? 11'hea : _GEN_2158; // @[RAM_ST.scala 32:46]
  assign _GEN_2160 = 11'heb == RADDR ? 11'heb : _GEN_2159; // @[RAM_ST.scala 32:46]
  assign _GEN_2161 = 11'hec == RADDR ? 11'hec : _GEN_2160; // @[RAM_ST.scala 32:46]
  assign _GEN_2162 = 11'hed == RADDR ? 11'hed : _GEN_2161; // @[RAM_ST.scala 32:46]
  assign _GEN_2163 = 11'hee == RADDR ? 11'hee : _GEN_2162; // @[RAM_ST.scala 32:46]
  assign _GEN_2164 = 11'hef == RADDR ? 11'hef : _GEN_2163; // @[RAM_ST.scala 32:46]
  assign _GEN_2165 = 11'hf0 == RADDR ? 11'hf0 : _GEN_2164; // @[RAM_ST.scala 32:46]
  assign _GEN_2166 = 11'hf1 == RADDR ? 11'hf1 : _GEN_2165; // @[RAM_ST.scala 32:46]
  assign _GEN_2167 = 11'hf2 == RADDR ? 11'hf2 : _GEN_2166; // @[RAM_ST.scala 32:46]
  assign _GEN_2168 = 11'hf3 == RADDR ? 11'hf3 : _GEN_2167; // @[RAM_ST.scala 32:46]
  assign _GEN_2169 = 11'hf4 == RADDR ? 11'hf4 : _GEN_2168; // @[RAM_ST.scala 32:46]
  assign _GEN_2170 = 11'hf5 == RADDR ? 11'hf5 : _GEN_2169; // @[RAM_ST.scala 32:46]
  assign _GEN_2171 = 11'hf6 == RADDR ? 11'hf6 : _GEN_2170; // @[RAM_ST.scala 32:46]
  assign _GEN_2172 = 11'hf7 == RADDR ? 11'hf7 : _GEN_2171; // @[RAM_ST.scala 32:46]
  assign _GEN_2173 = 11'hf8 == RADDR ? 11'hf8 : _GEN_2172; // @[RAM_ST.scala 32:46]
  assign _GEN_2174 = 11'hf9 == RADDR ? 11'hf9 : _GEN_2173; // @[RAM_ST.scala 32:46]
  assign _GEN_2175 = 11'hfa == RADDR ? 11'hfa : _GEN_2174; // @[RAM_ST.scala 32:46]
  assign _GEN_2176 = 11'hfb == RADDR ? 11'hfb : _GEN_2175; // @[RAM_ST.scala 32:46]
  assign _GEN_2177 = 11'hfc == RADDR ? 11'hfc : _GEN_2176; // @[RAM_ST.scala 32:46]
  assign _GEN_2178 = 11'hfd == RADDR ? 11'hfd : _GEN_2177; // @[RAM_ST.scala 32:46]
  assign _GEN_2179 = 11'hfe == RADDR ? 11'hfe : _GEN_2178; // @[RAM_ST.scala 32:46]
  assign _GEN_2180 = 11'hff == RADDR ? 11'hff : _GEN_2179; // @[RAM_ST.scala 32:46]
  assign _GEN_2181 = 11'h100 == RADDR ? 11'h100 : _GEN_2180; // @[RAM_ST.scala 32:46]
  assign _GEN_2182 = 11'h101 == RADDR ? 11'h101 : _GEN_2181; // @[RAM_ST.scala 32:46]
  assign _GEN_2183 = 11'h102 == RADDR ? 11'h102 : _GEN_2182; // @[RAM_ST.scala 32:46]
  assign _GEN_2184 = 11'h103 == RADDR ? 11'h103 : _GEN_2183; // @[RAM_ST.scala 32:46]
  assign _GEN_2185 = 11'h104 == RADDR ? 11'h104 : _GEN_2184; // @[RAM_ST.scala 32:46]
  assign _GEN_2186 = 11'h105 == RADDR ? 11'h105 : _GEN_2185; // @[RAM_ST.scala 32:46]
  assign _GEN_2187 = 11'h106 == RADDR ? 11'h106 : _GEN_2186; // @[RAM_ST.scala 32:46]
  assign _GEN_2188 = 11'h107 == RADDR ? 11'h107 : _GEN_2187; // @[RAM_ST.scala 32:46]
  assign _GEN_2189 = 11'h108 == RADDR ? 11'h108 : _GEN_2188; // @[RAM_ST.scala 32:46]
  assign _GEN_2190 = 11'h109 == RADDR ? 11'h109 : _GEN_2189; // @[RAM_ST.scala 32:46]
  assign _GEN_2191 = 11'h10a == RADDR ? 11'h10a : _GEN_2190; // @[RAM_ST.scala 32:46]
  assign _GEN_2192 = 11'h10b == RADDR ? 11'h10b : _GEN_2191; // @[RAM_ST.scala 32:46]
  assign _GEN_2193 = 11'h10c == RADDR ? 11'h10c : _GEN_2192; // @[RAM_ST.scala 32:46]
  assign _GEN_2194 = 11'h10d == RADDR ? 11'h10d : _GEN_2193; // @[RAM_ST.scala 32:46]
  assign _GEN_2195 = 11'h10e == RADDR ? 11'h10e : _GEN_2194; // @[RAM_ST.scala 32:46]
  assign _GEN_2196 = 11'h10f == RADDR ? 11'h10f : _GEN_2195; // @[RAM_ST.scala 32:46]
  assign _GEN_2197 = 11'h110 == RADDR ? 11'h110 : _GEN_2196; // @[RAM_ST.scala 32:46]
  assign _GEN_2198 = 11'h111 == RADDR ? 11'h111 : _GEN_2197; // @[RAM_ST.scala 32:46]
  assign _GEN_2199 = 11'h112 == RADDR ? 11'h112 : _GEN_2198; // @[RAM_ST.scala 32:46]
  assign _GEN_2200 = 11'h113 == RADDR ? 11'h113 : _GEN_2199; // @[RAM_ST.scala 32:46]
  assign _GEN_2201 = 11'h114 == RADDR ? 11'h114 : _GEN_2200; // @[RAM_ST.scala 32:46]
  assign _GEN_2202 = 11'h115 == RADDR ? 11'h115 : _GEN_2201; // @[RAM_ST.scala 32:46]
  assign _GEN_2203 = 11'h116 == RADDR ? 11'h116 : _GEN_2202; // @[RAM_ST.scala 32:46]
  assign _GEN_2204 = 11'h117 == RADDR ? 11'h117 : _GEN_2203; // @[RAM_ST.scala 32:46]
  assign _GEN_2205 = 11'h118 == RADDR ? 11'h118 : _GEN_2204; // @[RAM_ST.scala 32:46]
  assign _GEN_2206 = 11'h119 == RADDR ? 11'h119 : _GEN_2205; // @[RAM_ST.scala 32:46]
  assign _GEN_2207 = 11'h11a == RADDR ? 11'h11a : _GEN_2206; // @[RAM_ST.scala 32:46]
  assign _GEN_2208 = 11'h11b == RADDR ? 11'h11b : _GEN_2207; // @[RAM_ST.scala 32:46]
  assign _GEN_2209 = 11'h11c == RADDR ? 11'h11c : _GEN_2208; // @[RAM_ST.scala 32:46]
  assign _GEN_2210 = 11'h11d == RADDR ? 11'h11d : _GEN_2209; // @[RAM_ST.scala 32:46]
  assign _GEN_2211 = 11'h11e == RADDR ? 11'h11e : _GEN_2210; // @[RAM_ST.scala 32:46]
  assign _GEN_2212 = 11'h11f == RADDR ? 11'h11f : _GEN_2211; // @[RAM_ST.scala 32:46]
  assign _GEN_2213 = 11'h120 == RADDR ? 11'h120 : _GEN_2212; // @[RAM_ST.scala 32:46]
  assign _GEN_2214 = 11'h121 == RADDR ? 11'h121 : _GEN_2213; // @[RAM_ST.scala 32:46]
  assign _GEN_2215 = 11'h122 == RADDR ? 11'h122 : _GEN_2214; // @[RAM_ST.scala 32:46]
  assign _GEN_2216 = 11'h123 == RADDR ? 11'h123 : _GEN_2215; // @[RAM_ST.scala 32:46]
  assign _GEN_2217 = 11'h124 == RADDR ? 11'h124 : _GEN_2216; // @[RAM_ST.scala 32:46]
  assign _GEN_2218 = 11'h125 == RADDR ? 11'h125 : _GEN_2217; // @[RAM_ST.scala 32:46]
  assign _GEN_2219 = 11'h126 == RADDR ? 11'h126 : _GEN_2218; // @[RAM_ST.scala 32:46]
  assign _GEN_2220 = 11'h127 == RADDR ? 11'h127 : _GEN_2219; // @[RAM_ST.scala 32:46]
  assign _GEN_2221 = 11'h128 == RADDR ? 11'h128 : _GEN_2220; // @[RAM_ST.scala 32:46]
  assign _GEN_2222 = 11'h129 == RADDR ? 11'h129 : _GEN_2221; // @[RAM_ST.scala 32:46]
  assign _GEN_2223 = 11'h12a == RADDR ? 11'h12a : _GEN_2222; // @[RAM_ST.scala 32:46]
  assign _GEN_2224 = 11'h12b == RADDR ? 11'h12b : _GEN_2223; // @[RAM_ST.scala 32:46]
  assign _GEN_2225 = 11'h12c == RADDR ? 11'h12c : _GEN_2224; // @[RAM_ST.scala 32:46]
  assign _GEN_2226 = 11'h12d == RADDR ? 11'h12d : _GEN_2225; // @[RAM_ST.scala 32:46]
  assign _GEN_2227 = 11'h12e == RADDR ? 11'h12e : _GEN_2226; // @[RAM_ST.scala 32:46]
  assign _GEN_2228 = 11'h12f == RADDR ? 11'h12f : _GEN_2227; // @[RAM_ST.scala 32:46]
  assign _GEN_2229 = 11'h130 == RADDR ? 11'h130 : _GEN_2228; // @[RAM_ST.scala 32:46]
  assign _GEN_2230 = 11'h131 == RADDR ? 11'h131 : _GEN_2229; // @[RAM_ST.scala 32:46]
  assign _GEN_2231 = 11'h132 == RADDR ? 11'h132 : _GEN_2230; // @[RAM_ST.scala 32:46]
  assign _GEN_2232 = 11'h133 == RADDR ? 11'h133 : _GEN_2231; // @[RAM_ST.scala 32:46]
  assign _GEN_2233 = 11'h134 == RADDR ? 11'h134 : _GEN_2232; // @[RAM_ST.scala 32:46]
  assign _GEN_2234 = 11'h135 == RADDR ? 11'h135 : _GEN_2233; // @[RAM_ST.scala 32:46]
  assign _GEN_2235 = 11'h136 == RADDR ? 11'h136 : _GEN_2234; // @[RAM_ST.scala 32:46]
  assign _GEN_2236 = 11'h137 == RADDR ? 11'h137 : _GEN_2235; // @[RAM_ST.scala 32:46]
  assign _GEN_2237 = 11'h138 == RADDR ? 11'h138 : _GEN_2236; // @[RAM_ST.scala 32:46]
  assign _GEN_2238 = 11'h139 == RADDR ? 11'h139 : _GEN_2237; // @[RAM_ST.scala 32:46]
  assign _GEN_2239 = 11'h13a == RADDR ? 11'h13a : _GEN_2238; // @[RAM_ST.scala 32:46]
  assign _GEN_2240 = 11'h13b == RADDR ? 11'h13b : _GEN_2239; // @[RAM_ST.scala 32:46]
  assign _GEN_2241 = 11'h13c == RADDR ? 11'h13c : _GEN_2240; // @[RAM_ST.scala 32:46]
  assign _GEN_2242 = 11'h13d == RADDR ? 11'h13d : _GEN_2241; // @[RAM_ST.scala 32:46]
  assign _GEN_2243 = 11'h13e == RADDR ? 11'h13e : _GEN_2242; // @[RAM_ST.scala 32:46]
  assign _GEN_2244 = 11'h13f == RADDR ? 11'h13f : _GEN_2243; // @[RAM_ST.scala 32:46]
  assign _GEN_2245 = 11'h140 == RADDR ? 11'h140 : _GEN_2244; // @[RAM_ST.scala 32:46]
  assign _GEN_2246 = 11'h141 == RADDR ? 11'h141 : _GEN_2245; // @[RAM_ST.scala 32:46]
  assign _GEN_2247 = 11'h142 == RADDR ? 11'h142 : _GEN_2246; // @[RAM_ST.scala 32:46]
  assign _GEN_2248 = 11'h143 == RADDR ? 11'h143 : _GEN_2247; // @[RAM_ST.scala 32:46]
  assign _GEN_2249 = 11'h144 == RADDR ? 11'h144 : _GEN_2248; // @[RAM_ST.scala 32:46]
  assign _GEN_2250 = 11'h145 == RADDR ? 11'h145 : _GEN_2249; // @[RAM_ST.scala 32:46]
  assign _GEN_2251 = 11'h146 == RADDR ? 11'h146 : _GEN_2250; // @[RAM_ST.scala 32:46]
  assign _GEN_2252 = 11'h147 == RADDR ? 11'h147 : _GEN_2251; // @[RAM_ST.scala 32:46]
  assign _GEN_2253 = 11'h148 == RADDR ? 11'h148 : _GEN_2252; // @[RAM_ST.scala 32:46]
  assign _GEN_2254 = 11'h149 == RADDR ? 11'h149 : _GEN_2253; // @[RAM_ST.scala 32:46]
  assign _GEN_2255 = 11'h14a == RADDR ? 11'h14a : _GEN_2254; // @[RAM_ST.scala 32:46]
  assign _GEN_2256 = 11'h14b == RADDR ? 11'h14b : _GEN_2255; // @[RAM_ST.scala 32:46]
  assign _GEN_2257 = 11'h14c == RADDR ? 11'h14c : _GEN_2256; // @[RAM_ST.scala 32:46]
  assign _GEN_2258 = 11'h14d == RADDR ? 11'h14d : _GEN_2257; // @[RAM_ST.scala 32:46]
  assign _GEN_2259 = 11'h14e == RADDR ? 11'h14e : _GEN_2258; // @[RAM_ST.scala 32:46]
  assign _GEN_2260 = 11'h14f == RADDR ? 11'h14f : _GEN_2259; // @[RAM_ST.scala 32:46]
  assign _GEN_2261 = 11'h150 == RADDR ? 11'h150 : _GEN_2260; // @[RAM_ST.scala 32:46]
  assign _GEN_2262 = 11'h151 == RADDR ? 11'h151 : _GEN_2261; // @[RAM_ST.scala 32:46]
  assign _GEN_2263 = 11'h152 == RADDR ? 11'h152 : _GEN_2262; // @[RAM_ST.scala 32:46]
  assign _GEN_2264 = 11'h153 == RADDR ? 11'h153 : _GEN_2263; // @[RAM_ST.scala 32:46]
  assign _GEN_2265 = 11'h154 == RADDR ? 11'h154 : _GEN_2264; // @[RAM_ST.scala 32:46]
  assign _GEN_2266 = 11'h155 == RADDR ? 11'h155 : _GEN_2265; // @[RAM_ST.scala 32:46]
  assign _GEN_2267 = 11'h156 == RADDR ? 11'h156 : _GEN_2266; // @[RAM_ST.scala 32:46]
  assign _GEN_2268 = 11'h157 == RADDR ? 11'h157 : _GEN_2267; // @[RAM_ST.scala 32:46]
  assign _GEN_2269 = 11'h158 == RADDR ? 11'h158 : _GEN_2268; // @[RAM_ST.scala 32:46]
  assign _GEN_2270 = 11'h159 == RADDR ? 11'h159 : _GEN_2269; // @[RAM_ST.scala 32:46]
  assign _GEN_2271 = 11'h15a == RADDR ? 11'h15a : _GEN_2270; // @[RAM_ST.scala 32:46]
  assign _GEN_2272 = 11'h15b == RADDR ? 11'h15b : _GEN_2271; // @[RAM_ST.scala 32:46]
  assign _GEN_2273 = 11'h15c == RADDR ? 11'h15c : _GEN_2272; // @[RAM_ST.scala 32:46]
  assign _GEN_2274 = 11'h15d == RADDR ? 11'h15d : _GEN_2273; // @[RAM_ST.scala 32:46]
  assign _GEN_2275 = 11'h15e == RADDR ? 11'h15e : _GEN_2274; // @[RAM_ST.scala 32:46]
  assign _GEN_2276 = 11'h15f == RADDR ? 11'h15f : _GEN_2275; // @[RAM_ST.scala 32:46]
  assign _GEN_2277 = 11'h160 == RADDR ? 11'h160 : _GEN_2276; // @[RAM_ST.scala 32:46]
  assign _GEN_2278 = 11'h161 == RADDR ? 11'h161 : _GEN_2277; // @[RAM_ST.scala 32:46]
  assign _GEN_2279 = 11'h162 == RADDR ? 11'h162 : _GEN_2278; // @[RAM_ST.scala 32:46]
  assign _GEN_2280 = 11'h163 == RADDR ? 11'h163 : _GEN_2279; // @[RAM_ST.scala 32:46]
  assign _GEN_2281 = 11'h164 == RADDR ? 11'h164 : _GEN_2280; // @[RAM_ST.scala 32:46]
  assign _GEN_2282 = 11'h165 == RADDR ? 11'h165 : _GEN_2281; // @[RAM_ST.scala 32:46]
  assign _GEN_2283 = 11'h166 == RADDR ? 11'h166 : _GEN_2282; // @[RAM_ST.scala 32:46]
  assign _GEN_2284 = 11'h167 == RADDR ? 11'h167 : _GEN_2283; // @[RAM_ST.scala 32:46]
  assign _GEN_2285 = 11'h168 == RADDR ? 11'h168 : _GEN_2284; // @[RAM_ST.scala 32:46]
  assign _GEN_2286 = 11'h169 == RADDR ? 11'h169 : _GEN_2285; // @[RAM_ST.scala 32:46]
  assign _GEN_2287 = 11'h16a == RADDR ? 11'h16a : _GEN_2286; // @[RAM_ST.scala 32:46]
  assign _GEN_2288 = 11'h16b == RADDR ? 11'h16b : _GEN_2287; // @[RAM_ST.scala 32:46]
  assign _GEN_2289 = 11'h16c == RADDR ? 11'h16c : _GEN_2288; // @[RAM_ST.scala 32:46]
  assign _GEN_2290 = 11'h16d == RADDR ? 11'h16d : _GEN_2289; // @[RAM_ST.scala 32:46]
  assign _GEN_2291 = 11'h16e == RADDR ? 11'h16e : _GEN_2290; // @[RAM_ST.scala 32:46]
  assign _GEN_2292 = 11'h16f == RADDR ? 11'h16f : _GEN_2291; // @[RAM_ST.scala 32:46]
  assign _GEN_2293 = 11'h170 == RADDR ? 11'h170 : _GEN_2292; // @[RAM_ST.scala 32:46]
  assign _GEN_2294 = 11'h171 == RADDR ? 11'h171 : _GEN_2293; // @[RAM_ST.scala 32:46]
  assign _GEN_2295 = 11'h172 == RADDR ? 11'h172 : _GEN_2294; // @[RAM_ST.scala 32:46]
  assign _GEN_2296 = 11'h173 == RADDR ? 11'h173 : _GEN_2295; // @[RAM_ST.scala 32:46]
  assign _GEN_2297 = 11'h174 == RADDR ? 11'h174 : _GEN_2296; // @[RAM_ST.scala 32:46]
  assign _GEN_2298 = 11'h175 == RADDR ? 11'h175 : _GEN_2297; // @[RAM_ST.scala 32:46]
  assign _GEN_2299 = 11'h176 == RADDR ? 11'h176 : _GEN_2298; // @[RAM_ST.scala 32:46]
  assign _GEN_2300 = 11'h177 == RADDR ? 11'h177 : _GEN_2299; // @[RAM_ST.scala 32:46]
  assign _GEN_2301 = 11'h178 == RADDR ? 11'h178 : _GEN_2300; // @[RAM_ST.scala 32:46]
  assign _GEN_2302 = 11'h179 == RADDR ? 11'h179 : _GEN_2301; // @[RAM_ST.scala 32:46]
  assign _GEN_2303 = 11'h17a == RADDR ? 11'h17a : _GEN_2302; // @[RAM_ST.scala 32:46]
  assign _GEN_2304 = 11'h17b == RADDR ? 11'h17b : _GEN_2303; // @[RAM_ST.scala 32:46]
  assign _GEN_2305 = 11'h17c == RADDR ? 11'h17c : _GEN_2304; // @[RAM_ST.scala 32:46]
  assign _GEN_2306 = 11'h17d == RADDR ? 11'h17d : _GEN_2305; // @[RAM_ST.scala 32:46]
  assign _GEN_2307 = 11'h17e == RADDR ? 11'h17e : _GEN_2306; // @[RAM_ST.scala 32:46]
  assign _GEN_2308 = 11'h17f == RADDR ? 11'h17f : _GEN_2307; // @[RAM_ST.scala 32:46]
  assign _GEN_2309 = 11'h180 == RADDR ? 11'h180 : _GEN_2308; // @[RAM_ST.scala 32:46]
  assign _GEN_2310 = 11'h181 == RADDR ? 11'h181 : _GEN_2309; // @[RAM_ST.scala 32:46]
  assign _GEN_2311 = 11'h182 == RADDR ? 11'h182 : _GEN_2310; // @[RAM_ST.scala 32:46]
  assign _GEN_2312 = 11'h183 == RADDR ? 11'h183 : _GEN_2311; // @[RAM_ST.scala 32:46]
  assign _GEN_2313 = 11'h184 == RADDR ? 11'h184 : _GEN_2312; // @[RAM_ST.scala 32:46]
  assign _GEN_2314 = 11'h185 == RADDR ? 11'h185 : _GEN_2313; // @[RAM_ST.scala 32:46]
  assign _GEN_2315 = 11'h186 == RADDR ? 11'h186 : _GEN_2314; // @[RAM_ST.scala 32:46]
  assign _GEN_2316 = 11'h187 == RADDR ? 11'h187 : _GEN_2315; // @[RAM_ST.scala 32:46]
  assign _GEN_2317 = 11'h188 == RADDR ? 11'h188 : _GEN_2316; // @[RAM_ST.scala 32:46]
  assign _GEN_2318 = 11'h189 == RADDR ? 11'h189 : _GEN_2317; // @[RAM_ST.scala 32:46]
  assign _GEN_2319 = 11'h18a == RADDR ? 11'h18a : _GEN_2318; // @[RAM_ST.scala 32:46]
  assign _GEN_2320 = 11'h18b == RADDR ? 11'h18b : _GEN_2319; // @[RAM_ST.scala 32:46]
  assign _GEN_2321 = 11'h18c == RADDR ? 11'h18c : _GEN_2320; // @[RAM_ST.scala 32:46]
  assign _GEN_2322 = 11'h18d == RADDR ? 11'h18d : _GEN_2321; // @[RAM_ST.scala 32:46]
  assign _GEN_2323 = 11'h18e == RADDR ? 11'h18e : _GEN_2322; // @[RAM_ST.scala 32:46]
  assign _GEN_2324 = 11'h18f == RADDR ? 11'h18f : _GEN_2323; // @[RAM_ST.scala 32:46]
  assign _GEN_2325 = 11'h190 == RADDR ? 11'h190 : _GEN_2324; // @[RAM_ST.scala 32:46]
  assign _GEN_2326 = 11'h191 == RADDR ? 11'h191 : _GEN_2325; // @[RAM_ST.scala 32:46]
  assign _GEN_2327 = 11'h192 == RADDR ? 11'h192 : _GEN_2326; // @[RAM_ST.scala 32:46]
  assign _GEN_2328 = 11'h193 == RADDR ? 11'h193 : _GEN_2327; // @[RAM_ST.scala 32:46]
  assign _GEN_2329 = 11'h194 == RADDR ? 11'h194 : _GEN_2328; // @[RAM_ST.scala 32:46]
  assign _GEN_2330 = 11'h195 == RADDR ? 11'h195 : _GEN_2329; // @[RAM_ST.scala 32:46]
  assign _GEN_2331 = 11'h196 == RADDR ? 11'h196 : _GEN_2330; // @[RAM_ST.scala 32:46]
  assign _GEN_2332 = 11'h197 == RADDR ? 11'h197 : _GEN_2331; // @[RAM_ST.scala 32:46]
  assign _GEN_2333 = 11'h198 == RADDR ? 11'h198 : _GEN_2332; // @[RAM_ST.scala 32:46]
  assign _GEN_2334 = 11'h199 == RADDR ? 11'h199 : _GEN_2333; // @[RAM_ST.scala 32:46]
  assign _GEN_2335 = 11'h19a == RADDR ? 11'h19a : _GEN_2334; // @[RAM_ST.scala 32:46]
  assign _GEN_2336 = 11'h19b == RADDR ? 11'h19b : _GEN_2335; // @[RAM_ST.scala 32:46]
  assign _GEN_2337 = 11'h19c == RADDR ? 11'h19c : _GEN_2336; // @[RAM_ST.scala 32:46]
  assign _GEN_2338 = 11'h19d == RADDR ? 11'h19d : _GEN_2337; // @[RAM_ST.scala 32:46]
  assign _GEN_2339 = 11'h19e == RADDR ? 11'h19e : _GEN_2338; // @[RAM_ST.scala 32:46]
  assign _GEN_2340 = 11'h19f == RADDR ? 11'h19f : _GEN_2339; // @[RAM_ST.scala 32:46]
  assign _GEN_2341 = 11'h1a0 == RADDR ? 11'h1a0 : _GEN_2340; // @[RAM_ST.scala 32:46]
  assign _GEN_2342 = 11'h1a1 == RADDR ? 11'h1a1 : _GEN_2341; // @[RAM_ST.scala 32:46]
  assign _GEN_2343 = 11'h1a2 == RADDR ? 11'h1a2 : _GEN_2342; // @[RAM_ST.scala 32:46]
  assign _GEN_2344 = 11'h1a3 == RADDR ? 11'h1a3 : _GEN_2343; // @[RAM_ST.scala 32:46]
  assign _GEN_2345 = 11'h1a4 == RADDR ? 11'h1a4 : _GEN_2344; // @[RAM_ST.scala 32:46]
  assign _GEN_2346 = 11'h1a5 == RADDR ? 11'h1a5 : _GEN_2345; // @[RAM_ST.scala 32:46]
  assign _GEN_2347 = 11'h1a6 == RADDR ? 11'h1a6 : _GEN_2346; // @[RAM_ST.scala 32:46]
  assign _GEN_2348 = 11'h1a7 == RADDR ? 11'h1a7 : _GEN_2347; // @[RAM_ST.scala 32:46]
  assign _GEN_2349 = 11'h1a8 == RADDR ? 11'h1a8 : _GEN_2348; // @[RAM_ST.scala 32:46]
  assign _GEN_2350 = 11'h1a9 == RADDR ? 11'h1a9 : _GEN_2349; // @[RAM_ST.scala 32:46]
  assign _GEN_2351 = 11'h1aa == RADDR ? 11'h1aa : _GEN_2350; // @[RAM_ST.scala 32:46]
  assign _GEN_2352 = 11'h1ab == RADDR ? 11'h1ab : _GEN_2351; // @[RAM_ST.scala 32:46]
  assign _GEN_2353 = 11'h1ac == RADDR ? 11'h1ac : _GEN_2352; // @[RAM_ST.scala 32:46]
  assign _GEN_2354 = 11'h1ad == RADDR ? 11'h1ad : _GEN_2353; // @[RAM_ST.scala 32:46]
  assign _GEN_2355 = 11'h1ae == RADDR ? 11'h1ae : _GEN_2354; // @[RAM_ST.scala 32:46]
  assign _GEN_2356 = 11'h1af == RADDR ? 11'h1af : _GEN_2355; // @[RAM_ST.scala 32:46]
  assign _GEN_2357 = 11'h1b0 == RADDR ? 11'h1b0 : _GEN_2356; // @[RAM_ST.scala 32:46]
  assign _GEN_2358 = 11'h1b1 == RADDR ? 11'h1b1 : _GEN_2357; // @[RAM_ST.scala 32:46]
  assign _GEN_2359 = 11'h1b2 == RADDR ? 11'h1b2 : _GEN_2358; // @[RAM_ST.scala 32:46]
  assign _GEN_2360 = 11'h1b3 == RADDR ? 11'h1b3 : _GEN_2359; // @[RAM_ST.scala 32:46]
  assign _GEN_2361 = 11'h1b4 == RADDR ? 11'h1b4 : _GEN_2360; // @[RAM_ST.scala 32:46]
  assign _GEN_2362 = 11'h1b5 == RADDR ? 11'h1b5 : _GEN_2361; // @[RAM_ST.scala 32:46]
  assign _GEN_2363 = 11'h1b6 == RADDR ? 11'h1b6 : _GEN_2362; // @[RAM_ST.scala 32:46]
  assign _GEN_2364 = 11'h1b7 == RADDR ? 11'h1b7 : _GEN_2363; // @[RAM_ST.scala 32:46]
  assign _GEN_2365 = 11'h1b8 == RADDR ? 11'h1b8 : _GEN_2364; // @[RAM_ST.scala 32:46]
  assign _GEN_2366 = 11'h1b9 == RADDR ? 11'h1b9 : _GEN_2365; // @[RAM_ST.scala 32:46]
  assign _GEN_2367 = 11'h1ba == RADDR ? 11'h1ba : _GEN_2366; // @[RAM_ST.scala 32:46]
  assign _GEN_2368 = 11'h1bb == RADDR ? 11'h1bb : _GEN_2367; // @[RAM_ST.scala 32:46]
  assign _GEN_2369 = 11'h1bc == RADDR ? 11'h1bc : _GEN_2368; // @[RAM_ST.scala 32:46]
  assign _GEN_2370 = 11'h1bd == RADDR ? 11'h1bd : _GEN_2369; // @[RAM_ST.scala 32:46]
  assign _GEN_2371 = 11'h1be == RADDR ? 11'h1be : _GEN_2370; // @[RAM_ST.scala 32:46]
  assign _GEN_2372 = 11'h1bf == RADDR ? 11'h1bf : _GEN_2371; // @[RAM_ST.scala 32:46]
  assign _GEN_2373 = 11'h1c0 == RADDR ? 11'h1c0 : _GEN_2372; // @[RAM_ST.scala 32:46]
  assign _GEN_2374 = 11'h1c1 == RADDR ? 11'h1c1 : _GEN_2373; // @[RAM_ST.scala 32:46]
  assign _GEN_2375 = 11'h1c2 == RADDR ? 11'h1c2 : _GEN_2374; // @[RAM_ST.scala 32:46]
  assign _GEN_2376 = 11'h1c3 == RADDR ? 11'h1c3 : _GEN_2375; // @[RAM_ST.scala 32:46]
  assign _GEN_2377 = 11'h1c4 == RADDR ? 11'h1c4 : _GEN_2376; // @[RAM_ST.scala 32:46]
  assign _GEN_2378 = 11'h1c5 == RADDR ? 11'h1c5 : _GEN_2377; // @[RAM_ST.scala 32:46]
  assign _GEN_2379 = 11'h1c6 == RADDR ? 11'h1c6 : _GEN_2378; // @[RAM_ST.scala 32:46]
  assign _GEN_2380 = 11'h1c7 == RADDR ? 11'h1c7 : _GEN_2379; // @[RAM_ST.scala 32:46]
  assign _GEN_2381 = 11'h1c8 == RADDR ? 11'h1c8 : _GEN_2380; // @[RAM_ST.scala 32:46]
  assign _GEN_2382 = 11'h1c9 == RADDR ? 11'h1c9 : _GEN_2381; // @[RAM_ST.scala 32:46]
  assign _GEN_2383 = 11'h1ca == RADDR ? 11'h1ca : _GEN_2382; // @[RAM_ST.scala 32:46]
  assign _GEN_2384 = 11'h1cb == RADDR ? 11'h1cb : _GEN_2383; // @[RAM_ST.scala 32:46]
  assign _GEN_2385 = 11'h1cc == RADDR ? 11'h1cc : _GEN_2384; // @[RAM_ST.scala 32:46]
  assign _GEN_2386 = 11'h1cd == RADDR ? 11'h1cd : _GEN_2385; // @[RAM_ST.scala 32:46]
  assign _GEN_2387 = 11'h1ce == RADDR ? 11'h1ce : _GEN_2386; // @[RAM_ST.scala 32:46]
  assign _GEN_2388 = 11'h1cf == RADDR ? 11'h1cf : _GEN_2387; // @[RAM_ST.scala 32:46]
  assign _GEN_2389 = 11'h1d0 == RADDR ? 11'h1d0 : _GEN_2388; // @[RAM_ST.scala 32:46]
  assign _GEN_2390 = 11'h1d1 == RADDR ? 11'h1d1 : _GEN_2389; // @[RAM_ST.scala 32:46]
  assign _GEN_2391 = 11'h1d2 == RADDR ? 11'h1d2 : _GEN_2390; // @[RAM_ST.scala 32:46]
  assign _GEN_2392 = 11'h1d3 == RADDR ? 11'h1d3 : _GEN_2391; // @[RAM_ST.scala 32:46]
  assign _GEN_2393 = 11'h1d4 == RADDR ? 11'h1d4 : _GEN_2392; // @[RAM_ST.scala 32:46]
  assign _GEN_2394 = 11'h1d5 == RADDR ? 11'h1d5 : _GEN_2393; // @[RAM_ST.scala 32:46]
  assign _GEN_2395 = 11'h1d6 == RADDR ? 11'h1d6 : _GEN_2394; // @[RAM_ST.scala 32:46]
  assign _GEN_2396 = 11'h1d7 == RADDR ? 11'h1d7 : _GEN_2395; // @[RAM_ST.scala 32:46]
  assign _GEN_2397 = 11'h1d8 == RADDR ? 11'h1d8 : _GEN_2396; // @[RAM_ST.scala 32:46]
  assign _GEN_2398 = 11'h1d9 == RADDR ? 11'h1d9 : _GEN_2397; // @[RAM_ST.scala 32:46]
  assign _GEN_2399 = 11'h1da == RADDR ? 11'h1da : _GEN_2398; // @[RAM_ST.scala 32:46]
  assign _GEN_2400 = 11'h1db == RADDR ? 11'h1db : _GEN_2399; // @[RAM_ST.scala 32:46]
  assign _GEN_2401 = 11'h1dc == RADDR ? 11'h1dc : _GEN_2400; // @[RAM_ST.scala 32:46]
  assign _GEN_2402 = 11'h1dd == RADDR ? 11'h1dd : _GEN_2401; // @[RAM_ST.scala 32:46]
  assign _GEN_2403 = 11'h1de == RADDR ? 11'h1de : _GEN_2402; // @[RAM_ST.scala 32:46]
  assign _GEN_2404 = 11'h1df == RADDR ? 11'h1df : _GEN_2403; // @[RAM_ST.scala 32:46]
  assign _GEN_2405 = 11'h1e0 == RADDR ? 11'h1e0 : _GEN_2404; // @[RAM_ST.scala 32:46]
  assign _GEN_2406 = 11'h1e1 == RADDR ? 11'h1e1 : _GEN_2405; // @[RAM_ST.scala 32:46]
  assign _GEN_2407 = 11'h1e2 == RADDR ? 11'h1e2 : _GEN_2406; // @[RAM_ST.scala 32:46]
  assign _GEN_2408 = 11'h1e3 == RADDR ? 11'h1e3 : _GEN_2407; // @[RAM_ST.scala 32:46]
  assign _GEN_2409 = 11'h1e4 == RADDR ? 11'h1e4 : _GEN_2408; // @[RAM_ST.scala 32:46]
  assign _GEN_2410 = 11'h1e5 == RADDR ? 11'h1e5 : _GEN_2409; // @[RAM_ST.scala 32:46]
  assign _GEN_2411 = 11'h1e6 == RADDR ? 11'h1e6 : _GEN_2410; // @[RAM_ST.scala 32:46]
  assign _GEN_2412 = 11'h1e7 == RADDR ? 11'h1e7 : _GEN_2411; // @[RAM_ST.scala 32:46]
  assign _GEN_2413 = 11'h1e8 == RADDR ? 11'h1e8 : _GEN_2412; // @[RAM_ST.scala 32:46]
  assign _GEN_2414 = 11'h1e9 == RADDR ? 11'h1e9 : _GEN_2413; // @[RAM_ST.scala 32:46]
  assign _GEN_2415 = 11'h1ea == RADDR ? 11'h1ea : _GEN_2414; // @[RAM_ST.scala 32:46]
  assign _GEN_2416 = 11'h1eb == RADDR ? 11'h1eb : _GEN_2415; // @[RAM_ST.scala 32:46]
  assign _GEN_2417 = 11'h1ec == RADDR ? 11'h1ec : _GEN_2416; // @[RAM_ST.scala 32:46]
  assign _GEN_2418 = 11'h1ed == RADDR ? 11'h1ed : _GEN_2417; // @[RAM_ST.scala 32:46]
  assign _GEN_2419 = 11'h1ee == RADDR ? 11'h1ee : _GEN_2418; // @[RAM_ST.scala 32:46]
  assign _GEN_2420 = 11'h1ef == RADDR ? 11'h1ef : _GEN_2419; // @[RAM_ST.scala 32:46]
  assign _GEN_2421 = 11'h1f0 == RADDR ? 11'h1f0 : _GEN_2420; // @[RAM_ST.scala 32:46]
  assign _GEN_2422 = 11'h1f1 == RADDR ? 11'h1f1 : _GEN_2421; // @[RAM_ST.scala 32:46]
  assign _GEN_2423 = 11'h1f2 == RADDR ? 11'h1f2 : _GEN_2422; // @[RAM_ST.scala 32:46]
  assign _GEN_2424 = 11'h1f3 == RADDR ? 11'h1f3 : _GEN_2423; // @[RAM_ST.scala 32:46]
  assign _GEN_2425 = 11'h1f4 == RADDR ? 11'h1f4 : _GEN_2424; // @[RAM_ST.scala 32:46]
  assign _GEN_2426 = 11'h1f5 == RADDR ? 11'h1f5 : _GEN_2425; // @[RAM_ST.scala 32:46]
  assign _GEN_2427 = 11'h1f6 == RADDR ? 11'h1f6 : _GEN_2426; // @[RAM_ST.scala 32:46]
  assign _GEN_2428 = 11'h1f7 == RADDR ? 11'h1f7 : _GEN_2427; // @[RAM_ST.scala 32:46]
  assign _GEN_2429 = 11'h1f8 == RADDR ? 11'h1f8 : _GEN_2428; // @[RAM_ST.scala 32:46]
  assign _GEN_2430 = 11'h1f9 == RADDR ? 11'h1f9 : _GEN_2429; // @[RAM_ST.scala 32:46]
  assign _GEN_2431 = 11'h1fa == RADDR ? 11'h1fa : _GEN_2430; // @[RAM_ST.scala 32:46]
  assign _GEN_2432 = 11'h1fb == RADDR ? 11'h1fb : _GEN_2431; // @[RAM_ST.scala 32:46]
  assign _GEN_2433 = 11'h1fc == RADDR ? 11'h1fc : _GEN_2432; // @[RAM_ST.scala 32:46]
  assign _GEN_2434 = 11'h1fd == RADDR ? 11'h1fd : _GEN_2433; // @[RAM_ST.scala 32:46]
  assign _GEN_2435 = 11'h1fe == RADDR ? 11'h1fe : _GEN_2434; // @[RAM_ST.scala 32:46]
  assign _GEN_2436 = 11'h1ff == RADDR ? 11'h1ff : _GEN_2435; // @[RAM_ST.scala 32:46]
  assign _GEN_2437 = 11'h200 == RADDR ? 11'h200 : _GEN_2436; // @[RAM_ST.scala 32:46]
  assign _GEN_2438 = 11'h201 == RADDR ? 11'h201 : _GEN_2437; // @[RAM_ST.scala 32:46]
  assign _GEN_2439 = 11'h202 == RADDR ? 11'h202 : _GEN_2438; // @[RAM_ST.scala 32:46]
  assign _GEN_2440 = 11'h203 == RADDR ? 11'h203 : _GEN_2439; // @[RAM_ST.scala 32:46]
  assign _GEN_2441 = 11'h204 == RADDR ? 11'h204 : _GEN_2440; // @[RAM_ST.scala 32:46]
  assign _GEN_2442 = 11'h205 == RADDR ? 11'h205 : _GEN_2441; // @[RAM_ST.scala 32:46]
  assign _GEN_2443 = 11'h206 == RADDR ? 11'h206 : _GEN_2442; // @[RAM_ST.scala 32:46]
  assign _GEN_2444 = 11'h207 == RADDR ? 11'h207 : _GEN_2443; // @[RAM_ST.scala 32:46]
  assign _GEN_2445 = 11'h208 == RADDR ? 11'h208 : _GEN_2444; // @[RAM_ST.scala 32:46]
  assign _GEN_2446 = 11'h209 == RADDR ? 11'h209 : _GEN_2445; // @[RAM_ST.scala 32:46]
  assign _GEN_2447 = 11'h20a == RADDR ? 11'h20a : _GEN_2446; // @[RAM_ST.scala 32:46]
  assign _GEN_2448 = 11'h20b == RADDR ? 11'h20b : _GEN_2447; // @[RAM_ST.scala 32:46]
  assign _GEN_2449 = 11'h20c == RADDR ? 11'h20c : _GEN_2448; // @[RAM_ST.scala 32:46]
  assign _GEN_2450 = 11'h20d == RADDR ? 11'h20d : _GEN_2449; // @[RAM_ST.scala 32:46]
  assign _GEN_2451 = 11'h20e == RADDR ? 11'h20e : _GEN_2450; // @[RAM_ST.scala 32:46]
  assign _GEN_2452 = 11'h20f == RADDR ? 11'h20f : _GEN_2451; // @[RAM_ST.scala 32:46]
  assign _GEN_2453 = 11'h210 == RADDR ? 11'h210 : _GEN_2452; // @[RAM_ST.scala 32:46]
  assign _GEN_2454 = 11'h211 == RADDR ? 11'h211 : _GEN_2453; // @[RAM_ST.scala 32:46]
  assign _GEN_2455 = 11'h212 == RADDR ? 11'h212 : _GEN_2454; // @[RAM_ST.scala 32:46]
  assign _GEN_2456 = 11'h213 == RADDR ? 11'h213 : _GEN_2455; // @[RAM_ST.scala 32:46]
  assign _GEN_2457 = 11'h214 == RADDR ? 11'h214 : _GEN_2456; // @[RAM_ST.scala 32:46]
  assign _GEN_2458 = 11'h215 == RADDR ? 11'h215 : _GEN_2457; // @[RAM_ST.scala 32:46]
  assign _GEN_2459 = 11'h216 == RADDR ? 11'h216 : _GEN_2458; // @[RAM_ST.scala 32:46]
  assign _GEN_2460 = 11'h217 == RADDR ? 11'h217 : _GEN_2459; // @[RAM_ST.scala 32:46]
  assign _GEN_2461 = 11'h218 == RADDR ? 11'h218 : _GEN_2460; // @[RAM_ST.scala 32:46]
  assign _GEN_2462 = 11'h219 == RADDR ? 11'h219 : _GEN_2461; // @[RAM_ST.scala 32:46]
  assign _GEN_2463 = 11'h21a == RADDR ? 11'h21a : _GEN_2462; // @[RAM_ST.scala 32:46]
  assign _GEN_2464 = 11'h21b == RADDR ? 11'h21b : _GEN_2463; // @[RAM_ST.scala 32:46]
  assign _GEN_2465 = 11'h21c == RADDR ? 11'h21c : _GEN_2464; // @[RAM_ST.scala 32:46]
  assign _GEN_2466 = 11'h21d == RADDR ? 11'h21d : _GEN_2465; // @[RAM_ST.scala 32:46]
  assign _GEN_2467 = 11'h21e == RADDR ? 11'h21e : _GEN_2466; // @[RAM_ST.scala 32:46]
  assign _GEN_2468 = 11'h21f == RADDR ? 11'h21f : _GEN_2467; // @[RAM_ST.scala 32:46]
  assign _GEN_2469 = 11'h220 == RADDR ? 11'h220 : _GEN_2468; // @[RAM_ST.scala 32:46]
  assign _GEN_2470 = 11'h221 == RADDR ? 11'h221 : _GEN_2469; // @[RAM_ST.scala 32:46]
  assign _GEN_2471 = 11'h222 == RADDR ? 11'h222 : _GEN_2470; // @[RAM_ST.scala 32:46]
  assign _GEN_2472 = 11'h223 == RADDR ? 11'h223 : _GEN_2471; // @[RAM_ST.scala 32:46]
  assign _GEN_2473 = 11'h224 == RADDR ? 11'h224 : _GEN_2472; // @[RAM_ST.scala 32:46]
  assign _GEN_2474 = 11'h225 == RADDR ? 11'h225 : _GEN_2473; // @[RAM_ST.scala 32:46]
  assign _GEN_2475 = 11'h226 == RADDR ? 11'h226 : _GEN_2474; // @[RAM_ST.scala 32:46]
  assign _GEN_2476 = 11'h227 == RADDR ? 11'h227 : _GEN_2475; // @[RAM_ST.scala 32:46]
  assign _GEN_2477 = 11'h228 == RADDR ? 11'h228 : _GEN_2476; // @[RAM_ST.scala 32:46]
  assign _GEN_2478 = 11'h229 == RADDR ? 11'h229 : _GEN_2477; // @[RAM_ST.scala 32:46]
  assign _GEN_2479 = 11'h22a == RADDR ? 11'h22a : _GEN_2478; // @[RAM_ST.scala 32:46]
  assign _GEN_2480 = 11'h22b == RADDR ? 11'h22b : _GEN_2479; // @[RAM_ST.scala 32:46]
  assign _GEN_2481 = 11'h22c == RADDR ? 11'h22c : _GEN_2480; // @[RAM_ST.scala 32:46]
  assign _GEN_2482 = 11'h22d == RADDR ? 11'h22d : _GEN_2481; // @[RAM_ST.scala 32:46]
  assign _GEN_2483 = 11'h22e == RADDR ? 11'h22e : _GEN_2482; // @[RAM_ST.scala 32:46]
  assign _GEN_2484 = 11'h22f == RADDR ? 11'h22f : _GEN_2483; // @[RAM_ST.scala 32:46]
  assign _GEN_2485 = 11'h230 == RADDR ? 11'h230 : _GEN_2484; // @[RAM_ST.scala 32:46]
  assign _GEN_2486 = 11'h231 == RADDR ? 11'h231 : _GEN_2485; // @[RAM_ST.scala 32:46]
  assign _GEN_2487 = 11'h232 == RADDR ? 11'h232 : _GEN_2486; // @[RAM_ST.scala 32:46]
  assign _GEN_2488 = 11'h233 == RADDR ? 11'h233 : _GEN_2487; // @[RAM_ST.scala 32:46]
  assign _GEN_2489 = 11'h234 == RADDR ? 11'h234 : _GEN_2488; // @[RAM_ST.scala 32:46]
  assign _GEN_2490 = 11'h235 == RADDR ? 11'h235 : _GEN_2489; // @[RAM_ST.scala 32:46]
  assign _GEN_2491 = 11'h236 == RADDR ? 11'h236 : _GEN_2490; // @[RAM_ST.scala 32:46]
  assign _GEN_2492 = 11'h237 == RADDR ? 11'h237 : _GEN_2491; // @[RAM_ST.scala 32:46]
  assign _GEN_2493 = 11'h238 == RADDR ? 11'h238 : _GEN_2492; // @[RAM_ST.scala 32:46]
  assign _GEN_2494 = 11'h239 == RADDR ? 11'h239 : _GEN_2493; // @[RAM_ST.scala 32:46]
  assign _GEN_2495 = 11'h23a == RADDR ? 11'h23a : _GEN_2494; // @[RAM_ST.scala 32:46]
  assign _GEN_2496 = 11'h23b == RADDR ? 11'h23b : _GEN_2495; // @[RAM_ST.scala 32:46]
  assign _GEN_2497 = 11'h23c == RADDR ? 11'h23c : _GEN_2496; // @[RAM_ST.scala 32:46]
  assign _GEN_2498 = 11'h23d == RADDR ? 11'h23d : _GEN_2497; // @[RAM_ST.scala 32:46]
  assign _GEN_2499 = 11'h23e == RADDR ? 11'h23e : _GEN_2498; // @[RAM_ST.scala 32:46]
  assign _GEN_2500 = 11'h23f == RADDR ? 11'h23f : _GEN_2499; // @[RAM_ST.scala 32:46]
  assign _GEN_2501 = 11'h240 == RADDR ? 11'h240 : _GEN_2500; // @[RAM_ST.scala 32:46]
  assign _GEN_2502 = 11'h241 == RADDR ? 11'h241 : _GEN_2501; // @[RAM_ST.scala 32:46]
  assign _GEN_2503 = 11'h242 == RADDR ? 11'h242 : _GEN_2502; // @[RAM_ST.scala 32:46]
  assign _GEN_2504 = 11'h243 == RADDR ? 11'h243 : _GEN_2503; // @[RAM_ST.scala 32:46]
  assign _GEN_2505 = 11'h244 == RADDR ? 11'h244 : _GEN_2504; // @[RAM_ST.scala 32:46]
  assign _GEN_2506 = 11'h245 == RADDR ? 11'h245 : _GEN_2505; // @[RAM_ST.scala 32:46]
  assign _GEN_2507 = 11'h246 == RADDR ? 11'h246 : _GEN_2506; // @[RAM_ST.scala 32:46]
  assign _GEN_2508 = 11'h247 == RADDR ? 11'h247 : _GEN_2507; // @[RAM_ST.scala 32:46]
  assign _GEN_2509 = 11'h248 == RADDR ? 11'h248 : _GEN_2508; // @[RAM_ST.scala 32:46]
  assign _GEN_2510 = 11'h249 == RADDR ? 11'h249 : _GEN_2509; // @[RAM_ST.scala 32:46]
  assign _GEN_2511 = 11'h24a == RADDR ? 11'h24a : _GEN_2510; // @[RAM_ST.scala 32:46]
  assign _GEN_2512 = 11'h24b == RADDR ? 11'h24b : _GEN_2511; // @[RAM_ST.scala 32:46]
  assign _GEN_2513 = 11'h24c == RADDR ? 11'h24c : _GEN_2512; // @[RAM_ST.scala 32:46]
  assign _GEN_2514 = 11'h24d == RADDR ? 11'h24d : _GEN_2513; // @[RAM_ST.scala 32:46]
  assign _GEN_2515 = 11'h24e == RADDR ? 11'h24e : _GEN_2514; // @[RAM_ST.scala 32:46]
  assign _GEN_2516 = 11'h24f == RADDR ? 11'h24f : _GEN_2515; // @[RAM_ST.scala 32:46]
  assign _GEN_2517 = 11'h250 == RADDR ? 11'h250 : _GEN_2516; // @[RAM_ST.scala 32:46]
  assign _GEN_2518 = 11'h251 == RADDR ? 11'h251 : _GEN_2517; // @[RAM_ST.scala 32:46]
  assign _GEN_2519 = 11'h252 == RADDR ? 11'h252 : _GEN_2518; // @[RAM_ST.scala 32:46]
  assign _GEN_2520 = 11'h253 == RADDR ? 11'h253 : _GEN_2519; // @[RAM_ST.scala 32:46]
  assign _GEN_2521 = 11'h254 == RADDR ? 11'h254 : _GEN_2520; // @[RAM_ST.scala 32:46]
  assign _GEN_2522 = 11'h255 == RADDR ? 11'h255 : _GEN_2521; // @[RAM_ST.scala 32:46]
  assign _GEN_2523 = 11'h256 == RADDR ? 11'h256 : _GEN_2522; // @[RAM_ST.scala 32:46]
  assign _GEN_2524 = 11'h257 == RADDR ? 11'h257 : _GEN_2523; // @[RAM_ST.scala 32:46]
  assign _GEN_2525 = 11'h258 == RADDR ? 11'h258 : _GEN_2524; // @[RAM_ST.scala 32:46]
  assign _GEN_2526 = 11'h259 == RADDR ? 11'h259 : _GEN_2525; // @[RAM_ST.scala 32:46]
  assign _GEN_2527 = 11'h25a == RADDR ? 11'h25a : _GEN_2526; // @[RAM_ST.scala 32:46]
  assign _GEN_2528 = 11'h25b == RADDR ? 11'h25b : _GEN_2527; // @[RAM_ST.scala 32:46]
  assign _GEN_2529 = 11'h25c == RADDR ? 11'h25c : _GEN_2528; // @[RAM_ST.scala 32:46]
  assign _GEN_2530 = 11'h25d == RADDR ? 11'h25d : _GEN_2529; // @[RAM_ST.scala 32:46]
  assign _GEN_2531 = 11'h25e == RADDR ? 11'h25e : _GEN_2530; // @[RAM_ST.scala 32:46]
  assign _GEN_2532 = 11'h25f == RADDR ? 11'h25f : _GEN_2531; // @[RAM_ST.scala 32:46]
  assign _GEN_2533 = 11'h260 == RADDR ? 11'h260 : _GEN_2532; // @[RAM_ST.scala 32:46]
  assign _GEN_2534 = 11'h261 == RADDR ? 11'h261 : _GEN_2533; // @[RAM_ST.scala 32:46]
  assign _GEN_2535 = 11'h262 == RADDR ? 11'h262 : _GEN_2534; // @[RAM_ST.scala 32:46]
  assign _GEN_2536 = 11'h263 == RADDR ? 11'h263 : _GEN_2535; // @[RAM_ST.scala 32:46]
  assign _GEN_2537 = 11'h264 == RADDR ? 11'h264 : _GEN_2536; // @[RAM_ST.scala 32:46]
  assign _GEN_2538 = 11'h265 == RADDR ? 11'h265 : _GEN_2537; // @[RAM_ST.scala 32:46]
  assign _GEN_2539 = 11'h266 == RADDR ? 11'h266 : _GEN_2538; // @[RAM_ST.scala 32:46]
  assign _GEN_2540 = 11'h267 == RADDR ? 11'h267 : _GEN_2539; // @[RAM_ST.scala 32:46]
  assign _GEN_2541 = 11'h268 == RADDR ? 11'h268 : _GEN_2540; // @[RAM_ST.scala 32:46]
  assign _GEN_2542 = 11'h269 == RADDR ? 11'h269 : _GEN_2541; // @[RAM_ST.scala 32:46]
  assign _GEN_2543 = 11'h26a == RADDR ? 11'h26a : _GEN_2542; // @[RAM_ST.scala 32:46]
  assign _GEN_2544 = 11'h26b == RADDR ? 11'h26b : _GEN_2543; // @[RAM_ST.scala 32:46]
  assign _GEN_2545 = 11'h26c == RADDR ? 11'h26c : _GEN_2544; // @[RAM_ST.scala 32:46]
  assign _GEN_2546 = 11'h26d == RADDR ? 11'h26d : _GEN_2545; // @[RAM_ST.scala 32:46]
  assign _GEN_2547 = 11'h26e == RADDR ? 11'h26e : _GEN_2546; // @[RAM_ST.scala 32:46]
  assign _GEN_2548 = 11'h26f == RADDR ? 11'h26f : _GEN_2547; // @[RAM_ST.scala 32:46]
  assign _GEN_2549 = 11'h270 == RADDR ? 11'h270 : _GEN_2548; // @[RAM_ST.scala 32:46]
  assign _GEN_2550 = 11'h271 == RADDR ? 11'h271 : _GEN_2549; // @[RAM_ST.scala 32:46]
  assign _GEN_2551 = 11'h272 == RADDR ? 11'h272 : _GEN_2550; // @[RAM_ST.scala 32:46]
  assign _GEN_2552 = 11'h273 == RADDR ? 11'h273 : _GEN_2551; // @[RAM_ST.scala 32:46]
  assign _GEN_2553 = 11'h274 == RADDR ? 11'h274 : _GEN_2552; // @[RAM_ST.scala 32:46]
  assign _GEN_2554 = 11'h275 == RADDR ? 11'h275 : _GEN_2553; // @[RAM_ST.scala 32:46]
  assign _GEN_2555 = 11'h276 == RADDR ? 11'h276 : _GEN_2554; // @[RAM_ST.scala 32:46]
  assign _GEN_2556 = 11'h277 == RADDR ? 11'h277 : _GEN_2555; // @[RAM_ST.scala 32:46]
  assign _GEN_2557 = 11'h278 == RADDR ? 11'h278 : _GEN_2556; // @[RAM_ST.scala 32:46]
  assign _GEN_2558 = 11'h279 == RADDR ? 11'h279 : _GEN_2557; // @[RAM_ST.scala 32:46]
  assign _GEN_2559 = 11'h27a == RADDR ? 11'h27a : _GEN_2558; // @[RAM_ST.scala 32:46]
  assign _GEN_2560 = 11'h27b == RADDR ? 11'h27b : _GEN_2559; // @[RAM_ST.scala 32:46]
  assign _GEN_2561 = 11'h27c == RADDR ? 11'h27c : _GEN_2560; // @[RAM_ST.scala 32:46]
  assign _GEN_2562 = 11'h27d == RADDR ? 11'h27d : _GEN_2561; // @[RAM_ST.scala 32:46]
  assign _GEN_2563 = 11'h27e == RADDR ? 11'h27e : _GEN_2562; // @[RAM_ST.scala 32:46]
  assign _GEN_2564 = 11'h27f == RADDR ? 11'h27f : _GEN_2563; // @[RAM_ST.scala 32:46]
  assign _GEN_2565 = 11'h280 == RADDR ? 11'h280 : _GEN_2564; // @[RAM_ST.scala 32:46]
  assign _GEN_2566 = 11'h281 == RADDR ? 11'h281 : _GEN_2565; // @[RAM_ST.scala 32:46]
  assign _GEN_2567 = 11'h282 == RADDR ? 11'h282 : _GEN_2566; // @[RAM_ST.scala 32:46]
  assign _GEN_2568 = 11'h283 == RADDR ? 11'h283 : _GEN_2567; // @[RAM_ST.scala 32:46]
  assign _GEN_2569 = 11'h284 == RADDR ? 11'h284 : _GEN_2568; // @[RAM_ST.scala 32:46]
  assign _GEN_2570 = 11'h285 == RADDR ? 11'h285 : _GEN_2569; // @[RAM_ST.scala 32:46]
  assign _GEN_2571 = 11'h286 == RADDR ? 11'h286 : _GEN_2570; // @[RAM_ST.scala 32:46]
  assign _GEN_2572 = 11'h287 == RADDR ? 11'h287 : _GEN_2571; // @[RAM_ST.scala 32:46]
  assign _GEN_2573 = 11'h288 == RADDR ? 11'h288 : _GEN_2572; // @[RAM_ST.scala 32:46]
  assign _GEN_2574 = 11'h289 == RADDR ? 11'h289 : _GEN_2573; // @[RAM_ST.scala 32:46]
  assign _GEN_2575 = 11'h28a == RADDR ? 11'h28a : _GEN_2574; // @[RAM_ST.scala 32:46]
  assign _GEN_2576 = 11'h28b == RADDR ? 11'h28b : _GEN_2575; // @[RAM_ST.scala 32:46]
  assign _GEN_2577 = 11'h28c == RADDR ? 11'h28c : _GEN_2576; // @[RAM_ST.scala 32:46]
  assign _GEN_2578 = 11'h28d == RADDR ? 11'h28d : _GEN_2577; // @[RAM_ST.scala 32:46]
  assign _GEN_2579 = 11'h28e == RADDR ? 11'h28e : _GEN_2578; // @[RAM_ST.scala 32:46]
  assign _GEN_2580 = 11'h28f == RADDR ? 11'h28f : _GEN_2579; // @[RAM_ST.scala 32:46]
  assign _GEN_2581 = 11'h290 == RADDR ? 11'h290 : _GEN_2580; // @[RAM_ST.scala 32:46]
  assign _GEN_2582 = 11'h291 == RADDR ? 11'h291 : _GEN_2581; // @[RAM_ST.scala 32:46]
  assign _GEN_2583 = 11'h292 == RADDR ? 11'h292 : _GEN_2582; // @[RAM_ST.scala 32:46]
  assign _GEN_2584 = 11'h293 == RADDR ? 11'h293 : _GEN_2583; // @[RAM_ST.scala 32:46]
  assign _GEN_2585 = 11'h294 == RADDR ? 11'h294 : _GEN_2584; // @[RAM_ST.scala 32:46]
  assign _GEN_2586 = 11'h295 == RADDR ? 11'h295 : _GEN_2585; // @[RAM_ST.scala 32:46]
  assign _GEN_2587 = 11'h296 == RADDR ? 11'h296 : _GEN_2586; // @[RAM_ST.scala 32:46]
  assign _GEN_2588 = 11'h297 == RADDR ? 11'h297 : _GEN_2587; // @[RAM_ST.scala 32:46]
  assign _GEN_2589 = 11'h298 == RADDR ? 11'h298 : _GEN_2588; // @[RAM_ST.scala 32:46]
  assign _GEN_2590 = 11'h299 == RADDR ? 11'h299 : _GEN_2589; // @[RAM_ST.scala 32:46]
  assign _GEN_2591 = 11'h29a == RADDR ? 11'h29a : _GEN_2590; // @[RAM_ST.scala 32:46]
  assign _GEN_2592 = 11'h29b == RADDR ? 11'h29b : _GEN_2591; // @[RAM_ST.scala 32:46]
  assign _GEN_2593 = 11'h29c == RADDR ? 11'h29c : _GEN_2592; // @[RAM_ST.scala 32:46]
  assign _GEN_2594 = 11'h29d == RADDR ? 11'h29d : _GEN_2593; // @[RAM_ST.scala 32:46]
  assign _GEN_2595 = 11'h29e == RADDR ? 11'h29e : _GEN_2594; // @[RAM_ST.scala 32:46]
  assign _GEN_2596 = 11'h29f == RADDR ? 11'h29f : _GEN_2595; // @[RAM_ST.scala 32:46]
  assign _GEN_2597 = 11'h2a0 == RADDR ? 11'h2a0 : _GEN_2596; // @[RAM_ST.scala 32:46]
  assign _GEN_2598 = 11'h2a1 == RADDR ? 11'h2a1 : _GEN_2597; // @[RAM_ST.scala 32:46]
  assign _GEN_2599 = 11'h2a2 == RADDR ? 11'h2a2 : _GEN_2598; // @[RAM_ST.scala 32:46]
  assign _GEN_2600 = 11'h2a3 == RADDR ? 11'h2a3 : _GEN_2599; // @[RAM_ST.scala 32:46]
  assign _GEN_2601 = 11'h2a4 == RADDR ? 11'h2a4 : _GEN_2600; // @[RAM_ST.scala 32:46]
  assign _GEN_2602 = 11'h2a5 == RADDR ? 11'h2a5 : _GEN_2601; // @[RAM_ST.scala 32:46]
  assign _GEN_2603 = 11'h2a6 == RADDR ? 11'h2a6 : _GEN_2602; // @[RAM_ST.scala 32:46]
  assign _GEN_2604 = 11'h2a7 == RADDR ? 11'h2a7 : _GEN_2603; // @[RAM_ST.scala 32:46]
  assign _GEN_2605 = 11'h2a8 == RADDR ? 11'h2a8 : _GEN_2604; // @[RAM_ST.scala 32:46]
  assign _GEN_2606 = 11'h2a9 == RADDR ? 11'h2a9 : _GEN_2605; // @[RAM_ST.scala 32:46]
  assign _GEN_2607 = 11'h2aa == RADDR ? 11'h2aa : _GEN_2606; // @[RAM_ST.scala 32:46]
  assign _GEN_2608 = 11'h2ab == RADDR ? 11'h2ab : _GEN_2607; // @[RAM_ST.scala 32:46]
  assign _GEN_2609 = 11'h2ac == RADDR ? 11'h2ac : _GEN_2608; // @[RAM_ST.scala 32:46]
  assign _GEN_2610 = 11'h2ad == RADDR ? 11'h2ad : _GEN_2609; // @[RAM_ST.scala 32:46]
  assign _GEN_2611 = 11'h2ae == RADDR ? 11'h2ae : _GEN_2610; // @[RAM_ST.scala 32:46]
  assign _GEN_2612 = 11'h2af == RADDR ? 11'h2af : _GEN_2611; // @[RAM_ST.scala 32:46]
  assign _GEN_2613 = 11'h2b0 == RADDR ? 11'h2b0 : _GEN_2612; // @[RAM_ST.scala 32:46]
  assign _GEN_2614 = 11'h2b1 == RADDR ? 11'h2b1 : _GEN_2613; // @[RAM_ST.scala 32:46]
  assign _GEN_2615 = 11'h2b2 == RADDR ? 11'h2b2 : _GEN_2614; // @[RAM_ST.scala 32:46]
  assign _GEN_2616 = 11'h2b3 == RADDR ? 11'h2b3 : _GEN_2615; // @[RAM_ST.scala 32:46]
  assign _GEN_2617 = 11'h2b4 == RADDR ? 11'h2b4 : _GEN_2616; // @[RAM_ST.scala 32:46]
  assign _GEN_2618 = 11'h2b5 == RADDR ? 11'h2b5 : _GEN_2617; // @[RAM_ST.scala 32:46]
  assign _GEN_2619 = 11'h2b6 == RADDR ? 11'h2b6 : _GEN_2618; // @[RAM_ST.scala 32:46]
  assign _GEN_2620 = 11'h2b7 == RADDR ? 11'h2b7 : _GEN_2619; // @[RAM_ST.scala 32:46]
  assign _GEN_2621 = 11'h2b8 == RADDR ? 11'h2b8 : _GEN_2620; // @[RAM_ST.scala 32:46]
  assign _GEN_2622 = 11'h2b9 == RADDR ? 11'h2b9 : _GEN_2621; // @[RAM_ST.scala 32:46]
  assign _GEN_2623 = 11'h2ba == RADDR ? 11'h2ba : _GEN_2622; // @[RAM_ST.scala 32:46]
  assign _GEN_2624 = 11'h2bb == RADDR ? 11'h2bb : _GEN_2623; // @[RAM_ST.scala 32:46]
  assign _GEN_2625 = 11'h2bc == RADDR ? 11'h2bc : _GEN_2624; // @[RAM_ST.scala 32:46]
  assign _GEN_2626 = 11'h2bd == RADDR ? 11'h2bd : _GEN_2625; // @[RAM_ST.scala 32:46]
  assign _GEN_2627 = 11'h2be == RADDR ? 11'h2be : _GEN_2626; // @[RAM_ST.scala 32:46]
  assign _GEN_2628 = 11'h2bf == RADDR ? 11'h2bf : _GEN_2627; // @[RAM_ST.scala 32:46]
  assign _GEN_2629 = 11'h2c0 == RADDR ? 11'h2c0 : _GEN_2628; // @[RAM_ST.scala 32:46]
  assign _GEN_2630 = 11'h2c1 == RADDR ? 11'h2c1 : _GEN_2629; // @[RAM_ST.scala 32:46]
  assign _GEN_2631 = 11'h2c2 == RADDR ? 11'h2c2 : _GEN_2630; // @[RAM_ST.scala 32:46]
  assign _GEN_2632 = 11'h2c3 == RADDR ? 11'h2c3 : _GEN_2631; // @[RAM_ST.scala 32:46]
  assign _GEN_2633 = 11'h2c4 == RADDR ? 11'h2c4 : _GEN_2632; // @[RAM_ST.scala 32:46]
  assign _GEN_2634 = 11'h2c5 == RADDR ? 11'h2c5 : _GEN_2633; // @[RAM_ST.scala 32:46]
  assign _GEN_2635 = 11'h2c6 == RADDR ? 11'h2c6 : _GEN_2634; // @[RAM_ST.scala 32:46]
  assign _GEN_2636 = 11'h2c7 == RADDR ? 11'h2c7 : _GEN_2635; // @[RAM_ST.scala 32:46]
  assign _GEN_2637 = 11'h2c8 == RADDR ? 11'h2c8 : _GEN_2636; // @[RAM_ST.scala 32:46]
  assign _GEN_2638 = 11'h2c9 == RADDR ? 11'h2c9 : _GEN_2637; // @[RAM_ST.scala 32:46]
  assign _GEN_2639 = 11'h2ca == RADDR ? 11'h2ca : _GEN_2638; // @[RAM_ST.scala 32:46]
  assign _GEN_2640 = 11'h2cb == RADDR ? 11'h2cb : _GEN_2639; // @[RAM_ST.scala 32:46]
  assign _GEN_2641 = 11'h2cc == RADDR ? 11'h2cc : _GEN_2640; // @[RAM_ST.scala 32:46]
  assign _GEN_2642 = 11'h2cd == RADDR ? 11'h2cd : _GEN_2641; // @[RAM_ST.scala 32:46]
  assign _GEN_2643 = 11'h2ce == RADDR ? 11'h2ce : _GEN_2642; // @[RAM_ST.scala 32:46]
  assign _GEN_2644 = 11'h2cf == RADDR ? 11'h2cf : _GEN_2643; // @[RAM_ST.scala 32:46]
  assign _GEN_2645 = 11'h2d0 == RADDR ? 11'h2d0 : _GEN_2644; // @[RAM_ST.scala 32:46]
  assign _GEN_2646 = 11'h2d1 == RADDR ? 11'h2d1 : _GEN_2645; // @[RAM_ST.scala 32:46]
  assign _GEN_2647 = 11'h2d2 == RADDR ? 11'h2d2 : _GEN_2646; // @[RAM_ST.scala 32:46]
  assign _GEN_2648 = 11'h2d3 == RADDR ? 11'h2d3 : _GEN_2647; // @[RAM_ST.scala 32:46]
  assign _GEN_2649 = 11'h2d4 == RADDR ? 11'h2d4 : _GEN_2648; // @[RAM_ST.scala 32:46]
  assign _GEN_2650 = 11'h2d5 == RADDR ? 11'h2d5 : _GEN_2649; // @[RAM_ST.scala 32:46]
  assign _GEN_2651 = 11'h2d6 == RADDR ? 11'h2d6 : _GEN_2650; // @[RAM_ST.scala 32:46]
  assign _GEN_2652 = 11'h2d7 == RADDR ? 11'h2d7 : _GEN_2651; // @[RAM_ST.scala 32:46]
  assign _GEN_2653 = 11'h2d8 == RADDR ? 11'h2d8 : _GEN_2652; // @[RAM_ST.scala 32:46]
  assign _GEN_2654 = 11'h2d9 == RADDR ? 11'h2d9 : _GEN_2653; // @[RAM_ST.scala 32:46]
  assign _GEN_2655 = 11'h2da == RADDR ? 11'h2da : _GEN_2654; // @[RAM_ST.scala 32:46]
  assign _GEN_2656 = 11'h2db == RADDR ? 11'h2db : _GEN_2655; // @[RAM_ST.scala 32:46]
  assign _GEN_2657 = 11'h2dc == RADDR ? 11'h2dc : _GEN_2656; // @[RAM_ST.scala 32:46]
  assign _GEN_2658 = 11'h2dd == RADDR ? 11'h2dd : _GEN_2657; // @[RAM_ST.scala 32:46]
  assign _GEN_2659 = 11'h2de == RADDR ? 11'h2de : _GEN_2658; // @[RAM_ST.scala 32:46]
  assign _GEN_2660 = 11'h2df == RADDR ? 11'h2df : _GEN_2659; // @[RAM_ST.scala 32:46]
  assign _GEN_2661 = 11'h2e0 == RADDR ? 11'h2e0 : _GEN_2660; // @[RAM_ST.scala 32:46]
  assign _GEN_2662 = 11'h2e1 == RADDR ? 11'h2e1 : _GEN_2661; // @[RAM_ST.scala 32:46]
  assign _GEN_2663 = 11'h2e2 == RADDR ? 11'h2e2 : _GEN_2662; // @[RAM_ST.scala 32:46]
  assign _GEN_2664 = 11'h2e3 == RADDR ? 11'h2e3 : _GEN_2663; // @[RAM_ST.scala 32:46]
  assign _GEN_2665 = 11'h2e4 == RADDR ? 11'h2e4 : _GEN_2664; // @[RAM_ST.scala 32:46]
  assign _GEN_2666 = 11'h2e5 == RADDR ? 11'h2e5 : _GEN_2665; // @[RAM_ST.scala 32:46]
  assign _GEN_2667 = 11'h2e6 == RADDR ? 11'h2e6 : _GEN_2666; // @[RAM_ST.scala 32:46]
  assign _GEN_2668 = 11'h2e7 == RADDR ? 11'h2e7 : _GEN_2667; // @[RAM_ST.scala 32:46]
  assign _GEN_2669 = 11'h2e8 == RADDR ? 11'h2e8 : _GEN_2668; // @[RAM_ST.scala 32:46]
  assign _GEN_2670 = 11'h2e9 == RADDR ? 11'h2e9 : _GEN_2669; // @[RAM_ST.scala 32:46]
  assign _GEN_2671 = 11'h2ea == RADDR ? 11'h2ea : _GEN_2670; // @[RAM_ST.scala 32:46]
  assign _GEN_2672 = 11'h2eb == RADDR ? 11'h2eb : _GEN_2671; // @[RAM_ST.scala 32:46]
  assign _GEN_2673 = 11'h2ec == RADDR ? 11'h2ec : _GEN_2672; // @[RAM_ST.scala 32:46]
  assign _GEN_2674 = 11'h2ed == RADDR ? 11'h2ed : _GEN_2673; // @[RAM_ST.scala 32:46]
  assign _GEN_2675 = 11'h2ee == RADDR ? 11'h2ee : _GEN_2674; // @[RAM_ST.scala 32:46]
  assign _GEN_2676 = 11'h2ef == RADDR ? 11'h2ef : _GEN_2675; // @[RAM_ST.scala 32:46]
  assign _GEN_2677 = 11'h2f0 == RADDR ? 11'h2f0 : _GEN_2676; // @[RAM_ST.scala 32:46]
  assign _GEN_2678 = 11'h2f1 == RADDR ? 11'h2f1 : _GEN_2677; // @[RAM_ST.scala 32:46]
  assign _GEN_2679 = 11'h2f2 == RADDR ? 11'h2f2 : _GEN_2678; // @[RAM_ST.scala 32:46]
  assign _GEN_2680 = 11'h2f3 == RADDR ? 11'h2f3 : _GEN_2679; // @[RAM_ST.scala 32:46]
  assign _GEN_2681 = 11'h2f4 == RADDR ? 11'h2f4 : _GEN_2680; // @[RAM_ST.scala 32:46]
  assign _GEN_2682 = 11'h2f5 == RADDR ? 11'h2f5 : _GEN_2681; // @[RAM_ST.scala 32:46]
  assign _GEN_2683 = 11'h2f6 == RADDR ? 11'h2f6 : _GEN_2682; // @[RAM_ST.scala 32:46]
  assign _GEN_2684 = 11'h2f7 == RADDR ? 11'h2f7 : _GEN_2683; // @[RAM_ST.scala 32:46]
  assign _GEN_2685 = 11'h2f8 == RADDR ? 11'h2f8 : _GEN_2684; // @[RAM_ST.scala 32:46]
  assign _GEN_2686 = 11'h2f9 == RADDR ? 11'h2f9 : _GEN_2685; // @[RAM_ST.scala 32:46]
  assign _GEN_2687 = 11'h2fa == RADDR ? 11'h2fa : _GEN_2686; // @[RAM_ST.scala 32:46]
  assign _GEN_2688 = 11'h2fb == RADDR ? 11'h2fb : _GEN_2687; // @[RAM_ST.scala 32:46]
  assign _GEN_2689 = 11'h2fc == RADDR ? 11'h2fc : _GEN_2688; // @[RAM_ST.scala 32:46]
  assign _GEN_2690 = 11'h2fd == RADDR ? 11'h2fd : _GEN_2689; // @[RAM_ST.scala 32:46]
  assign _GEN_2691 = 11'h2fe == RADDR ? 11'h2fe : _GEN_2690; // @[RAM_ST.scala 32:46]
  assign _GEN_2692 = 11'h2ff == RADDR ? 11'h2ff : _GEN_2691; // @[RAM_ST.scala 32:46]
  assign _GEN_2693 = 11'h300 == RADDR ? 11'h300 : _GEN_2692; // @[RAM_ST.scala 32:46]
  assign _GEN_2694 = 11'h301 == RADDR ? 11'h301 : _GEN_2693; // @[RAM_ST.scala 32:46]
  assign _GEN_2695 = 11'h302 == RADDR ? 11'h302 : _GEN_2694; // @[RAM_ST.scala 32:46]
  assign _GEN_2696 = 11'h303 == RADDR ? 11'h303 : _GEN_2695; // @[RAM_ST.scala 32:46]
  assign _GEN_2697 = 11'h304 == RADDR ? 11'h304 : _GEN_2696; // @[RAM_ST.scala 32:46]
  assign _GEN_2698 = 11'h305 == RADDR ? 11'h305 : _GEN_2697; // @[RAM_ST.scala 32:46]
  assign _GEN_2699 = 11'h306 == RADDR ? 11'h306 : _GEN_2698; // @[RAM_ST.scala 32:46]
  assign _GEN_2700 = 11'h307 == RADDR ? 11'h307 : _GEN_2699; // @[RAM_ST.scala 32:46]
  assign _GEN_2701 = 11'h308 == RADDR ? 11'h308 : _GEN_2700; // @[RAM_ST.scala 32:46]
  assign _GEN_2702 = 11'h309 == RADDR ? 11'h309 : _GEN_2701; // @[RAM_ST.scala 32:46]
  assign _GEN_2703 = 11'h30a == RADDR ? 11'h30a : _GEN_2702; // @[RAM_ST.scala 32:46]
  assign _GEN_2704 = 11'h30b == RADDR ? 11'h30b : _GEN_2703; // @[RAM_ST.scala 32:46]
  assign _GEN_2705 = 11'h30c == RADDR ? 11'h30c : _GEN_2704; // @[RAM_ST.scala 32:46]
  assign _GEN_2706 = 11'h30d == RADDR ? 11'h30d : _GEN_2705; // @[RAM_ST.scala 32:46]
  assign _GEN_2707 = 11'h30e == RADDR ? 11'h30e : _GEN_2706; // @[RAM_ST.scala 32:46]
  assign _GEN_2708 = 11'h30f == RADDR ? 11'h30f : _GEN_2707; // @[RAM_ST.scala 32:46]
  assign _GEN_2709 = 11'h310 == RADDR ? 11'h310 : _GEN_2708; // @[RAM_ST.scala 32:46]
  assign _GEN_2710 = 11'h311 == RADDR ? 11'h311 : _GEN_2709; // @[RAM_ST.scala 32:46]
  assign _GEN_2711 = 11'h312 == RADDR ? 11'h312 : _GEN_2710; // @[RAM_ST.scala 32:46]
  assign _GEN_2712 = 11'h313 == RADDR ? 11'h313 : _GEN_2711; // @[RAM_ST.scala 32:46]
  assign _GEN_2713 = 11'h314 == RADDR ? 11'h314 : _GEN_2712; // @[RAM_ST.scala 32:46]
  assign _GEN_2714 = 11'h315 == RADDR ? 11'h315 : _GEN_2713; // @[RAM_ST.scala 32:46]
  assign _GEN_2715 = 11'h316 == RADDR ? 11'h316 : _GEN_2714; // @[RAM_ST.scala 32:46]
  assign _GEN_2716 = 11'h317 == RADDR ? 11'h317 : _GEN_2715; // @[RAM_ST.scala 32:46]
  assign _GEN_2717 = 11'h318 == RADDR ? 11'h318 : _GEN_2716; // @[RAM_ST.scala 32:46]
  assign _GEN_2718 = 11'h319 == RADDR ? 11'h319 : _GEN_2717; // @[RAM_ST.scala 32:46]
  assign _GEN_2719 = 11'h31a == RADDR ? 11'h31a : _GEN_2718; // @[RAM_ST.scala 32:46]
  assign _GEN_2720 = 11'h31b == RADDR ? 11'h31b : _GEN_2719; // @[RAM_ST.scala 32:46]
  assign _GEN_2721 = 11'h31c == RADDR ? 11'h31c : _GEN_2720; // @[RAM_ST.scala 32:46]
  assign _GEN_2722 = 11'h31d == RADDR ? 11'h31d : _GEN_2721; // @[RAM_ST.scala 32:46]
  assign _GEN_2723 = 11'h31e == RADDR ? 11'h31e : _GEN_2722; // @[RAM_ST.scala 32:46]
  assign _GEN_2724 = 11'h31f == RADDR ? 11'h31f : _GEN_2723; // @[RAM_ST.scala 32:46]
  assign _GEN_2725 = 11'h320 == RADDR ? 11'h320 : _GEN_2724; // @[RAM_ST.scala 32:46]
  assign _GEN_2726 = 11'h321 == RADDR ? 11'h321 : _GEN_2725; // @[RAM_ST.scala 32:46]
  assign _GEN_2727 = 11'h322 == RADDR ? 11'h322 : _GEN_2726; // @[RAM_ST.scala 32:46]
  assign _GEN_2728 = 11'h323 == RADDR ? 11'h323 : _GEN_2727; // @[RAM_ST.scala 32:46]
  assign _GEN_2729 = 11'h324 == RADDR ? 11'h324 : _GEN_2728; // @[RAM_ST.scala 32:46]
  assign _GEN_2730 = 11'h325 == RADDR ? 11'h325 : _GEN_2729; // @[RAM_ST.scala 32:46]
  assign _GEN_2731 = 11'h326 == RADDR ? 11'h326 : _GEN_2730; // @[RAM_ST.scala 32:46]
  assign _GEN_2732 = 11'h327 == RADDR ? 11'h327 : _GEN_2731; // @[RAM_ST.scala 32:46]
  assign _GEN_2733 = 11'h328 == RADDR ? 11'h328 : _GEN_2732; // @[RAM_ST.scala 32:46]
  assign _GEN_2734 = 11'h329 == RADDR ? 11'h329 : _GEN_2733; // @[RAM_ST.scala 32:46]
  assign _GEN_2735 = 11'h32a == RADDR ? 11'h32a : _GEN_2734; // @[RAM_ST.scala 32:46]
  assign _GEN_2736 = 11'h32b == RADDR ? 11'h32b : _GEN_2735; // @[RAM_ST.scala 32:46]
  assign _GEN_2737 = 11'h32c == RADDR ? 11'h32c : _GEN_2736; // @[RAM_ST.scala 32:46]
  assign _GEN_2738 = 11'h32d == RADDR ? 11'h32d : _GEN_2737; // @[RAM_ST.scala 32:46]
  assign _GEN_2739 = 11'h32e == RADDR ? 11'h32e : _GEN_2738; // @[RAM_ST.scala 32:46]
  assign _GEN_2740 = 11'h32f == RADDR ? 11'h32f : _GEN_2739; // @[RAM_ST.scala 32:46]
  assign _GEN_2741 = 11'h330 == RADDR ? 11'h330 : _GEN_2740; // @[RAM_ST.scala 32:46]
  assign _GEN_2742 = 11'h331 == RADDR ? 11'h331 : _GEN_2741; // @[RAM_ST.scala 32:46]
  assign _GEN_2743 = 11'h332 == RADDR ? 11'h332 : _GEN_2742; // @[RAM_ST.scala 32:46]
  assign _GEN_2744 = 11'h333 == RADDR ? 11'h333 : _GEN_2743; // @[RAM_ST.scala 32:46]
  assign _GEN_2745 = 11'h334 == RADDR ? 11'h334 : _GEN_2744; // @[RAM_ST.scala 32:46]
  assign _GEN_2746 = 11'h335 == RADDR ? 11'h335 : _GEN_2745; // @[RAM_ST.scala 32:46]
  assign _GEN_2747 = 11'h336 == RADDR ? 11'h336 : _GEN_2746; // @[RAM_ST.scala 32:46]
  assign _GEN_2748 = 11'h337 == RADDR ? 11'h337 : _GEN_2747; // @[RAM_ST.scala 32:46]
  assign _GEN_2749 = 11'h338 == RADDR ? 11'h338 : _GEN_2748; // @[RAM_ST.scala 32:46]
  assign _GEN_2750 = 11'h339 == RADDR ? 11'h339 : _GEN_2749; // @[RAM_ST.scala 32:46]
  assign _GEN_2751 = 11'h33a == RADDR ? 11'h33a : _GEN_2750; // @[RAM_ST.scala 32:46]
  assign _GEN_2752 = 11'h33b == RADDR ? 11'h33b : _GEN_2751; // @[RAM_ST.scala 32:46]
  assign _GEN_2753 = 11'h33c == RADDR ? 11'h33c : _GEN_2752; // @[RAM_ST.scala 32:46]
  assign _GEN_2754 = 11'h33d == RADDR ? 11'h33d : _GEN_2753; // @[RAM_ST.scala 32:46]
  assign _GEN_2755 = 11'h33e == RADDR ? 11'h33e : _GEN_2754; // @[RAM_ST.scala 32:46]
  assign _GEN_2756 = 11'h33f == RADDR ? 11'h33f : _GEN_2755; // @[RAM_ST.scala 32:46]
  assign _GEN_2757 = 11'h340 == RADDR ? 11'h340 : _GEN_2756; // @[RAM_ST.scala 32:46]
  assign _GEN_2758 = 11'h341 == RADDR ? 11'h341 : _GEN_2757; // @[RAM_ST.scala 32:46]
  assign _GEN_2759 = 11'h342 == RADDR ? 11'h342 : _GEN_2758; // @[RAM_ST.scala 32:46]
  assign _GEN_2760 = 11'h343 == RADDR ? 11'h343 : _GEN_2759; // @[RAM_ST.scala 32:46]
  assign _GEN_2761 = 11'h344 == RADDR ? 11'h344 : _GEN_2760; // @[RAM_ST.scala 32:46]
  assign _GEN_2762 = 11'h345 == RADDR ? 11'h345 : _GEN_2761; // @[RAM_ST.scala 32:46]
  assign _GEN_2763 = 11'h346 == RADDR ? 11'h346 : _GEN_2762; // @[RAM_ST.scala 32:46]
  assign _GEN_2764 = 11'h347 == RADDR ? 11'h347 : _GEN_2763; // @[RAM_ST.scala 32:46]
  assign _GEN_2765 = 11'h348 == RADDR ? 11'h348 : _GEN_2764; // @[RAM_ST.scala 32:46]
  assign _GEN_2766 = 11'h349 == RADDR ? 11'h349 : _GEN_2765; // @[RAM_ST.scala 32:46]
  assign _GEN_2767 = 11'h34a == RADDR ? 11'h34a : _GEN_2766; // @[RAM_ST.scala 32:46]
  assign _GEN_2768 = 11'h34b == RADDR ? 11'h34b : _GEN_2767; // @[RAM_ST.scala 32:46]
  assign _GEN_2769 = 11'h34c == RADDR ? 11'h34c : _GEN_2768; // @[RAM_ST.scala 32:46]
  assign _GEN_2770 = 11'h34d == RADDR ? 11'h34d : _GEN_2769; // @[RAM_ST.scala 32:46]
  assign _GEN_2771 = 11'h34e == RADDR ? 11'h34e : _GEN_2770; // @[RAM_ST.scala 32:46]
  assign _GEN_2772 = 11'h34f == RADDR ? 11'h34f : _GEN_2771; // @[RAM_ST.scala 32:46]
  assign _GEN_2773 = 11'h350 == RADDR ? 11'h350 : _GEN_2772; // @[RAM_ST.scala 32:46]
  assign _GEN_2774 = 11'h351 == RADDR ? 11'h351 : _GEN_2773; // @[RAM_ST.scala 32:46]
  assign _GEN_2775 = 11'h352 == RADDR ? 11'h352 : _GEN_2774; // @[RAM_ST.scala 32:46]
  assign _GEN_2776 = 11'h353 == RADDR ? 11'h353 : _GEN_2775; // @[RAM_ST.scala 32:46]
  assign _GEN_2777 = 11'h354 == RADDR ? 11'h354 : _GEN_2776; // @[RAM_ST.scala 32:46]
  assign _GEN_2778 = 11'h355 == RADDR ? 11'h355 : _GEN_2777; // @[RAM_ST.scala 32:46]
  assign _GEN_2779 = 11'h356 == RADDR ? 11'h356 : _GEN_2778; // @[RAM_ST.scala 32:46]
  assign _GEN_2780 = 11'h357 == RADDR ? 11'h357 : _GEN_2779; // @[RAM_ST.scala 32:46]
  assign _GEN_2781 = 11'h358 == RADDR ? 11'h358 : _GEN_2780; // @[RAM_ST.scala 32:46]
  assign _GEN_2782 = 11'h359 == RADDR ? 11'h359 : _GEN_2781; // @[RAM_ST.scala 32:46]
  assign _GEN_2783 = 11'h35a == RADDR ? 11'h35a : _GEN_2782; // @[RAM_ST.scala 32:46]
  assign _GEN_2784 = 11'h35b == RADDR ? 11'h35b : _GEN_2783; // @[RAM_ST.scala 32:46]
  assign _GEN_2785 = 11'h35c == RADDR ? 11'h35c : _GEN_2784; // @[RAM_ST.scala 32:46]
  assign _GEN_2786 = 11'h35d == RADDR ? 11'h35d : _GEN_2785; // @[RAM_ST.scala 32:46]
  assign _GEN_2787 = 11'h35e == RADDR ? 11'h35e : _GEN_2786; // @[RAM_ST.scala 32:46]
  assign _GEN_2788 = 11'h35f == RADDR ? 11'h35f : _GEN_2787; // @[RAM_ST.scala 32:46]
  assign _GEN_2789 = 11'h360 == RADDR ? 11'h360 : _GEN_2788; // @[RAM_ST.scala 32:46]
  assign _GEN_2790 = 11'h361 == RADDR ? 11'h361 : _GEN_2789; // @[RAM_ST.scala 32:46]
  assign _GEN_2791 = 11'h362 == RADDR ? 11'h362 : _GEN_2790; // @[RAM_ST.scala 32:46]
  assign _GEN_2792 = 11'h363 == RADDR ? 11'h363 : _GEN_2791; // @[RAM_ST.scala 32:46]
  assign _GEN_2793 = 11'h364 == RADDR ? 11'h364 : _GEN_2792; // @[RAM_ST.scala 32:46]
  assign _GEN_2794 = 11'h365 == RADDR ? 11'h365 : _GEN_2793; // @[RAM_ST.scala 32:46]
  assign _GEN_2795 = 11'h366 == RADDR ? 11'h366 : _GEN_2794; // @[RAM_ST.scala 32:46]
  assign _GEN_2796 = 11'h367 == RADDR ? 11'h367 : _GEN_2795; // @[RAM_ST.scala 32:46]
  assign _GEN_2797 = 11'h368 == RADDR ? 11'h368 : _GEN_2796; // @[RAM_ST.scala 32:46]
  assign _GEN_2798 = 11'h369 == RADDR ? 11'h369 : _GEN_2797; // @[RAM_ST.scala 32:46]
  assign _GEN_2799 = 11'h36a == RADDR ? 11'h36a : _GEN_2798; // @[RAM_ST.scala 32:46]
  assign _GEN_2800 = 11'h36b == RADDR ? 11'h36b : _GEN_2799; // @[RAM_ST.scala 32:46]
  assign _GEN_2801 = 11'h36c == RADDR ? 11'h36c : _GEN_2800; // @[RAM_ST.scala 32:46]
  assign _GEN_2802 = 11'h36d == RADDR ? 11'h36d : _GEN_2801; // @[RAM_ST.scala 32:46]
  assign _GEN_2803 = 11'h36e == RADDR ? 11'h36e : _GEN_2802; // @[RAM_ST.scala 32:46]
  assign _GEN_2804 = 11'h36f == RADDR ? 11'h36f : _GEN_2803; // @[RAM_ST.scala 32:46]
  assign _GEN_2805 = 11'h370 == RADDR ? 11'h370 : _GEN_2804; // @[RAM_ST.scala 32:46]
  assign _GEN_2806 = 11'h371 == RADDR ? 11'h371 : _GEN_2805; // @[RAM_ST.scala 32:46]
  assign _GEN_2807 = 11'h372 == RADDR ? 11'h372 : _GEN_2806; // @[RAM_ST.scala 32:46]
  assign _GEN_2808 = 11'h373 == RADDR ? 11'h373 : _GEN_2807; // @[RAM_ST.scala 32:46]
  assign _GEN_2809 = 11'h374 == RADDR ? 11'h374 : _GEN_2808; // @[RAM_ST.scala 32:46]
  assign _GEN_2810 = 11'h375 == RADDR ? 11'h375 : _GEN_2809; // @[RAM_ST.scala 32:46]
  assign _GEN_2811 = 11'h376 == RADDR ? 11'h376 : _GEN_2810; // @[RAM_ST.scala 32:46]
  assign _GEN_2812 = 11'h377 == RADDR ? 11'h377 : _GEN_2811; // @[RAM_ST.scala 32:46]
  assign _GEN_2813 = 11'h378 == RADDR ? 11'h378 : _GEN_2812; // @[RAM_ST.scala 32:46]
  assign _GEN_2814 = 11'h379 == RADDR ? 11'h379 : _GEN_2813; // @[RAM_ST.scala 32:46]
  assign _GEN_2815 = 11'h37a == RADDR ? 11'h37a : _GEN_2814; // @[RAM_ST.scala 32:46]
  assign _GEN_2816 = 11'h37b == RADDR ? 11'h37b : _GEN_2815; // @[RAM_ST.scala 32:46]
  assign _GEN_2817 = 11'h37c == RADDR ? 11'h37c : _GEN_2816; // @[RAM_ST.scala 32:46]
  assign _GEN_2818 = 11'h37d == RADDR ? 11'h37d : _GEN_2817; // @[RAM_ST.scala 32:46]
  assign _GEN_2819 = 11'h37e == RADDR ? 11'h37e : _GEN_2818; // @[RAM_ST.scala 32:46]
  assign _GEN_2820 = 11'h37f == RADDR ? 11'h37f : _GEN_2819; // @[RAM_ST.scala 32:46]
  assign _GEN_2821 = 11'h380 == RADDR ? 11'h380 : _GEN_2820; // @[RAM_ST.scala 32:46]
  assign _GEN_2822 = 11'h381 == RADDR ? 11'h381 : _GEN_2821; // @[RAM_ST.scala 32:46]
  assign _GEN_2823 = 11'h382 == RADDR ? 11'h382 : _GEN_2822; // @[RAM_ST.scala 32:46]
  assign _GEN_2824 = 11'h383 == RADDR ? 11'h383 : _GEN_2823; // @[RAM_ST.scala 32:46]
  assign _GEN_2825 = 11'h384 == RADDR ? 11'h384 : _GEN_2824; // @[RAM_ST.scala 32:46]
  assign _GEN_2826 = 11'h385 == RADDR ? 11'h385 : _GEN_2825; // @[RAM_ST.scala 32:46]
  assign _GEN_2827 = 11'h386 == RADDR ? 11'h386 : _GEN_2826; // @[RAM_ST.scala 32:46]
  assign _GEN_2828 = 11'h387 == RADDR ? 11'h387 : _GEN_2827; // @[RAM_ST.scala 32:46]
  assign _GEN_2829 = 11'h388 == RADDR ? 11'h388 : _GEN_2828; // @[RAM_ST.scala 32:46]
  assign _GEN_2830 = 11'h389 == RADDR ? 11'h389 : _GEN_2829; // @[RAM_ST.scala 32:46]
  assign _GEN_2831 = 11'h38a == RADDR ? 11'h38a : _GEN_2830; // @[RAM_ST.scala 32:46]
  assign _GEN_2832 = 11'h38b == RADDR ? 11'h38b : _GEN_2831; // @[RAM_ST.scala 32:46]
  assign _GEN_2833 = 11'h38c == RADDR ? 11'h38c : _GEN_2832; // @[RAM_ST.scala 32:46]
  assign _GEN_2834 = 11'h38d == RADDR ? 11'h38d : _GEN_2833; // @[RAM_ST.scala 32:46]
  assign _GEN_2835 = 11'h38e == RADDR ? 11'h38e : _GEN_2834; // @[RAM_ST.scala 32:46]
  assign _GEN_2836 = 11'h38f == RADDR ? 11'h38f : _GEN_2835; // @[RAM_ST.scala 32:46]
  assign _GEN_2837 = 11'h390 == RADDR ? 11'h390 : _GEN_2836; // @[RAM_ST.scala 32:46]
  assign _GEN_2838 = 11'h391 == RADDR ? 11'h391 : _GEN_2837; // @[RAM_ST.scala 32:46]
  assign _GEN_2839 = 11'h392 == RADDR ? 11'h392 : _GEN_2838; // @[RAM_ST.scala 32:46]
  assign _GEN_2840 = 11'h393 == RADDR ? 11'h393 : _GEN_2839; // @[RAM_ST.scala 32:46]
  assign _GEN_2841 = 11'h394 == RADDR ? 11'h394 : _GEN_2840; // @[RAM_ST.scala 32:46]
  assign _GEN_2842 = 11'h395 == RADDR ? 11'h395 : _GEN_2841; // @[RAM_ST.scala 32:46]
  assign _GEN_2843 = 11'h396 == RADDR ? 11'h396 : _GEN_2842; // @[RAM_ST.scala 32:46]
  assign _GEN_2844 = 11'h397 == RADDR ? 11'h397 : _GEN_2843; // @[RAM_ST.scala 32:46]
  assign _GEN_2845 = 11'h398 == RADDR ? 11'h398 : _GEN_2844; // @[RAM_ST.scala 32:46]
  assign _GEN_2846 = 11'h399 == RADDR ? 11'h399 : _GEN_2845; // @[RAM_ST.scala 32:46]
  assign _GEN_2847 = 11'h39a == RADDR ? 11'h39a : _GEN_2846; // @[RAM_ST.scala 32:46]
  assign _GEN_2848 = 11'h39b == RADDR ? 11'h39b : _GEN_2847; // @[RAM_ST.scala 32:46]
  assign _GEN_2849 = 11'h39c == RADDR ? 11'h39c : _GEN_2848; // @[RAM_ST.scala 32:46]
  assign _GEN_2850 = 11'h39d == RADDR ? 11'h39d : _GEN_2849; // @[RAM_ST.scala 32:46]
  assign _GEN_2851 = 11'h39e == RADDR ? 11'h39e : _GEN_2850; // @[RAM_ST.scala 32:46]
  assign _GEN_2852 = 11'h39f == RADDR ? 11'h39f : _GEN_2851; // @[RAM_ST.scala 32:46]
  assign _GEN_2853 = 11'h3a0 == RADDR ? 11'h3a0 : _GEN_2852; // @[RAM_ST.scala 32:46]
  assign _GEN_2854 = 11'h3a1 == RADDR ? 11'h3a1 : _GEN_2853; // @[RAM_ST.scala 32:46]
  assign _GEN_2855 = 11'h3a2 == RADDR ? 11'h3a2 : _GEN_2854; // @[RAM_ST.scala 32:46]
  assign _GEN_2856 = 11'h3a3 == RADDR ? 11'h3a3 : _GEN_2855; // @[RAM_ST.scala 32:46]
  assign _GEN_2857 = 11'h3a4 == RADDR ? 11'h3a4 : _GEN_2856; // @[RAM_ST.scala 32:46]
  assign _GEN_2858 = 11'h3a5 == RADDR ? 11'h3a5 : _GEN_2857; // @[RAM_ST.scala 32:46]
  assign _GEN_2859 = 11'h3a6 == RADDR ? 11'h3a6 : _GEN_2858; // @[RAM_ST.scala 32:46]
  assign _GEN_2860 = 11'h3a7 == RADDR ? 11'h3a7 : _GEN_2859; // @[RAM_ST.scala 32:46]
  assign _GEN_2861 = 11'h3a8 == RADDR ? 11'h3a8 : _GEN_2860; // @[RAM_ST.scala 32:46]
  assign _GEN_2862 = 11'h3a9 == RADDR ? 11'h3a9 : _GEN_2861; // @[RAM_ST.scala 32:46]
  assign _GEN_2863 = 11'h3aa == RADDR ? 11'h3aa : _GEN_2862; // @[RAM_ST.scala 32:46]
  assign _GEN_2864 = 11'h3ab == RADDR ? 11'h3ab : _GEN_2863; // @[RAM_ST.scala 32:46]
  assign _GEN_2865 = 11'h3ac == RADDR ? 11'h3ac : _GEN_2864; // @[RAM_ST.scala 32:46]
  assign _GEN_2866 = 11'h3ad == RADDR ? 11'h3ad : _GEN_2865; // @[RAM_ST.scala 32:46]
  assign _GEN_2867 = 11'h3ae == RADDR ? 11'h3ae : _GEN_2866; // @[RAM_ST.scala 32:46]
  assign _GEN_2868 = 11'h3af == RADDR ? 11'h3af : _GEN_2867; // @[RAM_ST.scala 32:46]
  assign _GEN_2869 = 11'h3b0 == RADDR ? 11'h3b0 : _GEN_2868; // @[RAM_ST.scala 32:46]
  assign _GEN_2870 = 11'h3b1 == RADDR ? 11'h3b1 : _GEN_2869; // @[RAM_ST.scala 32:46]
  assign _GEN_2871 = 11'h3b2 == RADDR ? 11'h3b2 : _GEN_2870; // @[RAM_ST.scala 32:46]
  assign _GEN_2872 = 11'h3b3 == RADDR ? 11'h3b3 : _GEN_2871; // @[RAM_ST.scala 32:46]
  assign _GEN_2873 = 11'h3b4 == RADDR ? 11'h3b4 : _GEN_2872; // @[RAM_ST.scala 32:46]
  assign _GEN_2874 = 11'h3b5 == RADDR ? 11'h3b5 : _GEN_2873; // @[RAM_ST.scala 32:46]
  assign _GEN_2875 = 11'h3b6 == RADDR ? 11'h3b6 : _GEN_2874; // @[RAM_ST.scala 32:46]
  assign _GEN_2876 = 11'h3b7 == RADDR ? 11'h3b7 : _GEN_2875; // @[RAM_ST.scala 32:46]
  assign _GEN_2877 = 11'h3b8 == RADDR ? 11'h3b8 : _GEN_2876; // @[RAM_ST.scala 32:46]
  assign _GEN_2878 = 11'h3b9 == RADDR ? 11'h3b9 : _GEN_2877; // @[RAM_ST.scala 32:46]
  assign _GEN_2879 = 11'h3ba == RADDR ? 11'h3ba : _GEN_2878; // @[RAM_ST.scala 32:46]
  assign _GEN_2880 = 11'h3bb == RADDR ? 11'h3bb : _GEN_2879; // @[RAM_ST.scala 32:46]
  assign _GEN_2881 = 11'h3bc == RADDR ? 11'h3bc : _GEN_2880; // @[RAM_ST.scala 32:46]
  assign _GEN_2882 = 11'h3bd == RADDR ? 11'h3bd : _GEN_2881; // @[RAM_ST.scala 32:46]
  assign _GEN_2883 = 11'h3be == RADDR ? 11'h3be : _GEN_2882; // @[RAM_ST.scala 32:46]
  assign _GEN_2884 = 11'h3bf == RADDR ? 11'h3bf : _GEN_2883; // @[RAM_ST.scala 32:46]
  assign _GEN_2885 = 11'h3c0 == RADDR ? 11'h3c0 : _GEN_2884; // @[RAM_ST.scala 32:46]
  assign _GEN_2886 = 11'h3c1 == RADDR ? 11'h3c1 : _GEN_2885; // @[RAM_ST.scala 32:46]
  assign _GEN_2887 = 11'h3c2 == RADDR ? 11'h3c2 : _GEN_2886; // @[RAM_ST.scala 32:46]
  assign _GEN_2888 = 11'h3c3 == RADDR ? 11'h3c3 : _GEN_2887; // @[RAM_ST.scala 32:46]
  assign _GEN_2889 = 11'h3c4 == RADDR ? 11'h3c4 : _GEN_2888; // @[RAM_ST.scala 32:46]
  assign _GEN_2890 = 11'h3c5 == RADDR ? 11'h3c5 : _GEN_2889; // @[RAM_ST.scala 32:46]
  assign _GEN_2891 = 11'h3c6 == RADDR ? 11'h3c6 : _GEN_2890; // @[RAM_ST.scala 32:46]
  assign _GEN_2892 = 11'h3c7 == RADDR ? 11'h3c7 : _GEN_2891; // @[RAM_ST.scala 32:46]
  assign _GEN_2893 = 11'h3c8 == RADDR ? 11'h3c8 : _GEN_2892; // @[RAM_ST.scala 32:46]
  assign _GEN_2894 = 11'h3c9 == RADDR ? 11'h3c9 : _GEN_2893; // @[RAM_ST.scala 32:46]
  assign _GEN_2895 = 11'h3ca == RADDR ? 11'h3ca : _GEN_2894; // @[RAM_ST.scala 32:46]
  assign _GEN_2896 = 11'h3cb == RADDR ? 11'h3cb : _GEN_2895; // @[RAM_ST.scala 32:46]
  assign _GEN_2897 = 11'h3cc == RADDR ? 11'h3cc : _GEN_2896; // @[RAM_ST.scala 32:46]
  assign _GEN_2898 = 11'h3cd == RADDR ? 11'h3cd : _GEN_2897; // @[RAM_ST.scala 32:46]
  assign _GEN_2899 = 11'h3ce == RADDR ? 11'h3ce : _GEN_2898; // @[RAM_ST.scala 32:46]
  assign _GEN_2900 = 11'h3cf == RADDR ? 11'h3cf : _GEN_2899; // @[RAM_ST.scala 32:46]
  assign _GEN_2901 = 11'h3d0 == RADDR ? 11'h3d0 : _GEN_2900; // @[RAM_ST.scala 32:46]
  assign _GEN_2902 = 11'h3d1 == RADDR ? 11'h3d1 : _GEN_2901; // @[RAM_ST.scala 32:46]
  assign _GEN_2903 = 11'h3d2 == RADDR ? 11'h3d2 : _GEN_2902; // @[RAM_ST.scala 32:46]
  assign _GEN_2904 = 11'h3d3 == RADDR ? 11'h3d3 : _GEN_2903; // @[RAM_ST.scala 32:46]
  assign _GEN_2905 = 11'h3d4 == RADDR ? 11'h3d4 : _GEN_2904; // @[RAM_ST.scala 32:46]
  assign _GEN_2906 = 11'h3d5 == RADDR ? 11'h3d5 : _GEN_2905; // @[RAM_ST.scala 32:46]
  assign _GEN_2907 = 11'h3d6 == RADDR ? 11'h3d6 : _GEN_2906; // @[RAM_ST.scala 32:46]
  assign _GEN_2908 = 11'h3d7 == RADDR ? 11'h3d7 : _GEN_2907; // @[RAM_ST.scala 32:46]
  assign _GEN_2909 = 11'h3d8 == RADDR ? 11'h3d8 : _GEN_2908; // @[RAM_ST.scala 32:46]
  assign _GEN_2910 = 11'h3d9 == RADDR ? 11'h3d9 : _GEN_2909; // @[RAM_ST.scala 32:46]
  assign _GEN_2911 = 11'h3da == RADDR ? 11'h3da : _GEN_2910; // @[RAM_ST.scala 32:46]
  assign _GEN_2912 = 11'h3db == RADDR ? 11'h3db : _GEN_2911; // @[RAM_ST.scala 32:46]
  assign _GEN_2913 = 11'h3dc == RADDR ? 11'h3dc : _GEN_2912; // @[RAM_ST.scala 32:46]
  assign _GEN_2914 = 11'h3dd == RADDR ? 11'h3dd : _GEN_2913; // @[RAM_ST.scala 32:46]
  assign _GEN_2915 = 11'h3de == RADDR ? 11'h3de : _GEN_2914; // @[RAM_ST.scala 32:46]
  assign _GEN_2916 = 11'h3df == RADDR ? 11'h3df : _GEN_2915; // @[RAM_ST.scala 32:46]
  assign _GEN_2917 = 11'h3e0 == RADDR ? 11'h3e0 : _GEN_2916; // @[RAM_ST.scala 32:46]
  assign _GEN_2918 = 11'h3e1 == RADDR ? 11'h3e1 : _GEN_2917; // @[RAM_ST.scala 32:46]
  assign _GEN_2919 = 11'h3e2 == RADDR ? 11'h3e2 : _GEN_2918; // @[RAM_ST.scala 32:46]
  assign _GEN_2920 = 11'h3e3 == RADDR ? 11'h3e3 : _GEN_2919; // @[RAM_ST.scala 32:46]
  assign _GEN_2921 = 11'h3e4 == RADDR ? 11'h3e4 : _GEN_2920; // @[RAM_ST.scala 32:46]
  assign _GEN_2922 = 11'h3e5 == RADDR ? 11'h3e5 : _GEN_2921; // @[RAM_ST.scala 32:46]
  assign _GEN_2923 = 11'h3e6 == RADDR ? 11'h3e6 : _GEN_2922; // @[RAM_ST.scala 32:46]
  assign _GEN_2924 = 11'h3e7 == RADDR ? 11'h3e7 : _GEN_2923; // @[RAM_ST.scala 32:46]
  assign _GEN_2925 = 11'h3e8 == RADDR ? 11'h3e8 : _GEN_2924; // @[RAM_ST.scala 32:46]
  assign _GEN_2926 = 11'h3e9 == RADDR ? 11'h3e9 : _GEN_2925; // @[RAM_ST.scala 32:46]
  assign _GEN_2927 = 11'h3ea == RADDR ? 11'h3ea : _GEN_2926; // @[RAM_ST.scala 32:46]
  assign _GEN_2928 = 11'h3eb == RADDR ? 11'h3eb : _GEN_2927; // @[RAM_ST.scala 32:46]
  assign _GEN_2929 = 11'h3ec == RADDR ? 11'h3ec : _GEN_2928; // @[RAM_ST.scala 32:46]
  assign _GEN_2930 = 11'h3ed == RADDR ? 11'h3ed : _GEN_2929; // @[RAM_ST.scala 32:46]
  assign _GEN_2931 = 11'h3ee == RADDR ? 11'h3ee : _GEN_2930; // @[RAM_ST.scala 32:46]
  assign _GEN_2932 = 11'h3ef == RADDR ? 11'h3ef : _GEN_2931; // @[RAM_ST.scala 32:46]
  assign _GEN_2933 = 11'h3f0 == RADDR ? 11'h3f0 : _GEN_2932; // @[RAM_ST.scala 32:46]
  assign _GEN_2934 = 11'h3f1 == RADDR ? 11'h3f1 : _GEN_2933; // @[RAM_ST.scala 32:46]
  assign _GEN_2935 = 11'h3f2 == RADDR ? 11'h3f2 : _GEN_2934; // @[RAM_ST.scala 32:46]
  assign _GEN_2936 = 11'h3f3 == RADDR ? 11'h3f3 : _GEN_2935; // @[RAM_ST.scala 32:46]
  assign _GEN_2937 = 11'h3f4 == RADDR ? 11'h3f4 : _GEN_2936; // @[RAM_ST.scala 32:46]
  assign _GEN_2938 = 11'h3f5 == RADDR ? 11'h3f5 : _GEN_2937; // @[RAM_ST.scala 32:46]
  assign _GEN_2939 = 11'h3f6 == RADDR ? 11'h3f6 : _GEN_2938; // @[RAM_ST.scala 32:46]
  assign _GEN_2940 = 11'h3f7 == RADDR ? 11'h3f7 : _GEN_2939; // @[RAM_ST.scala 32:46]
  assign _GEN_2941 = 11'h3f8 == RADDR ? 11'h3f8 : _GEN_2940; // @[RAM_ST.scala 32:46]
  assign _GEN_2942 = 11'h3f9 == RADDR ? 11'h3f9 : _GEN_2941; // @[RAM_ST.scala 32:46]
  assign _GEN_2943 = 11'h3fa == RADDR ? 11'h3fa : _GEN_2942; // @[RAM_ST.scala 32:46]
  assign _GEN_2944 = 11'h3fb == RADDR ? 11'h3fb : _GEN_2943; // @[RAM_ST.scala 32:46]
  assign _GEN_2945 = 11'h3fc == RADDR ? 11'h3fc : _GEN_2944; // @[RAM_ST.scala 32:46]
  assign _GEN_2946 = 11'h3fd == RADDR ? 11'h3fd : _GEN_2945; // @[RAM_ST.scala 32:46]
  assign _GEN_2947 = 11'h3fe == RADDR ? 11'h3fe : _GEN_2946; // @[RAM_ST.scala 32:46]
  assign _GEN_2948 = 11'h3ff == RADDR ? 11'h3ff : _GEN_2947; // @[RAM_ST.scala 32:46]
  assign _GEN_2949 = 11'h400 == RADDR ? 11'h400 : _GEN_2948; // @[RAM_ST.scala 32:46]
  assign _GEN_2950 = 11'h401 == RADDR ? 11'h401 : _GEN_2949; // @[RAM_ST.scala 32:46]
  assign _GEN_2951 = 11'h402 == RADDR ? 11'h402 : _GEN_2950; // @[RAM_ST.scala 32:46]
  assign _GEN_2952 = 11'h403 == RADDR ? 11'h403 : _GEN_2951; // @[RAM_ST.scala 32:46]
  assign _GEN_2953 = 11'h404 == RADDR ? 11'h404 : _GEN_2952; // @[RAM_ST.scala 32:46]
  assign _GEN_2954 = 11'h405 == RADDR ? 11'h405 : _GEN_2953; // @[RAM_ST.scala 32:46]
  assign _GEN_2955 = 11'h406 == RADDR ? 11'h406 : _GEN_2954; // @[RAM_ST.scala 32:46]
  assign _GEN_2956 = 11'h407 == RADDR ? 11'h407 : _GEN_2955; // @[RAM_ST.scala 32:46]
  assign _GEN_2957 = 11'h408 == RADDR ? 11'h408 : _GEN_2956; // @[RAM_ST.scala 32:46]
  assign _GEN_2958 = 11'h409 == RADDR ? 11'h409 : _GEN_2957; // @[RAM_ST.scala 32:46]
  assign _GEN_2959 = 11'h40a == RADDR ? 11'h40a : _GEN_2958; // @[RAM_ST.scala 32:46]
  assign _GEN_2960 = 11'h40b == RADDR ? 11'h40b : _GEN_2959; // @[RAM_ST.scala 32:46]
  assign _GEN_2961 = 11'h40c == RADDR ? 11'h40c : _GEN_2960; // @[RAM_ST.scala 32:46]
  assign _GEN_2962 = 11'h40d == RADDR ? 11'h40d : _GEN_2961; // @[RAM_ST.scala 32:46]
  assign _GEN_2963 = 11'h40e == RADDR ? 11'h40e : _GEN_2962; // @[RAM_ST.scala 32:46]
  assign _GEN_2964 = 11'h40f == RADDR ? 11'h40f : _GEN_2963; // @[RAM_ST.scala 32:46]
  assign _GEN_2965 = 11'h410 == RADDR ? 11'h410 : _GEN_2964; // @[RAM_ST.scala 32:46]
  assign _GEN_2966 = 11'h411 == RADDR ? 11'h411 : _GEN_2965; // @[RAM_ST.scala 32:46]
  assign _GEN_2967 = 11'h412 == RADDR ? 11'h412 : _GEN_2966; // @[RAM_ST.scala 32:46]
  assign _GEN_2968 = 11'h413 == RADDR ? 11'h413 : _GEN_2967; // @[RAM_ST.scala 32:46]
  assign _GEN_2969 = 11'h414 == RADDR ? 11'h414 : _GEN_2968; // @[RAM_ST.scala 32:46]
  assign _GEN_2970 = 11'h415 == RADDR ? 11'h415 : _GEN_2969; // @[RAM_ST.scala 32:46]
  assign _GEN_2971 = 11'h416 == RADDR ? 11'h416 : _GEN_2970; // @[RAM_ST.scala 32:46]
  assign _GEN_2972 = 11'h417 == RADDR ? 11'h417 : _GEN_2971; // @[RAM_ST.scala 32:46]
  assign _GEN_2973 = 11'h418 == RADDR ? 11'h418 : _GEN_2972; // @[RAM_ST.scala 32:46]
  assign _GEN_2974 = 11'h419 == RADDR ? 11'h419 : _GEN_2973; // @[RAM_ST.scala 32:46]
  assign _GEN_2975 = 11'h41a == RADDR ? 11'h41a : _GEN_2974; // @[RAM_ST.scala 32:46]
  assign _GEN_2976 = 11'h41b == RADDR ? 11'h41b : _GEN_2975; // @[RAM_ST.scala 32:46]
  assign _GEN_2977 = 11'h41c == RADDR ? 11'h41c : _GEN_2976; // @[RAM_ST.scala 32:46]
  assign _GEN_2978 = 11'h41d == RADDR ? 11'h41d : _GEN_2977; // @[RAM_ST.scala 32:46]
  assign _GEN_2979 = 11'h41e == RADDR ? 11'h41e : _GEN_2978; // @[RAM_ST.scala 32:46]
  assign _GEN_2980 = 11'h41f == RADDR ? 11'h41f : _GEN_2979; // @[RAM_ST.scala 32:46]
  assign _GEN_2981 = 11'h420 == RADDR ? 11'h420 : _GEN_2980; // @[RAM_ST.scala 32:46]
  assign _GEN_2982 = 11'h421 == RADDR ? 11'h421 : _GEN_2981; // @[RAM_ST.scala 32:46]
  assign _GEN_2983 = 11'h422 == RADDR ? 11'h422 : _GEN_2982; // @[RAM_ST.scala 32:46]
  assign _GEN_2984 = 11'h423 == RADDR ? 11'h423 : _GEN_2983; // @[RAM_ST.scala 32:46]
  assign _GEN_2985 = 11'h424 == RADDR ? 11'h424 : _GEN_2984; // @[RAM_ST.scala 32:46]
  assign _GEN_2986 = 11'h425 == RADDR ? 11'h425 : _GEN_2985; // @[RAM_ST.scala 32:46]
  assign _GEN_2987 = 11'h426 == RADDR ? 11'h426 : _GEN_2986; // @[RAM_ST.scala 32:46]
  assign _GEN_2988 = 11'h427 == RADDR ? 11'h427 : _GEN_2987; // @[RAM_ST.scala 32:46]
  assign _GEN_2989 = 11'h428 == RADDR ? 11'h428 : _GEN_2988; // @[RAM_ST.scala 32:46]
  assign _GEN_2990 = 11'h429 == RADDR ? 11'h429 : _GEN_2989; // @[RAM_ST.scala 32:46]
  assign _GEN_2991 = 11'h42a == RADDR ? 11'h42a : _GEN_2990; // @[RAM_ST.scala 32:46]
  assign _GEN_2992 = 11'h42b == RADDR ? 11'h42b : _GEN_2991; // @[RAM_ST.scala 32:46]
  assign _GEN_2993 = 11'h42c == RADDR ? 11'h42c : _GEN_2992; // @[RAM_ST.scala 32:46]
  assign _GEN_2994 = 11'h42d == RADDR ? 11'h42d : _GEN_2993; // @[RAM_ST.scala 32:46]
  assign _GEN_2995 = 11'h42e == RADDR ? 11'h42e : _GEN_2994; // @[RAM_ST.scala 32:46]
  assign _GEN_2996 = 11'h42f == RADDR ? 11'h42f : _GEN_2995; // @[RAM_ST.scala 32:46]
  assign _GEN_2997 = 11'h430 == RADDR ? 11'h430 : _GEN_2996; // @[RAM_ST.scala 32:46]
  assign _GEN_2998 = 11'h431 == RADDR ? 11'h431 : _GEN_2997; // @[RAM_ST.scala 32:46]
  assign _GEN_2999 = 11'h432 == RADDR ? 11'h432 : _GEN_2998; // @[RAM_ST.scala 32:46]
  assign _GEN_3000 = 11'h433 == RADDR ? 11'h433 : _GEN_2999; // @[RAM_ST.scala 32:46]
  assign _GEN_3001 = 11'h434 == RADDR ? 11'h434 : _GEN_3000; // @[RAM_ST.scala 32:46]
  assign _GEN_3002 = 11'h435 == RADDR ? 11'h435 : _GEN_3001; // @[RAM_ST.scala 32:46]
  assign _GEN_3003 = 11'h436 == RADDR ? 11'h436 : _GEN_3002; // @[RAM_ST.scala 32:46]
  assign _GEN_3004 = 11'h437 == RADDR ? 11'h437 : _GEN_3003; // @[RAM_ST.scala 32:46]
  assign _GEN_3005 = 11'h438 == RADDR ? 11'h438 : _GEN_3004; // @[RAM_ST.scala 32:46]
  assign _GEN_3006 = 11'h439 == RADDR ? 11'h439 : _GEN_3005; // @[RAM_ST.scala 32:46]
  assign _GEN_3007 = 11'h43a == RADDR ? 11'h43a : _GEN_3006; // @[RAM_ST.scala 32:46]
  assign _GEN_3008 = 11'h43b == RADDR ? 11'h43b : _GEN_3007; // @[RAM_ST.scala 32:46]
  assign _GEN_3009 = 11'h43c == RADDR ? 11'h43c : _GEN_3008; // @[RAM_ST.scala 32:46]
  assign _GEN_3010 = 11'h43d == RADDR ? 11'h43d : _GEN_3009; // @[RAM_ST.scala 32:46]
  assign _GEN_3011 = 11'h43e == RADDR ? 11'h43e : _GEN_3010; // @[RAM_ST.scala 32:46]
  assign _GEN_3012 = 11'h43f == RADDR ? 11'h43f : _GEN_3011; // @[RAM_ST.scala 32:46]
  assign _GEN_3013 = 11'h440 == RADDR ? 11'h440 : _GEN_3012; // @[RAM_ST.scala 32:46]
  assign _GEN_3014 = 11'h441 == RADDR ? 11'h441 : _GEN_3013; // @[RAM_ST.scala 32:46]
  assign _GEN_3015 = 11'h442 == RADDR ? 11'h442 : _GEN_3014; // @[RAM_ST.scala 32:46]
  assign _GEN_3016 = 11'h443 == RADDR ? 11'h443 : _GEN_3015; // @[RAM_ST.scala 32:46]
  assign _GEN_3017 = 11'h444 == RADDR ? 11'h444 : _GEN_3016; // @[RAM_ST.scala 32:46]
  assign _GEN_3018 = 11'h445 == RADDR ? 11'h445 : _GEN_3017; // @[RAM_ST.scala 32:46]
  assign _GEN_3019 = 11'h446 == RADDR ? 11'h446 : _GEN_3018; // @[RAM_ST.scala 32:46]
  assign _GEN_3020 = 11'h447 == RADDR ? 11'h447 : _GEN_3019; // @[RAM_ST.scala 32:46]
  assign _GEN_3021 = 11'h448 == RADDR ? 11'h448 : _GEN_3020; // @[RAM_ST.scala 32:46]
  assign _GEN_3022 = 11'h449 == RADDR ? 11'h449 : _GEN_3021; // @[RAM_ST.scala 32:46]
  assign _GEN_3023 = 11'h44a == RADDR ? 11'h44a : _GEN_3022; // @[RAM_ST.scala 32:46]
  assign _GEN_3024 = 11'h44b == RADDR ? 11'h44b : _GEN_3023; // @[RAM_ST.scala 32:46]
  assign _GEN_3025 = 11'h44c == RADDR ? 11'h44c : _GEN_3024; // @[RAM_ST.scala 32:46]
  assign _GEN_3026 = 11'h44d == RADDR ? 11'h44d : _GEN_3025; // @[RAM_ST.scala 32:46]
  assign _GEN_3027 = 11'h44e == RADDR ? 11'h44e : _GEN_3026; // @[RAM_ST.scala 32:46]
  assign _GEN_3028 = 11'h44f == RADDR ? 11'h44f : _GEN_3027; // @[RAM_ST.scala 32:46]
  assign _GEN_3029 = 11'h450 == RADDR ? 11'h450 : _GEN_3028; // @[RAM_ST.scala 32:46]
  assign _GEN_3030 = 11'h451 == RADDR ? 11'h451 : _GEN_3029; // @[RAM_ST.scala 32:46]
  assign _GEN_3031 = 11'h452 == RADDR ? 11'h452 : _GEN_3030; // @[RAM_ST.scala 32:46]
  assign _GEN_3032 = 11'h453 == RADDR ? 11'h453 : _GEN_3031; // @[RAM_ST.scala 32:46]
  assign _GEN_3033 = 11'h454 == RADDR ? 11'h454 : _GEN_3032; // @[RAM_ST.scala 32:46]
  assign _GEN_3034 = 11'h455 == RADDR ? 11'h455 : _GEN_3033; // @[RAM_ST.scala 32:46]
  assign _GEN_3035 = 11'h456 == RADDR ? 11'h456 : _GEN_3034; // @[RAM_ST.scala 32:46]
  assign _GEN_3036 = 11'h457 == RADDR ? 11'h457 : _GEN_3035; // @[RAM_ST.scala 32:46]
  assign _GEN_3037 = 11'h458 == RADDR ? 11'h458 : _GEN_3036; // @[RAM_ST.scala 32:46]
  assign _GEN_3038 = 11'h459 == RADDR ? 11'h459 : _GEN_3037; // @[RAM_ST.scala 32:46]
  assign _GEN_3039 = 11'h45a == RADDR ? 11'h45a : _GEN_3038; // @[RAM_ST.scala 32:46]
  assign _GEN_3040 = 11'h45b == RADDR ? 11'h45b : _GEN_3039; // @[RAM_ST.scala 32:46]
  assign _GEN_3041 = 11'h45c == RADDR ? 11'h45c : _GEN_3040; // @[RAM_ST.scala 32:46]
  assign _GEN_3042 = 11'h45d == RADDR ? 11'h45d : _GEN_3041; // @[RAM_ST.scala 32:46]
  assign _GEN_3043 = 11'h45e == RADDR ? 11'h45e : _GEN_3042; // @[RAM_ST.scala 32:46]
  assign _GEN_3044 = 11'h45f == RADDR ? 11'h45f : _GEN_3043; // @[RAM_ST.scala 32:46]
  assign _GEN_3045 = 11'h460 == RADDR ? 11'h460 : _GEN_3044; // @[RAM_ST.scala 32:46]
  assign _GEN_3046 = 11'h461 == RADDR ? 11'h461 : _GEN_3045; // @[RAM_ST.scala 32:46]
  assign _GEN_3047 = 11'h462 == RADDR ? 11'h462 : _GEN_3046; // @[RAM_ST.scala 32:46]
  assign _GEN_3048 = 11'h463 == RADDR ? 11'h463 : _GEN_3047; // @[RAM_ST.scala 32:46]
  assign _GEN_3049 = 11'h464 == RADDR ? 11'h464 : _GEN_3048; // @[RAM_ST.scala 32:46]
  assign _GEN_3050 = 11'h465 == RADDR ? 11'h465 : _GEN_3049; // @[RAM_ST.scala 32:46]
  assign _GEN_3051 = 11'h466 == RADDR ? 11'h466 : _GEN_3050; // @[RAM_ST.scala 32:46]
  assign _GEN_3052 = 11'h467 == RADDR ? 11'h467 : _GEN_3051; // @[RAM_ST.scala 32:46]
  assign _GEN_3053 = 11'h468 == RADDR ? 11'h468 : _GEN_3052; // @[RAM_ST.scala 32:46]
  assign _GEN_3054 = 11'h469 == RADDR ? 11'h469 : _GEN_3053; // @[RAM_ST.scala 32:46]
  assign _GEN_3055 = 11'h46a == RADDR ? 11'h46a : _GEN_3054; // @[RAM_ST.scala 32:46]
  assign _GEN_3056 = 11'h46b == RADDR ? 11'h46b : _GEN_3055; // @[RAM_ST.scala 32:46]
  assign _GEN_3057 = 11'h46c == RADDR ? 11'h46c : _GEN_3056; // @[RAM_ST.scala 32:46]
  assign _GEN_3058 = 11'h46d == RADDR ? 11'h46d : _GEN_3057; // @[RAM_ST.scala 32:46]
  assign _GEN_3059 = 11'h46e == RADDR ? 11'h46e : _GEN_3058; // @[RAM_ST.scala 32:46]
  assign _GEN_3060 = 11'h46f == RADDR ? 11'h46f : _GEN_3059; // @[RAM_ST.scala 32:46]
  assign _GEN_3061 = 11'h470 == RADDR ? 11'h470 : _GEN_3060; // @[RAM_ST.scala 32:46]
  assign _GEN_3062 = 11'h471 == RADDR ? 11'h471 : _GEN_3061; // @[RAM_ST.scala 32:46]
  assign _GEN_3063 = 11'h472 == RADDR ? 11'h472 : _GEN_3062; // @[RAM_ST.scala 32:46]
  assign _GEN_3064 = 11'h473 == RADDR ? 11'h473 : _GEN_3063; // @[RAM_ST.scala 32:46]
  assign _GEN_3065 = 11'h474 == RADDR ? 11'h474 : _GEN_3064; // @[RAM_ST.scala 32:46]
  assign _GEN_3066 = 11'h475 == RADDR ? 11'h475 : _GEN_3065; // @[RAM_ST.scala 32:46]
  assign _GEN_3067 = 11'h476 == RADDR ? 11'h476 : _GEN_3066; // @[RAM_ST.scala 32:46]
  assign _GEN_3068 = 11'h477 == RADDR ? 11'h477 : _GEN_3067; // @[RAM_ST.scala 32:46]
  assign _GEN_3069 = 11'h478 == RADDR ? 11'h478 : _GEN_3068; // @[RAM_ST.scala 32:46]
  assign _GEN_3070 = 11'h479 == RADDR ? 11'h479 : _GEN_3069; // @[RAM_ST.scala 32:46]
  assign _GEN_3071 = 11'h47a == RADDR ? 11'h47a : _GEN_3070; // @[RAM_ST.scala 32:46]
  assign _GEN_3072 = 11'h47b == RADDR ? 11'h47b : _GEN_3071; // @[RAM_ST.scala 32:46]
  assign _GEN_3073 = 11'h47c == RADDR ? 11'h47c : _GEN_3072; // @[RAM_ST.scala 32:46]
  assign _GEN_3074 = 11'h47d == RADDR ? 11'h47d : _GEN_3073; // @[RAM_ST.scala 32:46]
  assign _GEN_3075 = 11'h47e == RADDR ? 11'h47e : _GEN_3074; // @[RAM_ST.scala 32:46]
  assign _GEN_3076 = 11'h47f == RADDR ? 11'h47f : _GEN_3075; // @[RAM_ST.scala 32:46]
  assign _GEN_3077 = 11'h480 == RADDR ? 11'h480 : _GEN_3076; // @[RAM_ST.scala 32:46]
  assign _GEN_3078 = 11'h481 == RADDR ? 11'h481 : _GEN_3077; // @[RAM_ST.scala 32:46]
  assign _GEN_3079 = 11'h482 == RADDR ? 11'h482 : _GEN_3078; // @[RAM_ST.scala 32:46]
  assign _GEN_3080 = 11'h483 == RADDR ? 11'h483 : _GEN_3079; // @[RAM_ST.scala 32:46]
  assign _GEN_3081 = 11'h484 == RADDR ? 11'h484 : _GEN_3080; // @[RAM_ST.scala 32:46]
  assign _GEN_3082 = 11'h485 == RADDR ? 11'h485 : _GEN_3081; // @[RAM_ST.scala 32:46]
  assign _GEN_3083 = 11'h486 == RADDR ? 11'h486 : _GEN_3082; // @[RAM_ST.scala 32:46]
  assign _GEN_3084 = 11'h487 == RADDR ? 11'h487 : _GEN_3083; // @[RAM_ST.scala 32:46]
  assign _GEN_3085 = 11'h488 == RADDR ? 11'h488 : _GEN_3084; // @[RAM_ST.scala 32:46]
  assign _GEN_3086 = 11'h489 == RADDR ? 11'h489 : _GEN_3085; // @[RAM_ST.scala 32:46]
  assign _GEN_3087 = 11'h48a == RADDR ? 11'h48a : _GEN_3086; // @[RAM_ST.scala 32:46]
  assign _GEN_3088 = 11'h48b == RADDR ? 11'h48b : _GEN_3087; // @[RAM_ST.scala 32:46]
  assign _GEN_3089 = 11'h48c == RADDR ? 11'h48c : _GEN_3088; // @[RAM_ST.scala 32:46]
  assign _GEN_3090 = 11'h48d == RADDR ? 11'h48d : _GEN_3089; // @[RAM_ST.scala 32:46]
  assign _GEN_3091 = 11'h48e == RADDR ? 11'h48e : _GEN_3090; // @[RAM_ST.scala 32:46]
  assign _GEN_3092 = 11'h48f == RADDR ? 11'h48f : _GEN_3091; // @[RAM_ST.scala 32:46]
  assign _GEN_3093 = 11'h490 == RADDR ? 11'h490 : _GEN_3092; // @[RAM_ST.scala 32:46]
  assign _GEN_3094 = 11'h491 == RADDR ? 11'h491 : _GEN_3093; // @[RAM_ST.scala 32:46]
  assign _GEN_3095 = 11'h492 == RADDR ? 11'h492 : _GEN_3094; // @[RAM_ST.scala 32:46]
  assign _GEN_3096 = 11'h493 == RADDR ? 11'h493 : _GEN_3095; // @[RAM_ST.scala 32:46]
  assign _GEN_3097 = 11'h494 == RADDR ? 11'h494 : _GEN_3096; // @[RAM_ST.scala 32:46]
  assign _GEN_3098 = 11'h495 == RADDR ? 11'h495 : _GEN_3097; // @[RAM_ST.scala 32:46]
  assign _GEN_3099 = 11'h496 == RADDR ? 11'h496 : _GEN_3098; // @[RAM_ST.scala 32:46]
  assign _GEN_3100 = 11'h497 == RADDR ? 11'h497 : _GEN_3099; // @[RAM_ST.scala 32:46]
  assign _GEN_3101 = 11'h498 == RADDR ? 11'h498 : _GEN_3100; // @[RAM_ST.scala 32:46]
  assign _GEN_3102 = 11'h499 == RADDR ? 11'h499 : _GEN_3101; // @[RAM_ST.scala 32:46]
  assign _GEN_3103 = 11'h49a == RADDR ? 11'h49a : _GEN_3102; // @[RAM_ST.scala 32:46]
  assign _GEN_3104 = 11'h49b == RADDR ? 11'h49b : _GEN_3103; // @[RAM_ST.scala 32:46]
  assign _GEN_3105 = 11'h49c == RADDR ? 11'h49c : _GEN_3104; // @[RAM_ST.scala 32:46]
  assign _GEN_3106 = 11'h49d == RADDR ? 11'h49d : _GEN_3105; // @[RAM_ST.scala 32:46]
  assign _GEN_3107 = 11'h49e == RADDR ? 11'h49e : _GEN_3106; // @[RAM_ST.scala 32:46]
  assign _GEN_3108 = 11'h49f == RADDR ? 11'h49f : _GEN_3107; // @[RAM_ST.scala 32:46]
  assign _GEN_3109 = 11'h4a0 == RADDR ? 11'h4a0 : _GEN_3108; // @[RAM_ST.scala 32:46]
  assign _GEN_3110 = 11'h4a1 == RADDR ? 11'h4a1 : _GEN_3109; // @[RAM_ST.scala 32:46]
  assign _GEN_3111 = 11'h4a2 == RADDR ? 11'h4a2 : _GEN_3110; // @[RAM_ST.scala 32:46]
  assign _GEN_3112 = 11'h4a3 == RADDR ? 11'h4a3 : _GEN_3111; // @[RAM_ST.scala 32:46]
  assign _GEN_3113 = 11'h4a4 == RADDR ? 11'h4a4 : _GEN_3112; // @[RAM_ST.scala 32:46]
  assign _GEN_3114 = 11'h4a5 == RADDR ? 11'h4a5 : _GEN_3113; // @[RAM_ST.scala 32:46]
  assign _GEN_3115 = 11'h4a6 == RADDR ? 11'h4a6 : _GEN_3114; // @[RAM_ST.scala 32:46]
  assign _GEN_3116 = 11'h4a7 == RADDR ? 11'h4a7 : _GEN_3115; // @[RAM_ST.scala 32:46]
  assign _GEN_3117 = 11'h4a8 == RADDR ? 11'h4a8 : _GEN_3116; // @[RAM_ST.scala 32:46]
  assign _GEN_3118 = 11'h4a9 == RADDR ? 11'h4a9 : _GEN_3117; // @[RAM_ST.scala 32:46]
  assign _GEN_3119 = 11'h4aa == RADDR ? 11'h4aa : _GEN_3118; // @[RAM_ST.scala 32:46]
  assign _GEN_3120 = 11'h4ab == RADDR ? 11'h4ab : _GEN_3119; // @[RAM_ST.scala 32:46]
  assign _GEN_3121 = 11'h4ac == RADDR ? 11'h4ac : _GEN_3120; // @[RAM_ST.scala 32:46]
  assign _GEN_3122 = 11'h4ad == RADDR ? 11'h4ad : _GEN_3121; // @[RAM_ST.scala 32:46]
  assign _GEN_3123 = 11'h4ae == RADDR ? 11'h4ae : _GEN_3122; // @[RAM_ST.scala 32:46]
  assign _GEN_3124 = 11'h4af == RADDR ? 11'h4af : _GEN_3123; // @[RAM_ST.scala 32:46]
  assign _GEN_3125 = 11'h4b0 == RADDR ? 11'h4b0 : _GEN_3124; // @[RAM_ST.scala 32:46]
  assign _GEN_3126 = 11'h4b1 == RADDR ? 11'h4b1 : _GEN_3125; // @[RAM_ST.scala 32:46]
  assign _GEN_3127 = 11'h4b2 == RADDR ? 11'h4b2 : _GEN_3126; // @[RAM_ST.scala 32:46]
  assign _GEN_3128 = 11'h4b3 == RADDR ? 11'h4b3 : _GEN_3127; // @[RAM_ST.scala 32:46]
  assign _GEN_3129 = 11'h4b4 == RADDR ? 11'h4b4 : _GEN_3128; // @[RAM_ST.scala 32:46]
  assign _GEN_3130 = 11'h4b5 == RADDR ? 11'h4b5 : _GEN_3129; // @[RAM_ST.scala 32:46]
  assign _GEN_3131 = 11'h4b6 == RADDR ? 11'h4b6 : _GEN_3130; // @[RAM_ST.scala 32:46]
  assign _GEN_3132 = 11'h4b7 == RADDR ? 11'h4b7 : _GEN_3131; // @[RAM_ST.scala 32:46]
  assign _GEN_3133 = 11'h4b8 == RADDR ? 11'h4b8 : _GEN_3132; // @[RAM_ST.scala 32:46]
  assign _GEN_3134 = 11'h4b9 == RADDR ? 11'h4b9 : _GEN_3133; // @[RAM_ST.scala 32:46]
  assign _GEN_3135 = 11'h4ba == RADDR ? 11'h4ba : _GEN_3134; // @[RAM_ST.scala 32:46]
  assign _GEN_3136 = 11'h4bb == RADDR ? 11'h4bb : _GEN_3135; // @[RAM_ST.scala 32:46]
  assign _GEN_3137 = 11'h4bc == RADDR ? 11'h4bc : _GEN_3136; // @[RAM_ST.scala 32:46]
  assign _GEN_3138 = 11'h4bd == RADDR ? 11'h4bd : _GEN_3137; // @[RAM_ST.scala 32:46]
  assign _GEN_3139 = 11'h4be == RADDR ? 11'h4be : _GEN_3138; // @[RAM_ST.scala 32:46]
  assign _GEN_3140 = 11'h4bf == RADDR ? 11'h4bf : _GEN_3139; // @[RAM_ST.scala 32:46]
  assign _GEN_3141 = 11'h4c0 == RADDR ? 11'h4c0 : _GEN_3140; // @[RAM_ST.scala 32:46]
  assign _GEN_3142 = 11'h4c1 == RADDR ? 11'h4c1 : _GEN_3141; // @[RAM_ST.scala 32:46]
  assign _GEN_3143 = 11'h4c2 == RADDR ? 11'h4c2 : _GEN_3142; // @[RAM_ST.scala 32:46]
  assign _GEN_3144 = 11'h4c3 == RADDR ? 11'h4c3 : _GEN_3143; // @[RAM_ST.scala 32:46]
  assign _GEN_3145 = 11'h4c4 == RADDR ? 11'h4c4 : _GEN_3144; // @[RAM_ST.scala 32:46]
  assign _GEN_3146 = 11'h4c5 == RADDR ? 11'h4c5 : _GEN_3145; // @[RAM_ST.scala 32:46]
  assign _GEN_3147 = 11'h4c6 == RADDR ? 11'h4c6 : _GEN_3146; // @[RAM_ST.scala 32:46]
  assign _GEN_3148 = 11'h4c7 == RADDR ? 11'h4c7 : _GEN_3147; // @[RAM_ST.scala 32:46]
  assign _GEN_3149 = 11'h4c8 == RADDR ? 11'h4c8 : _GEN_3148; // @[RAM_ST.scala 32:46]
  assign _GEN_3150 = 11'h4c9 == RADDR ? 11'h4c9 : _GEN_3149; // @[RAM_ST.scala 32:46]
  assign _GEN_3151 = 11'h4ca == RADDR ? 11'h4ca : _GEN_3150; // @[RAM_ST.scala 32:46]
  assign _GEN_3152 = 11'h4cb == RADDR ? 11'h4cb : _GEN_3151; // @[RAM_ST.scala 32:46]
  assign _GEN_3153 = 11'h4cc == RADDR ? 11'h4cc : _GEN_3152; // @[RAM_ST.scala 32:46]
  assign _GEN_3154 = 11'h4cd == RADDR ? 11'h4cd : _GEN_3153; // @[RAM_ST.scala 32:46]
  assign _GEN_3155 = 11'h4ce == RADDR ? 11'h4ce : _GEN_3154; // @[RAM_ST.scala 32:46]
  assign _GEN_3156 = 11'h4cf == RADDR ? 11'h4cf : _GEN_3155; // @[RAM_ST.scala 32:46]
  assign _GEN_3157 = 11'h4d0 == RADDR ? 11'h4d0 : _GEN_3156; // @[RAM_ST.scala 32:46]
  assign _GEN_3158 = 11'h4d1 == RADDR ? 11'h4d1 : _GEN_3157; // @[RAM_ST.scala 32:46]
  assign _GEN_3159 = 11'h4d2 == RADDR ? 11'h4d2 : _GEN_3158; // @[RAM_ST.scala 32:46]
  assign _GEN_3160 = 11'h4d3 == RADDR ? 11'h4d3 : _GEN_3159; // @[RAM_ST.scala 32:46]
  assign _GEN_3161 = 11'h4d4 == RADDR ? 11'h4d4 : _GEN_3160; // @[RAM_ST.scala 32:46]
  assign _GEN_3162 = 11'h4d5 == RADDR ? 11'h4d5 : _GEN_3161; // @[RAM_ST.scala 32:46]
  assign _GEN_3163 = 11'h4d6 == RADDR ? 11'h4d6 : _GEN_3162; // @[RAM_ST.scala 32:46]
  assign _GEN_3164 = 11'h4d7 == RADDR ? 11'h4d7 : _GEN_3163; // @[RAM_ST.scala 32:46]
  assign _GEN_3165 = 11'h4d8 == RADDR ? 11'h4d8 : _GEN_3164; // @[RAM_ST.scala 32:46]
  assign _GEN_3166 = 11'h4d9 == RADDR ? 11'h4d9 : _GEN_3165; // @[RAM_ST.scala 32:46]
  assign _GEN_3167 = 11'h4da == RADDR ? 11'h4da : _GEN_3166; // @[RAM_ST.scala 32:46]
  assign _GEN_3168 = 11'h4db == RADDR ? 11'h4db : _GEN_3167; // @[RAM_ST.scala 32:46]
  assign _GEN_3169 = 11'h4dc == RADDR ? 11'h4dc : _GEN_3168; // @[RAM_ST.scala 32:46]
  assign _GEN_3170 = 11'h4dd == RADDR ? 11'h4dd : _GEN_3169; // @[RAM_ST.scala 32:46]
  assign _GEN_3171 = 11'h4de == RADDR ? 11'h4de : _GEN_3170; // @[RAM_ST.scala 32:46]
  assign _GEN_3172 = 11'h4df == RADDR ? 11'h4df : _GEN_3171; // @[RAM_ST.scala 32:46]
  assign _GEN_3173 = 11'h4e0 == RADDR ? 11'h4e0 : _GEN_3172; // @[RAM_ST.scala 32:46]
  assign _GEN_3174 = 11'h4e1 == RADDR ? 11'h4e1 : _GEN_3173; // @[RAM_ST.scala 32:46]
  assign _GEN_3175 = 11'h4e2 == RADDR ? 11'h4e2 : _GEN_3174; // @[RAM_ST.scala 32:46]
  assign _GEN_3176 = 11'h4e3 == RADDR ? 11'h4e3 : _GEN_3175; // @[RAM_ST.scala 32:46]
  assign _GEN_3177 = 11'h4e4 == RADDR ? 11'h4e4 : _GEN_3176; // @[RAM_ST.scala 32:46]
  assign _GEN_3178 = 11'h4e5 == RADDR ? 11'h4e5 : _GEN_3177; // @[RAM_ST.scala 32:46]
  assign _GEN_3179 = 11'h4e6 == RADDR ? 11'h4e6 : _GEN_3178; // @[RAM_ST.scala 32:46]
  assign _GEN_3180 = 11'h4e7 == RADDR ? 11'h4e7 : _GEN_3179; // @[RAM_ST.scala 32:46]
  assign _GEN_3181 = 11'h4e8 == RADDR ? 11'h4e8 : _GEN_3180; // @[RAM_ST.scala 32:46]
  assign _GEN_3182 = 11'h4e9 == RADDR ? 11'h4e9 : _GEN_3181; // @[RAM_ST.scala 32:46]
  assign _GEN_3183 = 11'h4ea == RADDR ? 11'h4ea : _GEN_3182; // @[RAM_ST.scala 32:46]
  assign _GEN_3184 = 11'h4eb == RADDR ? 11'h4eb : _GEN_3183; // @[RAM_ST.scala 32:46]
  assign _GEN_3185 = 11'h4ec == RADDR ? 11'h4ec : _GEN_3184; // @[RAM_ST.scala 32:46]
  assign _GEN_3186 = 11'h4ed == RADDR ? 11'h4ed : _GEN_3185; // @[RAM_ST.scala 32:46]
  assign _GEN_3187 = 11'h4ee == RADDR ? 11'h4ee : _GEN_3186; // @[RAM_ST.scala 32:46]
  assign _GEN_3188 = 11'h4ef == RADDR ? 11'h4ef : _GEN_3187; // @[RAM_ST.scala 32:46]
  assign _GEN_3189 = 11'h4f0 == RADDR ? 11'h4f0 : _GEN_3188; // @[RAM_ST.scala 32:46]
  assign _GEN_3190 = 11'h4f1 == RADDR ? 11'h4f1 : _GEN_3189; // @[RAM_ST.scala 32:46]
  assign _GEN_3191 = 11'h4f2 == RADDR ? 11'h4f2 : _GEN_3190; // @[RAM_ST.scala 32:46]
  assign _GEN_3192 = 11'h4f3 == RADDR ? 11'h4f3 : _GEN_3191; // @[RAM_ST.scala 32:46]
  assign _GEN_3193 = 11'h4f4 == RADDR ? 11'h4f4 : _GEN_3192; // @[RAM_ST.scala 32:46]
  assign _GEN_3194 = 11'h4f5 == RADDR ? 11'h4f5 : _GEN_3193; // @[RAM_ST.scala 32:46]
  assign _GEN_3195 = 11'h4f6 == RADDR ? 11'h4f6 : _GEN_3194; // @[RAM_ST.scala 32:46]
  assign _GEN_3196 = 11'h4f7 == RADDR ? 11'h4f7 : _GEN_3195; // @[RAM_ST.scala 32:46]
  assign _GEN_3197 = 11'h4f8 == RADDR ? 11'h4f8 : _GEN_3196; // @[RAM_ST.scala 32:46]
  assign _GEN_3198 = 11'h4f9 == RADDR ? 11'h4f9 : _GEN_3197; // @[RAM_ST.scala 32:46]
  assign _GEN_3199 = 11'h4fa == RADDR ? 11'h4fa : _GEN_3198; // @[RAM_ST.scala 32:46]
  assign _GEN_3200 = 11'h4fb == RADDR ? 11'h4fb : _GEN_3199; // @[RAM_ST.scala 32:46]
  assign _GEN_3201 = 11'h4fc == RADDR ? 11'h4fc : _GEN_3200; // @[RAM_ST.scala 32:46]
  assign _GEN_3202 = 11'h4fd == RADDR ? 11'h4fd : _GEN_3201; // @[RAM_ST.scala 32:46]
  assign _GEN_3203 = 11'h4fe == RADDR ? 11'h4fe : _GEN_3202; // @[RAM_ST.scala 32:46]
  assign _GEN_3204 = 11'h4ff == RADDR ? 11'h4ff : _GEN_3203; // @[RAM_ST.scala 32:46]
  assign _GEN_3205 = 11'h500 == RADDR ? 11'h500 : _GEN_3204; // @[RAM_ST.scala 32:46]
  assign _GEN_3206 = 11'h501 == RADDR ? 11'h501 : _GEN_3205; // @[RAM_ST.scala 32:46]
  assign _GEN_3207 = 11'h502 == RADDR ? 11'h502 : _GEN_3206; // @[RAM_ST.scala 32:46]
  assign _GEN_3208 = 11'h503 == RADDR ? 11'h503 : _GEN_3207; // @[RAM_ST.scala 32:46]
  assign _GEN_3209 = 11'h504 == RADDR ? 11'h504 : _GEN_3208; // @[RAM_ST.scala 32:46]
  assign _GEN_3210 = 11'h505 == RADDR ? 11'h505 : _GEN_3209; // @[RAM_ST.scala 32:46]
  assign _GEN_3211 = 11'h506 == RADDR ? 11'h506 : _GEN_3210; // @[RAM_ST.scala 32:46]
  assign _GEN_3212 = 11'h507 == RADDR ? 11'h507 : _GEN_3211; // @[RAM_ST.scala 32:46]
  assign _GEN_3213 = 11'h508 == RADDR ? 11'h508 : _GEN_3212; // @[RAM_ST.scala 32:46]
  assign _GEN_3214 = 11'h509 == RADDR ? 11'h509 : _GEN_3213; // @[RAM_ST.scala 32:46]
  assign _GEN_3215 = 11'h50a == RADDR ? 11'h50a : _GEN_3214; // @[RAM_ST.scala 32:46]
  assign _GEN_3216 = 11'h50b == RADDR ? 11'h50b : _GEN_3215; // @[RAM_ST.scala 32:46]
  assign _GEN_3217 = 11'h50c == RADDR ? 11'h50c : _GEN_3216; // @[RAM_ST.scala 32:46]
  assign _GEN_3218 = 11'h50d == RADDR ? 11'h50d : _GEN_3217; // @[RAM_ST.scala 32:46]
  assign _GEN_3219 = 11'h50e == RADDR ? 11'h50e : _GEN_3218; // @[RAM_ST.scala 32:46]
  assign _GEN_3220 = 11'h50f == RADDR ? 11'h50f : _GEN_3219; // @[RAM_ST.scala 32:46]
  assign _GEN_3221 = 11'h510 == RADDR ? 11'h510 : _GEN_3220; // @[RAM_ST.scala 32:46]
  assign _GEN_3222 = 11'h511 == RADDR ? 11'h511 : _GEN_3221; // @[RAM_ST.scala 32:46]
  assign _GEN_3223 = 11'h512 == RADDR ? 11'h512 : _GEN_3222; // @[RAM_ST.scala 32:46]
  assign _GEN_3224 = 11'h513 == RADDR ? 11'h513 : _GEN_3223; // @[RAM_ST.scala 32:46]
  assign _GEN_3225 = 11'h514 == RADDR ? 11'h514 : _GEN_3224; // @[RAM_ST.scala 32:46]
  assign _GEN_3226 = 11'h515 == RADDR ? 11'h515 : _GEN_3225; // @[RAM_ST.scala 32:46]
  assign _GEN_3227 = 11'h516 == RADDR ? 11'h516 : _GEN_3226; // @[RAM_ST.scala 32:46]
  assign _GEN_3228 = 11'h517 == RADDR ? 11'h517 : _GEN_3227; // @[RAM_ST.scala 32:46]
  assign _GEN_3229 = 11'h518 == RADDR ? 11'h518 : _GEN_3228; // @[RAM_ST.scala 32:46]
  assign _GEN_3230 = 11'h519 == RADDR ? 11'h519 : _GEN_3229; // @[RAM_ST.scala 32:46]
  assign _GEN_3231 = 11'h51a == RADDR ? 11'h51a : _GEN_3230; // @[RAM_ST.scala 32:46]
  assign _GEN_3232 = 11'h51b == RADDR ? 11'h51b : _GEN_3231; // @[RAM_ST.scala 32:46]
  assign _GEN_3233 = 11'h51c == RADDR ? 11'h51c : _GEN_3232; // @[RAM_ST.scala 32:46]
  assign _GEN_3234 = 11'h51d == RADDR ? 11'h51d : _GEN_3233; // @[RAM_ST.scala 32:46]
  assign _GEN_3235 = 11'h51e == RADDR ? 11'h51e : _GEN_3234; // @[RAM_ST.scala 32:46]
  assign _GEN_3236 = 11'h51f == RADDR ? 11'h51f : _GEN_3235; // @[RAM_ST.scala 32:46]
  assign _GEN_3237 = 11'h520 == RADDR ? 11'h520 : _GEN_3236; // @[RAM_ST.scala 32:46]
  assign _GEN_3238 = 11'h521 == RADDR ? 11'h521 : _GEN_3237; // @[RAM_ST.scala 32:46]
  assign _GEN_3239 = 11'h522 == RADDR ? 11'h522 : _GEN_3238; // @[RAM_ST.scala 32:46]
  assign _GEN_3240 = 11'h523 == RADDR ? 11'h523 : _GEN_3239; // @[RAM_ST.scala 32:46]
  assign _GEN_3241 = 11'h524 == RADDR ? 11'h524 : _GEN_3240; // @[RAM_ST.scala 32:46]
  assign _GEN_3242 = 11'h525 == RADDR ? 11'h525 : _GEN_3241; // @[RAM_ST.scala 32:46]
  assign _GEN_3243 = 11'h526 == RADDR ? 11'h526 : _GEN_3242; // @[RAM_ST.scala 32:46]
  assign _GEN_3244 = 11'h527 == RADDR ? 11'h527 : _GEN_3243; // @[RAM_ST.scala 32:46]
  assign _GEN_3245 = 11'h528 == RADDR ? 11'h528 : _GEN_3244; // @[RAM_ST.scala 32:46]
  assign _GEN_3246 = 11'h529 == RADDR ? 11'h529 : _GEN_3245; // @[RAM_ST.scala 32:46]
  assign _GEN_3247 = 11'h52a == RADDR ? 11'h52a : _GEN_3246; // @[RAM_ST.scala 32:46]
  assign _GEN_3248 = 11'h52b == RADDR ? 11'h52b : _GEN_3247; // @[RAM_ST.scala 32:46]
  assign _GEN_3249 = 11'h52c == RADDR ? 11'h52c : _GEN_3248; // @[RAM_ST.scala 32:46]
  assign _GEN_3250 = 11'h52d == RADDR ? 11'h52d : _GEN_3249; // @[RAM_ST.scala 32:46]
  assign _GEN_3251 = 11'h52e == RADDR ? 11'h52e : _GEN_3250; // @[RAM_ST.scala 32:46]
  assign _GEN_3252 = 11'h52f == RADDR ? 11'h52f : _GEN_3251; // @[RAM_ST.scala 32:46]
  assign _GEN_3253 = 11'h530 == RADDR ? 11'h530 : _GEN_3252; // @[RAM_ST.scala 32:46]
  assign _GEN_3254 = 11'h531 == RADDR ? 11'h531 : _GEN_3253; // @[RAM_ST.scala 32:46]
  assign _GEN_3255 = 11'h532 == RADDR ? 11'h532 : _GEN_3254; // @[RAM_ST.scala 32:46]
  assign _GEN_3256 = 11'h533 == RADDR ? 11'h533 : _GEN_3255; // @[RAM_ST.scala 32:46]
  assign _GEN_3257 = 11'h534 == RADDR ? 11'h534 : _GEN_3256; // @[RAM_ST.scala 32:46]
  assign _GEN_3258 = 11'h535 == RADDR ? 11'h535 : _GEN_3257; // @[RAM_ST.scala 32:46]
  assign _GEN_3259 = 11'h536 == RADDR ? 11'h536 : _GEN_3258; // @[RAM_ST.scala 32:46]
  assign _GEN_3260 = 11'h537 == RADDR ? 11'h537 : _GEN_3259; // @[RAM_ST.scala 32:46]
  assign _GEN_3261 = 11'h538 == RADDR ? 11'h538 : _GEN_3260; // @[RAM_ST.scala 32:46]
  assign _GEN_3262 = 11'h539 == RADDR ? 11'h539 : _GEN_3261; // @[RAM_ST.scala 32:46]
  assign _GEN_3263 = 11'h53a == RADDR ? 11'h53a : _GEN_3262; // @[RAM_ST.scala 32:46]
  assign _GEN_3264 = 11'h53b == RADDR ? 11'h53b : _GEN_3263; // @[RAM_ST.scala 32:46]
  assign _GEN_3265 = 11'h53c == RADDR ? 11'h53c : _GEN_3264; // @[RAM_ST.scala 32:46]
  assign _GEN_3266 = 11'h53d == RADDR ? 11'h53d : _GEN_3265; // @[RAM_ST.scala 32:46]
  assign _GEN_3267 = 11'h53e == RADDR ? 11'h53e : _GEN_3266; // @[RAM_ST.scala 32:46]
  assign _GEN_3268 = 11'h53f == RADDR ? 11'h53f : _GEN_3267; // @[RAM_ST.scala 32:46]
  assign _GEN_3269 = 11'h540 == RADDR ? 11'h540 : _GEN_3268; // @[RAM_ST.scala 32:46]
  assign _GEN_3270 = 11'h541 == RADDR ? 11'h541 : _GEN_3269; // @[RAM_ST.scala 32:46]
  assign _GEN_3271 = 11'h542 == RADDR ? 11'h542 : _GEN_3270; // @[RAM_ST.scala 32:46]
  assign _GEN_3272 = 11'h543 == RADDR ? 11'h543 : _GEN_3271; // @[RAM_ST.scala 32:46]
  assign _GEN_3273 = 11'h544 == RADDR ? 11'h544 : _GEN_3272; // @[RAM_ST.scala 32:46]
  assign _GEN_3274 = 11'h545 == RADDR ? 11'h545 : _GEN_3273; // @[RAM_ST.scala 32:46]
  assign _GEN_3275 = 11'h546 == RADDR ? 11'h546 : _GEN_3274; // @[RAM_ST.scala 32:46]
  assign _GEN_3276 = 11'h547 == RADDR ? 11'h547 : _GEN_3275; // @[RAM_ST.scala 32:46]
  assign _GEN_3277 = 11'h548 == RADDR ? 11'h548 : _GEN_3276; // @[RAM_ST.scala 32:46]
  assign _GEN_3278 = 11'h549 == RADDR ? 11'h549 : _GEN_3277; // @[RAM_ST.scala 32:46]
  assign _GEN_3279 = 11'h54a == RADDR ? 11'h54a : _GEN_3278; // @[RAM_ST.scala 32:46]
  assign _GEN_3280 = 11'h54b == RADDR ? 11'h54b : _GEN_3279; // @[RAM_ST.scala 32:46]
  assign _GEN_3281 = 11'h54c == RADDR ? 11'h54c : _GEN_3280; // @[RAM_ST.scala 32:46]
  assign _GEN_3282 = 11'h54d == RADDR ? 11'h54d : _GEN_3281; // @[RAM_ST.scala 32:46]
  assign _GEN_3283 = 11'h54e == RADDR ? 11'h54e : _GEN_3282; // @[RAM_ST.scala 32:46]
  assign _GEN_3284 = 11'h54f == RADDR ? 11'h54f : _GEN_3283; // @[RAM_ST.scala 32:46]
  assign _GEN_3285 = 11'h550 == RADDR ? 11'h550 : _GEN_3284; // @[RAM_ST.scala 32:46]
  assign _GEN_3286 = 11'h551 == RADDR ? 11'h551 : _GEN_3285; // @[RAM_ST.scala 32:46]
  assign _GEN_3287 = 11'h552 == RADDR ? 11'h552 : _GEN_3286; // @[RAM_ST.scala 32:46]
  assign _GEN_3288 = 11'h553 == RADDR ? 11'h553 : _GEN_3287; // @[RAM_ST.scala 32:46]
  assign _GEN_3289 = 11'h554 == RADDR ? 11'h554 : _GEN_3288; // @[RAM_ST.scala 32:46]
  assign _GEN_3290 = 11'h555 == RADDR ? 11'h555 : _GEN_3289; // @[RAM_ST.scala 32:46]
  assign _GEN_3291 = 11'h556 == RADDR ? 11'h556 : _GEN_3290; // @[RAM_ST.scala 32:46]
  assign _GEN_3292 = 11'h557 == RADDR ? 11'h557 : _GEN_3291; // @[RAM_ST.scala 32:46]
  assign _GEN_3293 = 11'h558 == RADDR ? 11'h558 : _GEN_3292; // @[RAM_ST.scala 32:46]
  assign _GEN_3294 = 11'h559 == RADDR ? 11'h559 : _GEN_3293; // @[RAM_ST.scala 32:46]
  assign _GEN_3295 = 11'h55a == RADDR ? 11'h55a : _GEN_3294; // @[RAM_ST.scala 32:46]
  assign _GEN_3296 = 11'h55b == RADDR ? 11'h55b : _GEN_3295; // @[RAM_ST.scala 32:46]
  assign _GEN_3297 = 11'h55c == RADDR ? 11'h55c : _GEN_3296; // @[RAM_ST.scala 32:46]
  assign _GEN_3298 = 11'h55d == RADDR ? 11'h55d : _GEN_3297; // @[RAM_ST.scala 32:46]
  assign _GEN_3299 = 11'h55e == RADDR ? 11'h55e : _GEN_3298; // @[RAM_ST.scala 32:46]
  assign _GEN_3300 = 11'h55f == RADDR ? 11'h55f : _GEN_3299; // @[RAM_ST.scala 32:46]
  assign _GEN_3301 = 11'h560 == RADDR ? 11'h560 : _GEN_3300; // @[RAM_ST.scala 32:46]
  assign _GEN_3302 = 11'h561 == RADDR ? 11'h561 : _GEN_3301; // @[RAM_ST.scala 32:46]
  assign _GEN_3303 = 11'h562 == RADDR ? 11'h562 : _GEN_3302; // @[RAM_ST.scala 32:46]
  assign _GEN_3304 = 11'h563 == RADDR ? 11'h563 : _GEN_3303; // @[RAM_ST.scala 32:46]
  assign _GEN_3305 = 11'h564 == RADDR ? 11'h564 : _GEN_3304; // @[RAM_ST.scala 32:46]
  assign _GEN_3306 = 11'h565 == RADDR ? 11'h565 : _GEN_3305; // @[RAM_ST.scala 32:46]
  assign _GEN_3307 = 11'h566 == RADDR ? 11'h566 : _GEN_3306; // @[RAM_ST.scala 32:46]
  assign _GEN_3308 = 11'h567 == RADDR ? 11'h567 : _GEN_3307; // @[RAM_ST.scala 32:46]
  assign _GEN_3309 = 11'h568 == RADDR ? 11'h568 : _GEN_3308; // @[RAM_ST.scala 32:46]
  assign _GEN_3310 = 11'h569 == RADDR ? 11'h569 : _GEN_3309; // @[RAM_ST.scala 32:46]
  assign _GEN_3311 = 11'h56a == RADDR ? 11'h56a : _GEN_3310; // @[RAM_ST.scala 32:46]
  assign _GEN_3312 = 11'h56b == RADDR ? 11'h56b : _GEN_3311; // @[RAM_ST.scala 32:46]
  assign _GEN_3313 = 11'h56c == RADDR ? 11'h56c : _GEN_3312; // @[RAM_ST.scala 32:46]
  assign _GEN_3314 = 11'h56d == RADDR ? 11'h56d : _GEN_3313; // @[RAM_ST.scala 32:46]
  assign _GEN_3315 = 11'h56e == RADDR ? 11'h56e : _GEN_3314; // @[RAM_ST.scala 32:46]
  assign _GEN_3316 = 11'h56f == RADDR ? 11'h56f : _GEN_3315; // @[RAM_ST.scala 32:46]
  assign _GEN_3317 = 11'h570 == RADDR ? 11'h570 : _GEN_3316; // @[RAM_ST.scala 32:46]
  assign _GEN_3318 = 11'h571 == RADDR ? 11'h571 : _GEN_3317; // @[RAM_ST.scala 32:46]
  assign _GEN_3319 = 11'h572 == RADDR ? 11'h572 : _GEN_3318; // @[RAM_ST.scala 32:46]
  assign _GEN_3320 = 11'h573 == RADDR ? 11'h573 : _GEN_3319; // @[RAM_ST.scala 32:46]
  assign _GEN_3321 = 11'h574 == RADDR ? 11'h574 : _GEN_3320; // @[RAM_ST.scala 32:46]
  assign _GEN_3322 = 11'h575 == RADDR ? 11'h575 : _GEN_3321; // @[RAM_ST.scala 32:46]
  assign _GEN_3323 = 11'h576 == RADDR ? 11'h576 : _GEN_3322; // @[RAM_ST.scala 32:46]
  assign _GEN_3324 = 11'h577 == RADDR ? 11'h577 : _GEN_3323; // @[RAM_ST.scala 32:46]
  assign _GEN_3325 = 11'h578 == RADDR ? 11'h578 : _GEN_3324; // @[RAM_ST.scala 32:46]
  assign _GEN_3326 = 11'h579 == RADDR ? 11'h579 : _GEN_3325; // @[RAM_ST.scala 32:46]
  assign _GEN_3327 = 11'h57a == RADDR ? 11'h57a : _GEN_3326; // @[RAM_ST.scala 32:46]
  assign _GEN_3328 = 11'h57b == RADDR ? 11'h57b : _GEN_3327; // @[RAM_ST.scala 32:46]
  assign _GEN_3329 = 11'h57c == RADDR ? 11'h57c : _GEN_3328; // @[RAM_ST.scala 32:46]
  assign _GEN_3330 = 11'h57d == RADDR ? 11'h57d : _GEN_3329; // @[RAM_ST.scala 32:46]
  assign _GEN_3331 = 11'h57e == RADDR ? 11'h57e : _GEN_3330; // @[RAM_ST.scala 32:46]
  assign _GEN_3332 = 11'h57f == RADDR ? 11'h57f : _GEN_3331; // @[RAM_ST.scala 32:46]
  assign _GEN_3333 = 11'h580 == RADDR ? 11'h580 : _GEN_3332; // @[RAM_ST.scala 32:46]
  assign _GEN_3334 = 11'h581 == RADDR ? 11'h581 : _GEN_3333; // @[RAM_ST.scala 32:46]
  assign _GEN_3335 = 11'h582 == RADDR ? 11'h582 : _GEN_3334; // @[RAM_ST.scala 32:46]
  assign _GEN_3336 = 11'h583 == RADDR ? 11'h583 : _GEN_3335; // @[RAM_ST.scala 32:46]
  assign _GEN_3337 = 11'h584 == RADDR ? 11'h584 : _GEN_3336; // @[RAM_ST.scala 32:46]
  assign _GEN_3338 = 11'h585 == RADDR ? 11'h585 : _GEN_3337; // @[RAM_ST.scala 32:46]
  assign _GEN_3339 = 11'h586 == RADDR ? 11'h586 : _GEN_3338; // @[RAM_ST.scala 32:46]
  assign _GEN_3340 = 11'h587 == RADDR ? 11'h587 : _GEN_3339; // @[RAM_ST.scala 32:46]
  assign _GEN_3341 = 11'h588 == RADDR ? 11'h588 : _GEN_3340; // @[RAM_ST.scala 32:46]
  assign _GEN_3342 = 11'h589 == RADDR ? 11'h589 : _GEN_3341; // @[RAM_ST.scala 32:46]
  assign _GEN_3343 = 11'h58a == RADDR ? 11'h58a : _GEN_3342; // @[RAM_ST.scala 32:46]
  assign _GEN_3344 = 11'h58b == RADDR ? 11'h58b : _GEN_3343; // @[RAM_ST.scala 32:46]
  assign _GEN_3345 = 11'h58c == RADDR ? 11'h58c : _GEN_3344; // @[RAM_ST.scala 32:46]
  assign _GEN_3346 = 11'h58d == RADDR ? 11'h58d : _GEN_3345; // @[RAM_ST.scala 32:46]
  assign _GEN_3347 = 11'h58e == RADDR ? 11'h58e : _GEN_3346; // @[RAM_ST.scala 32:46]
  assign _GEN_3348 = 11'h58f == RADDR ? 11'h58f : _GEN_3347; // @[RAM_ST.scala 32:46]
  assign _GEN_3349 = 11'h590 == RADDR ? 11'h590 : _GEN_3348; // @[RAM_ST.scala 32:46]
  assign _GEN_3350 = 11'h591 == RADDR ? 11'h591 : _GEN_3349; // @[RAM_ST.scala 32:46]
  assign _GEN_3351 = 11'h592 == RADDR ? 11'h592 : _GEN_3350; // @[RAM_ST.scala 32:46]
  assign _GEN_3352 = 11'h593 == RADDR ? 11'h593 : _GEN_3351; // @[RAM_ST.scala 32:46]
  assign _GEN_3353 = 11'h594 == RADDR ? 11'h594 : _GEN_3352; // @[RAM_ST.scala 32:46]
  assign _GEN_3354 = 11'h595 == RADDR ? 11'h595 : _GEN_3353; // @[RAM_ST.scala 32:46]
  assign _GEN_3355 = 11'h596 == RADDR ? 11'h596 : _GEN_3354; // @[RAM_ST.scala 32:46]
  assign _GEN_3356 = 11'h597 == RADDR ? 11'h597 : _GEN_3355; // @[RAM_ST.scala 32:46]
  assign _GEN_3357 = 11'h598 == RADDR ? 11'h598 : _GEN_3356; // @[RAM_ST.scala 32:46]
  assign _GEN_3358 = 11'h599 == RADDR ? 11'h599 : _GEN_3357; // @[RAM_ST.scala 32:46]
  assign _GEN_3359 = 11'h59a == RADDR ? 11'h59a : _GEN_3358; // @[RAM_ST.scala 32:46]
  assign _GEN_3360 = 11'h59b == RADDR ? 11'h59b : _GEN_3359; // @[RAM_ST.scala 32:46]
  assign _GEN_3361 = 11'h59c == RADDR ? 11'h59c : _GEN_3360; // @[RAM_ST.scala 32:46]
  assign _GEN_3362 = 11'h59d == RADDR ? 11'h59d : _GEN_3361; // @[RAM_ST.scala 32:46]
  assign _GEN_3363 = 11'h59e == RADDR ? 11'h59e : _GEN_3362; // @[RAM_ST.scala 32:46]
  assign _GEN_3364 = 11'h59f == RADDR ? 11'h59f : _GEN_3363; // @[RAM_ST.scala 32:46]
  assign _GEN_3365 = 11'h5a0 == RADDR ? 11'h5a0 : _GEN_3364; // @[RAM_ST.scala 32:46]
  assign _GEN_3366 = 11'h5a1 == RADDR ? 11'h5a1 : _GEN_3365; // @[RAM_ST.scala 32:46]
  assign _GEN_3367 = 11'h5a2 == RADDR ? 11'h5a2 : _GEN_3366; // @[RAM_ST.scala 32:46]
  assign _GEN_3368 = 11'h5a3 == RADDR ? 11'h5a3 : _GEN_3367; // @[RAM_ST.scala 32:46]
  assign _GEN_3369 = 11'h5a4 == RADDR ? 11'h5a4 : _GEN_3368; // @[RAM_ST.scala 32:46]
  assign _GEN_3370 = 11'h5a5 == RADDR ? 11'h5a5 : _GEN_3369; // @[RAM_ST.scala 32:46]
  assign _GEN_3371 = 11'h5a6 == RADDR ? 11'h5a6 : _GEN_3370; // @[RAM_ST.scala 32:46]
  assign _GEN_3372 = 11'h5a7 == RADDR ? 11'h5a7 : _GEN_3371; // @[RAM_ST.scala 32:46]
  assign _GEN_3373 = 11'h5a8 == RADDR ? 11'h5a8 : _GEN_3372; // @[RAM_ST.scala 32:46]
  assign _GEN_3374 = 11'h5a9 == RADDR ? 11'h5a9 : _GEN_3373; // @[RAM_ST.scala 32:46]
  assign _GEN_3375 = 11'h5aa == RADDR ? 11'h5aa : _GEN_3374; // @[RAM_ST.scala 32:46]
  assign _GEN_3376 = 11'h5ab == RADDR ? 11'h5ab : _GEN_3375; // @[RAM_ST.scala 32:46]
  assign _GEN_3377 = 11'h5ac == RADDR ? 11'h5ac : _GEN_3376; // @[RAM_ST.scala 32:46]
  assign _GEN_3378 = 11'h5ad == RADDR ? 11'h5ad : _GEN_3377; // @[RAM_ST.scala 32:46]
  assign _GEN_3379 = 11'h5ae == RADDR ? 11'h5ae : _GEN_3378; // @[RAM_ST.scala 32:46]
  assign _GEN_3380 = 11'h5af == RADDR ? 11'h5af : _GEN_3379; // @[RAM_ST.scala 32:46]
  assign _GEN_3381 = 11'h5b0 == RADDR ? 11'h5b0 : _GEN_3380; // @[RAM_ST.scala 32:46]
  assign _GEN_3382 = 11'h5b1 == RADDR ? 11'h5b1 : _GEN_3381; // @[RAM_ST.scala 32:46]
  assign _GEN_3383 = 11'h5b2 == RADDR ? 11'h5b2 : _GEN_3382; // @[RAM_ST.scala 32:46]
  assign _GEN_3384 = 11'h5b3 == RADDR ? 11'h5b3 : _GEN_3383; // @[RAM_ST.scala 32:46]
  assign _GEN_3385 = 11'h5b4 == RADDR ? 11'h5b4 : _GEN_3384; // @[RAM_ST.scala 32:46]
  assign _GEN_3386 = 11'h5b5 == RADDR ? 11'h5b5 : _GEN_3385; // @[RAM_ST.scala 32:46]
  assign _GEN_3387 = 11'h5b6 == RADDR ? 11'h5b6 : _GEN_3386; // @[RAM_ST.scala 32:46]
  assign _GEN_3388 = 11'h5b7 == RADDR ? 11'h5b7 : _GEN_3387; // @[RAM_ST.scala 32:46]
  assign _GEN_3389 = 11'h5b8 == RADDR ? 11'h5b8 : _GEN_3388; // @[RAM_ST.scala 32:46]
  assign _GEN_3390 = 11'h5b9 == RADDR ? 11'h5b9 : _GEN_3389; // @[RAM_ST.scala 32:46]
  assign _GEN_3391 = 11'h5ba == RADDR ? 11'h5ba : _GEN_3390; // @[RAM_ST.scala 32:46]
  assign _GEN_3392 = 11'h5bb == RADDR ? 11'h5bb : _GEN_3391; // @[RAM_ST.scala 32:46]
  assign _GEN_3393 = 11'h5bc == RADDR ? 11'h5bc : _GEN_3392; // @[RAM_ST.scala 32:46]
  assign _GEN_3394 = 11'h5bd == RADDR ? 11'h5bd : _GEN_3393; // @[RAM_ST.scala 32:46]
  assign _GEN_3395 = 11'h5be == RADDR ? 11'h5be : _GEN_3394; // @[RAM_ST.scala 32:46]
  assign _GEN_3396 = 11'h5bf == RADDR ? 11'h5bf : _GEN_3395; // @[RAM_ST.scala 32:46]
  assign _GEN_3397 = 11'h5c0 == RADDR ? 11'h5c0 : _GEN_3396; // @[RAM_ST.scala 32:46]
  assign _GEN_3398 = 11'h5c1 == RADDR ? 11'h5c1 : _GEN_3397; // @[RAM_ST.scala 32:46]
  assign _GEN_3399 = 11'h5c2 == RADDR ? 11'h5c2 : _GEN_3398; // @[RAM_ST.scala 32:46]
  assign _GEN_3400 = 11'h5c3 == RADDR ? 11'h5c3 : _GEN_3399; // @[RAM_ST.scala 32:46]
  assign _GEN_3401 = 11'h5c4 == RADDR ? 11'h5c4 : _GEN_3400; // @[RAM_ST.scala 32:46]
  assign _GEN_3402 = 11'h5c5 == RADDR ? 11'h5c5 : _GEN_3401; // @[RAM_ST.scala 32:46]
  assign _GEN_3403 = 11'h5c6 == RADDR ? 11'h5c6 : _GEN_3402; // @[RAM_ST.scala 32:46]
  assign _GEN_3404 = 11'h5c7 == RADDR ? 11'h5c7 : _GEN_3403; // @[RAM_ST.scala 32:46]
  assign _GEN_3405 = 11'h5c8 == RADDR ? 11'h5c8 : _GEN_3404; // @[RAM_ST.scala 32:46]
  assign _GEN_3406 = 11'h5c9 == RADDR ? 11'h5c9 : _GEN_3405; // @[RAM_ST.scala 32:46]
  assign _GEN_3407 = 11'h5ca == RADDR ? 11'h5ca : _GEN_3406; // @[RAM_ST.scala 32:46]
  assign _GEN_3408 = 11'h5cb == RADDR ? 11'h5cb : _GEN_3407; // @[RAM_ST.scala 32:46]
  assign _GEN_3409 = 11'h5cc == RADDR ? 11'h5cc : _GEN_3408; // @[RAM_ST.scala 32:46]
  assign _GEN_3410 = 11'h5cd == RADDR ? 11'h5cd : _GEN_3409; // @[RAM_ST.scala 32:46]
  assign _GEN_3411 = 11'h5ce == RADDR ? 11'h5ce : _GEN_3410; // @[RAM_ST.scala 32:46]
  assign _GEN_3412 = 11'h5cf == RADDR ? 11'h5cf : _GEN_3411; // @[RAM_ST.scala 32:46]
  assign _GEN_3413 = 11'h5d0 == RADDR ? 11'h5d0 : _GEN_3412; // @[RAM_ST.scala 32:46]
  assign _GEN_3414 = 11'h5d1 == RADDR ? 11'h5d1 : _GEN_3413; // @[RAM_ST.scala 32:46]
  assign _GEN_3415 = 11'h5d2 == RADDR ? 11'h5d2 : _GEN_3414; // @[RAM_ST.scala 32:46]
  assign _GEN_3416 = 11'h5d3 == RADDR ? 11'h5d3 : _GEN_3415; // @[RAM_ST.scala 32:46]
  assign _GEN_3417 = 11'h5d4 == RADDR ? 11'h5d4 : _GEN_3416; // @[RAM_ST.scala 32:46]
  assign _GEN_3418 = 11'h5d5 == RADDR ? 11'h5d5 : _GEN_3417; // @[RAM_ST.scala 32:46]
  assign _GEN_3419 = 11'h5d6 == RADDR ? 11'h5d6 : _GEN_3418; // @[RAM_ST.scala 32:46]
  assign _GEN_3420 = 11'h5d7 == RADDR ? 11'h5d7 : _GEN_3419; // @[RAM_ST.scala 32:46]
  assign _GEN_3421 = 11'h5d8 == RADDR ? 11'h5d8 : _GEN_3420; // @[RAM_ST.scala 32:46]
  assign _GEN_3422 = 11'h5d9 == RADDR ? 11'h5d9 : _GEN_3421; // @[RAM_ST.scala 32:46]
  assign _GEN_3423 = 11'h5da == RADDR ? 11'h5da : _GEN_3422; // @[RAM_ST.scala 32:46]
  assign _GEN_3424 = 11'h5db == RADDR ? 11'h5db : _GEN_3423; // @[RAM_ST.scala 32:46]
  assign _GEN_3425 = 11'h5dc == RADDR ? 11'h5dc : _GEN_3424; // @[RAM_ST.scala 32:46]
  assign _GEN_3426 = 11'h5dd == RADDR ? 11'h5dd : _GEN_3425; // @[RAM_ST.scala 32:46]
  assign _GEN_3427 = 11'h5de == RADDR ? 11'h5de : _GEN_3426; // @[RAM_ST.scala 32:46]
  assign _GEN_3428 = 11'h5df == RADDR ? 11'h5df : _GEN_3427; // @[RAM_ST.scala 32:46]
  assign _GEN_3429 = 11'h5e0 == RADDR ? 11'h5e0 : _GEN_3428; // @[RAM_ST.scala 32:46]
  assign _GEN_3430 = 11'h5e1 == RADDR ? 11'h5e1 : _GEN_3429; // @[RAM_ST.scala 32:46]
  assign _GEN_3431 = 11'h5e2 == RADDR ? 11'h5e2 : _GEN_3430; // @[RAM_ST.scala 32:46]
  assign _GEN_3432 = 11'h5e3 == RADDR ? 11'h5e3 : _GEN_3431; // @[RAM_ST.scala 32:46]
  assign _GEN_3433 = 11'h5e4 == RADDR ? 11'h5e4 : _GEN_3432; // @[RAM_ST.scala 32:46]
  assign _GEN_3434 = 11'h5e5 == RADDR ? 11'h5e5 : _GEN_3433; // @[RAM_ST.scala 32:46]
  assign _GEN_3435 = 11'h5e6 == RADDR ? 11'h5e6 : _GEN_3434; // @[RAM_ST.scala 32:46]
  assign _GEN_3436 = 11'h5e7 == RADDR ? 11'h5e7 : _GEN_3435; // @[RAM_ST.scala 32:46]
  assign _GEN_3437 = 11'h5e8 == RADDR ? 11'h5e8 : _GEN_3436; // @[RAM_ST.scala 32:46]
  assign _GEN_3438 = 11'h5e9 == RADDR ? 11'h5e9 : _GEN_3437; // @[RAM_ST.scala 32:46]
  assign _GEN_3439 = 11'h5ea == RADDR ? 11'h5ea : _GEN_3438; // @[RAM_ST.scala 32:46]
  assign _GEN_3440 = 11'h5eb == RADDR ? 11'h5eb : _GEN_3439; // @[RAM_ST.scala 32:46]
  assign _GEN_3441 = 11'h5ec == RADDR ? 11'h5ec : _GEN_3440; // @[RAM_ST.scala 32:46]
  assign _GEN_3442 = 11'h5ed == RADDR ? 11'h5ed : _GEN_3441; // @[RAM_ST.scala 32:46]
  assign _GEN_3443 = 11'h5ee == RADDR ? 11'h5ee : _GEN_3442; // @[RAM_ST.scala 32:46]
  assign _GEN_3444 = 11'h5ef == RADDR ? 11'h5ef : _GEN_3443; // @[RAM_ST.scala 32:46]
  assign _GEN_3445 = 11'h5f0 == RADDR ? 11'h5f0 : _GEN_3444; // @[RAM_ST.scala 32:46]
  assign _GEN_3446 = 11'h5f1 == RADDR ? 11'h5f1 : _GEN_3445; // @[RAM_ST.scala 32:46]
  assign _GEN_3447 = 11'h5f2 == RADDR ? 11'h5f2 : _GEN_3446; // @[RAM_ST.scala 32:46]
  assign _GEN_3448 = 11'h5f3 == RADDR ? 11'h5f3 : _GEN_3447; // @[RAM_ST.scala 32:46]
  assign _GEN_3449 = 11'h5f4 == RADDR ? 11'h5f4 : _GEN_3448; // @[RAM_ST.scala 32:46]
  assign _GEN_3450 = 11'h5f5 == RADDR ? 11'h5f5 : _GEN_3449; // @[RAM_ST.scala 32:46]
  assign _GEN_3451 = 11'h5f6 == RADDR ? 11'h5f6 : _GEN_3450; // @[RAM_ST.scala 32:46]
  assign _GEN_3452 = 11'h5f7 == RADDR ? 11'h5f7 : _GEN_3451; // @[RAM_ST.scala 32:46]
  assign _GEN_3453 = 11'h5f8 == RADDR ? 11'h5f8 : _GEN_3452; // @[RAM_ST.scala 32:46]
  assign _GEN_3454 = 11'h5f9 == RADDR ? 11'h5f9 : _GEN_3453; // @[RAM_ST.scala 32:46]
  assign _GEN_3455 = 11'h5fa == RADDR ? 11'h5fa : _GEN_3454; // @[RAM_ST.scala 32:46]
  assign _GEN_3456 = 11'h5fb == RADDR ? 11'h5fb : _GEN_3455; // @[RAM_ST.scala 32:46]
  assign _GEN_3457 = 11'h5fc == RADDR ? 11'h5fc : _GEN_3456; // @[RAM_ST.scala 32:46]
  assign _GEN_3458 = 11'h5fd == RADDR ? 11'h5fd : _GEN_3457; // @[RAM_ST.scala 32:46]
  assign _GEN_3459 = 11'h5fe == RADDR ? 11'h5fe : _GEN_3458; // @[RAM_ST.scala 32:46]
  assign _GEN_3460 = 11'h5ff == RADDR ? 11'h5ff : _GEN_3459; // @[RAM_ST.scala 32:46]
  assign _GEN_3461 = 11'h600 == RADDR ? 11'h600 : _GEN_3460; // @[RAM_ST.scala 32:46]
  assign _GEN_3462 = 11'h601 == RADDR ? 11'h601 : _GEN_3461; // @[RAM_ST.scala 32:46]
  assign _GEN_3463 = 11'h602 == RADDR ? 11'h602 : _GEN_3462; // @[RAM_ST.scala 32:46]
  assign _GEN_3464 = 11'h603 == RADDR ? 11'h603 : _GEN_3463; // @[RAM_ST.scala 32:46]
  assign _GEN_3465 = 11'h604 == RADDR ? 11'h604 : _GEN_3464; // @[RAM_ST.scala 32:46]
  assign _GEN_3466 = 11'h605 == RADDR ? 11'h605 : _GEN_3465; // @[RAM_ST.scala 32:46]
  assign _GEN_3467 = 11'h606 == RADDR ? 11'h606 : _GEN_3466; // @[RAM_ST.scala 32:46]
  assign _GEN_3468 = 11'h607 == RADDR ? 11'h607 : _GEN_3467; // @[RAM_ST.scala 32:46]
  assign _GEN_3469 = 11'h608 == RADDR ? 11'h608 : _GEN_3468; // @[RAM_ST.scala 32:46]
  assign _GEN_3470 = 11'h609 == RADDR ? 11'h609 : _GEN_3469; // @[RAM_ST.scala 32:46]
  assign _GEN_3471 = 11'h60a == RADDR ? 11'h60a : _GEN_3470; // @[RAM_ST.scala 32:46]
  assign _GEN_3472 = 11'h60b == RADDR ? 11'h60b : _GEN_3471; // @[RAM_ST.scala 32:46]
  assign _GEN_3473 = 11'h60c == RADDR ? 11'h60c : _GEN_3472; // @[RAM_ST.scala 32:46]
  assign _GEN_3474 = 11'h60d == RADDR ? 11'h60d : _GEN_3473; // @[RAM_ST.scala 32:46]
  assign _GEN_3475 = 11'h60e == RADDR ? 11'h60e : _GEN_3474; // @[RAM_ST.scala 32:46]
  assign _GEN_3476 = 11'h60f == RADDR ? 11'h60f : _GEN_3475; // @[RAM_ST.scala 32:46]
  assign _GEN_3477 = 11'h610 == RADDR ? 11'h610 : _GEN_3476; // @[RAM_ST.scala 32:46]
  assign _GEN_3478 = 11'h611 == RADDR ? 11'h611 : _GEN_3477; // @[RAM_ST.scala 32:46]
  assign _GEN_3479 = 11'h612 == RADDR ? 11'h612 : _GEN_3478; // @[RAM_ST.scala 32:46]
  assign _GEN_3480 = 11'h613 == RADDR ? 11'h613 : _GEN_3479; // @[RAM_ST.scala 32:46]
  assign _GEN_3481 = 11'h614 == RADDR ? 11'h614 : _GEN_3480; // @[RAM_ST.scala 32:46]
  assign _GEN_3482 = 11'h615 == RADDR ? 11'h615 : _GEN_3481; // @[RAM_ST.scala 32:46]
  assign _GEN_3483 = 11'h616 == RADDR ? 11'h616 : _GEN_3482; // @[RAM_ST.scala 32:46]
  assign _GEN_3484 = 11'h617 == RADDR ? 11'h617 : _GEN_3483; // @[RAM_ST.scala 32:46]
  assign _GEN_3485 = 11'h618 == RADDR ? 11'h618 : _GEN_3484; // @[RAM_ST.scala 32:46]
  assign _GEN_3486 = 11'h619 == RADDR ? 11'h619 : _GEN_3485; // @[RAM_ST.scala 32:46]
  assign _GEN_3487 = 11'h61a == RADDR ? 11'h61a : _GEN_3486; // @[RAM_ST.scala 32:46]
  assign _GEN_3488 = 11'h61b == RADDR ? 11'h61b : _GEN_3487; // @[RAM_ST.scala 32:46]
  assign _GEN_3489 = 11'h61c == RADDR ? 11'h61c : _GEN_3488; // @[RAM_ST.scala 32:46]
  assign _GEN_3490 = 11'h61d == RADDR ? 11'h61d : _GEN_3489; // @[RAM_ST.scala 32:46]
  assign _GEN_3491 = 11'h61e == RADDR ? 11'h61e : _GEN_3490; // @[RAM_ST.scala 32:46]
  assign _GEN_3492 = 11'h61f == RADDR ? 11'h61f : _GEN_3491; // @[RAM_ST.scala 32:46]
  assign _GEN_3493 = 11'h620 == RADDR ? 11'h620 : _GEN_3492; // @[RAM_ST.scala 32:46]
  assign _GEN_3494 = 11'h621 == RADDR ? 11'h621 : _GEN_3493; // @[RAM_ST.scala 32:46]
  assign _GEN_3495 = 11'h622 == RADDR ? 11'h622 : _GEN_3494; // @[RAM_ST.scala 32:46]
  assign _GEN_3496 = 11'h623 == RADDR ? 11'h623 : _GEN_3495; // @[RAM_ST.scala 32:46]
  assign _GEN_3497 = 11'h624 == RADDR ? 11'h624 : _GEN_3496; // @[RAM_ST.scala 32:46]
  assign _GEN_3498 = 11'h625 == RADDR ? 11'h625 : _GEN_3497; // @[RAM_ST.scala 32:46]
  assign _GEN_3499 = 11'h626 == RADDR ? 11'h626 : _GEN_3498; // @[RAM_ST.scala 32:46]
  assign _GEN_3500 = 11'h627 == RADDR ? 11'h627 : _GEN_3499; // @[RAM_ST.scala 32:46]
  assign _GEN_3501 = 11'h628 == RADDR ? 11'h628 : _GEN_3500; // @[RAM_ST.scala 32:46]
  assign _GEN_3502 = 11'h629 == RADDR ? 11'h629 : _GEN_3501; // @[RAM_ST.scala 32:46]
  assign _GEN_3503 = 11'h62a == RADDR ? 11'h62a : _GEN_3502; // @[RAM_ST.scala 32:46]
  assign _GEN_3504 = 11'h62b == RADDR ? 11'h62b : _GEN_3503; // @[RAM_ST.scala 32:46]
  assign _GEN_3505 = 11'h62c == RADDR ? 11'h62c : _GEN_3504; // @[RAM_ST.scala 32:46]
  assign _GEN_3506 = 11'h62d == RADDR ? 11'h62d : _GEN_3505; // @[RAM_ST.scala 32:46]
  assign _GEN_3507 = 11'h62e == RADDR ? 11'h62e : _GEN_3506; // @[RAM_ST.scala 32:46]
  assign _GEN_3508 = 11'h62f == RADDR ? 11'h62f : _GEN_3507; // @[RAM_ST.scala 32:46]
  assign _GEN_3509 = 11'h630 == RADDR ? 11'h630 : _GEN_3508; // @[RAM_ST.scala 32:46]
  assign _GEN_3510 = 11'h631 == RADDR ? 11'h631 : _GEN_3509; // @[RAM_ST.scala 32:46]
  assign _GEN_3511 = 11'h632 == RADDR ? 11'h632 : _GEN_3510; // @[RAM_ST.scala 32:46]
  assign _GEN_3512 = 11'h633 == RADDR ? 11'h633 : _GEN_3511; // @[RAM_ST.scala 32:46]
  assign _GEN_3513 = 11'h634 == RADDR ? 11'h634 : _GEN_3512; // @[RAM_ST.scala 32:46]
  assign _GEN_3514 = 11'h635 == RADDR ? 11'h635 : _GEN_3513; // @[RAM_ST.scala 32:46]
  assign _GEN_3515 = 11'h636 == RADDR ? 11'h636 : _GEN_3514; // @[RAM_ST.scala 32:46]
  assign _GEN_3516 = 11'h637 == RADDR ? 11'h637 : _GEN_3515; // @[RAM_ST.scala 32:46]
  assign _GEN_3517 = 11'h638 == RADDR ? 11'h638 : _GEN_3516; // @[RAM_ST.scala 32:46]
  assign _GEN_3518 = 11'h639 == RADDR ? 11'h639 : _GEN_3517; // @[RAM_ST.scala 32:46]
  assign _GEN_3519 = 11'h63a == RADDR ? 11'h63a : _GEN_3518; // @[RAM_ST.scala 32:46]
  assign _GEN_3520 = 11'h63b == RADDR ? 11'h63b : _GEN_3519; // @[RAM_ST.scala 32:46]
  assign _GEN_3521 = 11'h63c == RADDR ? 11'h63c : _GEN_3520; // @[RAM_ST.scala 32:46]
  assign _GEN_3522 = 11'h63d == RADDR ? 11'h63d : _GEN_3521; // @[RAM_ST.scala 32:46]
  assign _GEN_3523 = 11'h63e == RADDR ? 11'h63e : _GEN_3522; // @[RAM_ST.scala 32:46]
  assign _GEN_3524 = 11'h63f == RADDR ? 11'h63f : _GEN_3523; // @[RAM_ST.scala 32:46]
  assign _GEN_3525 = 11'h640 == RADDR ? 11'h640 : _GEN_3524; // @[RAM_ST.scala 32:46]
  assign _GEN_3526 = 11'h641 == RADDR ? 11'h641 : _GEN_3525; // @[RAM_ST.scala 32:46]
  assign _GEN_3527 = 11'h642 == RADDR ? 11'h642 : _GEN_3526; // @[RAM_ST.scala 32:46]
  assign _GEN_3528 = 11'h643 == RADDR ? 11'h643 : _GEN_3527; // @[RAM_ST.scala 32:46]
  assign _GEN_3529 = 11'h644 == RADDR ? 11'h644 : _GEN_3528; // @[RAM_ST.scala 32:46]
  assign _GEN_3530 = 11'h645 == RADDR ? 11'h645 : _GEN_3529; // @[RAM_ST.scala 32:46]
  assign _GEN_3531 = 11'h646 == RADDR ? 11'h646 : _GEN_3530; // @[RAM_ST.scala 32:46]
  assign _GEN_3532 = 11'h647 == RADDR ? 11'h647 : _GEN_3531; // @[RAM_ST.scala 32:46]
  assign _GEN_3533 = 11'h648 == RADDR ? 11'h648 : _GEN_3532; // @[RAM_ST.scala 32:46]
  assign _GEN_3534 = 11'h649 == RADDR ? 11'h649 : _GEN_3533; // @[RAM_ST.scala 32:46]
  assign _GEN_3535 = 11'h64a == RADDR ? 11'h64a : _GEN_3534; // @[RAM_ST.scala 32:46]
  assign _GEN_3536 = 11'h64b == RADDR ? 11'h64b : _GEN_3535; // @[RAM_ST.scala 32:46]
  assign _GEN_3537 = 11'h64c == RADDR ? 11'h64c : _GEN_3536; // @[RAM_ST.scala 32:46]
  assign _GEN_3538 = 11'h64d == RADDR ? 11'h64d : _GEN_3537; // @[RAM_ST.scala 32:46]
  assign _GEN_3539 = 11'h64e == RADDR ? 11'h64e : _GEN_3538; // @[RAM_ST.scala 32:46]
  assign _GEN_3540 = 11'h64f == RADDR ? 11'h64f : _GEN_3539; // @[RAM_ST.scala 32:46]
  assign _GEN_3541 = 11'h650 == RADDR ? 11'h650 : _GEN_3540; // @[RAM_ST.scala 32:46]
  assign _GEN_3542 = 11'h651 == RADDR ? 11'h651 : _GEN_3541; // @[RAM_ST.scala 32:46]
  assign _GEN_3543 = 11'h652 == RADDR ? 11'h652 : _GEN_3542; // @[RAM_ST.scala 32:46]
  assign _GEN_3544 = 11'h653 == RADDR ? 11'h653 : _GEN_3543; // @[RAM_ST.scala 32:46]
  assign _GEN_3545 = 11'h654 == RADDR ? 11'h654 : _GEN_3544; // @[RAM_ST.scala 32:46]
  assign _GEN_3546 = 11'h655 == RADDR ? 11'h655 : _GEN_3545; // @[RAM_ST.scala 32:46]
  assign _GEN_3547 = 11'h656 == RADDR ? 11'h656 : _GEN_3546; // @[RAM_ST.scala 32:46]
  assign _GEN_3548 = 11'h657 == RADDR ? 11'h657 : _GEN_3547; // @[RAM_ST.scala 32:46]
  assign _GEN_3549 = 11'h658 == RADDR ? 11'h658 : _GEN_3548; // @[RAM_ST.scala 32:46]
  assign _GEN_3550 = 11'h659 == RADDR ? 11'h659 : _GEN_3549; // @[RAM_ST.scala 32:46]
  assign _GEN_3551 = 11'h65a == RADDR ? 11'h65a : _GEN_3550; // @[RAM_ST.scala 32:46]
  assign _GEN_3552 = 11'h65b == RADDR ? 11'h65b : _GEN_3551; // @[RAM_ST.scala 32:46]
  assign _GEN_3553 = 11'h65c == RADDR ? 11'h65c : _GEN_3552; // @[RAM_ST.scala 32:46]
  assign _GEN_3554 = 11'h65d == RADDR ? 11'h65d : _GEN_3553; // @[RAM_ST.scala 32:46]
  assign _GEN_3555 = 11'h65e == RADDR ? 11'h65e : _GEN_3554; // @[RAM_ST.scala 32:46]
  assign _GEN_3556 = 11'h65f == RADDR ? 11'h65f : _GEN_3555; // @[RAM_ST.scala 32:46]
  assign _GEN_3557 = 11'h660 == RADDR ? 11'h660 : _GEN_3556; // @[RAM_ST.scala 32:46]
  assign _GEN_3558 = 11'h661 == RADDR ? 11'h661 : _GEN_3557; // @[RAM_ST.scala 32:46]
  assign _GEN_3559 = 11'h662 == RADDR ? 11'h662 : _GEN_3558; // @[RAM_ST.scala 32:46]
  assign _GEN_3560 = 11'h663 == RADDR ? 11'h663 : _GEN_3559; // @[RAM_ST.scala 32:46]
  assign _GEN_3561 = 11'h664 == RADDR ? 11'h664 : _GEN_3560; // @[RAM_ST.scala 32:46]
  assign _GEN_3562 = 11'h665 == RADDR ? 11'h665 : _GEN_3561; // @[RAM_ST.scala 32:46]
  assign _GEN_3563 = 11'h666 == RADDR ? 11'h666 : _GEN_3562; // @[RAM_ST.scala 32:46]
  assign _GEN_3564 = 11'h667 == RADDR ? 11'h667 : _GEN_3563; // @[RAM_ST.scala 32:46]
  assign _GEN_3565 = 11'h668 == RADDR ? 11'h668 : _GEN_3564; // @[RAM_ST.scala 32:46]
  assign _GEN_3566 = 11'h669 == RADDR ? 11'h669 : _GEN_3565; // @[RAM_ST.scala 32:46]
  assign _GEN_3567 = 11'h66a == RADDR ? 11'h66a : _GEN_3566; // @[RAM_ST.scala 32:46]
  assign _GEN_3568 = 11'h66b == RADDR ? 11'h66b : _GEN_3567; // @[RAM_ST.scala 32:46]
  assign _GEN_3569 = 11'h66c == RADDR ? 11'h66c : _GEN_3568; // @[RAM_ST.scala 32:46]
  assign _GEN_3570 = 11'h66d == RADDR ? 11'h66d : _GEN_3569; // @[RAM_ST.scala 32:46]
  assign _GEN_3571 = 11'h66e == RADDR ? 11'h66e : _GEN_3570; // @[RAM_ST.scala 32:46]
  assign _GEN_3572 = 11'h66f == RADDR ? 11'h66f : _GEN_3571; // @[RAM_ST.scala 32:46]
  assign _GEN_3573 = 11'h670 == RADDR ? 11'h670 : _GEN_3572; // @[RAM_ST.scala 32:46]
  assign _GEN_3574 = 11'h671 == RADDR ? 11'h671 : _GEN_3573; // @[RAM_ST.scala 32:46]
  assign _GEN_3575 = 11'h672 == RADDR ? 11'h672 : _GEN_3574; // @[RAM_ST.scala 32:46]
  assign _GEN_3576 = 11'h673 == RADDR ? 11'h673 : _GEN_3575; // @[RAM_ST.scala 32:46]
  assign _GEN_3577 = 11'h674 == RADDR ? 11'h674 : _GEN_3576; // @[RAM_ST.scala 32:46]
  assign _GEN_3578 = 11'h675 == RADDR ? 11'h675 : _GEN_3577; // @[RAM_ST.scala 32:46]
  assign _GEN_3579 = 11'h676 == RADDR ? 11'h676 : _GEN_3578; // @[RAM_ST.scala 32:46]
  assign _GEN_3580 = 11'h677 == RADDR ? 11'h677 : _GEN_3579; // @[RAM_ST.scala 32:46]
  assign _GEN_3581 = 11'h678 == RADDR ? 11'h678 : _GEN_3580; // @[RAM_ST.scala 32:46]
  assign _GEN_3582 = 11'h679 == RADDR ? 11'h679 : _GEN_3581; // @[RAM_ST.scala 32:46]
  assign _GEN_3583 = 11'h67a == RADDR ? 11'h67a : _GEN_3582; // @[RAM_ST.scala 32:46]
  assign _GEN_3584 = 11'h67b == RADDR ? 11'h67b : _GEN_3583; // @[RAM_ST.scala 32:46]
  assign _GEN_3585 = 11'h67c == RADDR ? 11'h67c : _GEN_3584; // @[RAM_ST.scala 32:46]
  assign _GEN_3586 = 11'h67d == RADDR ? 11'h67d : _GEN_3585; // @[RAM_ST.scala 32:46]
  assign _GEN_3587 = 11'h67e == RADDR ? 11'h67e : _GEN_3586; // @[RAM_ST.scala 32:46]
  assign _GEN_3588 = 11'h67f == RADDR ? 11'h67f : _GEN_3587; // @[RAM_ST.scala 32:46]
  assign _GEN_3589 = 11'h680 == RADDR ? 11'h680 : _GEN_3588; // @[RAM_ST.scala 32:46]
  assign _GEN_3590 = 11'h681 == RADDR ? 11'h681 : _GEN_3589; // @[RAM_ST.scala 32:46]
  assign _GEN_3591 = 11'h682 == RADDR ? 11'h682 : _GEN_3590; // @[RAM_ST.scala 32:46]
  assign _GEN_3592 = 11'h683 == RADDR ? 11'h683 : _GEN_3591; // @[RAM_ST.scala 32:46]
  assign _GEN_3593 = 11'h684 == RADDR ? 11'h684 : _GEN_3592; // @[RAM_ST.scala 32:46]
  assign _GEN_3594 = 11'h685 == RADDR ? 11'h685 : _GEN_3593; // @[RAM_ST.scala 32:46]
  assign _GEN_3595 = 11'h686 == RADDR ? 11'h686 : _GEN_3594; // @[RAM_ST.scala 32:46]
  assign _GEN_3596 = 11'h687 == RADDR ? 11'h687 : _GEN_3595; // @[RAM_ST.scala 32:46]
  assign _GEN_3597 = 11'h688 == RADDR ? 11'h688 : _GEN_3596; // @[RAM_ST.scala 32:46]
  assign _GEN_3598 = 11'h689 == RADDR ? 11'h689 : _GEN_3597; // @[RAM_ST.scala 32:46]
  assign _GEN_3599 = 11'h68a == RADDR ? 11'h68a : _GEN_3598; // @[RAM_ST.scala 32:46]
  assign _GEN_3600 = 11'h68b == RADDR ? 11'h68b : _GEN_3599; // @[RAM_ST.scala 32:46]
  assign _GEN_3601 = 11'h68c == RADDR ? 11'h68c : _GEN_3600; // @[RAM_ST.scala 32:46]
  assign _GEN_3602 = 11'h68d == RADDR ? 11'h68d : _GEN_3601; // @[RAM_ST.scala 32:46]
  assign _GEN_3603 = 11'h68e == RADDR ? 11'h68e : _GEN_3602; // @[RAM_ST.scala 32:46]
  assign _GEN_3604 = 11'h68f == RADDR ? 11'h68f : _GEN_3603; // @[RAM_ST.scala 32:46]
  assign _GEN_3605 = 11'h690 == RADDR ? 11'h690 : _GEN_3604; // @[RAM_ST.scala 32:46]
  assign _GEN_3606 = 11'h691 == RADDR ? 11'h691 : _GEN_3605; // @[RAM_ST.scala 32:46]
  assign _GEN_3607 = 11'h692 == RADDR ? 11'h692 : _GEN_3606; // @[RAM_ST.scala 32:46]
  assign _GEN_3608 = 11'h693 == RADDR ? 11'h693 : _GEN_3607; // @[RAM_ST.scala 32:46]
  assign _GEN_3609 = 11'h694 == RADDR ? 11'h694 : _GEN_3608; // @[RAM_ST.scala 32:46]
  assign _GEN_3610 = 11'h695 == RADDR ? 11'h695 : _GEN_3609; // @[RAM_ST.scala 32:46]
  assign _GEN_3611 = 11'h696 == RADDR ? 11'h696 : _GEN_3610; // @[RAM_ST.scala 32:46]
  assign _GEN_3612 = 11'h697 == RADDR ? 11'h697 : _GEN_3611; // @[RAM_ST.scala 32:46]
  assign _GEN_3613 = 11'h698 == RADDR ? 11'h698 : _GEN_3612; // @[RAM_ST.scala 32:46]
  assign _GEN_3614 = 11'h699 == RADDR ? 11'h699 : _GEN_3613; // @[RAM_ST.scala 32:46]
  assign _GEN_3615 = 11'h69a == RADDR ? 11'h69a : _GEN_3614; // @[RAM_ST.scala 32:46]
  assign _GEN_3616 = 11'h69b == RADDR ? 11'h69b : _GEN_3615; // @[RAM_ST.scala 32:46]
  assign _GEN_3617 = 11'h69c == RADDR ? 11'h69c : _GEN_3616; // @[RAM_ST.scala 32:46]
  assign _GEN_3618 = 11'h69d == RADDR ? 11'h69d : _GEN_3617; // @[RAM_ST.scala 32:46]
  assign _GEN_3619 = 11'h69e == RADDR ? 11'h69e : _GEN_3618; // @[RAM_ST.scala 32:46]
  assign _GEN_3620 = 11'h69f == RADDR ? 11'h69f : _GEN_3619; // @[RAM_ST.scala 32:46]
  assign _GEN_3621 = 11'h6a0 == RADDR ? 11'h6a0 : _GEN_3620; // @[RAM_ST.scala 32:46]
  assign _GEN_3622 = 11'h6a1 == RADDR ? 11'h6a1 : _GEN_3621; // @[RAM_ST.scala 32:46]
  assign _GEN_3623 = 11'h6a2 == RADDR ? 11'h6a2 : _GEN_3622; // @[RAM_ST.scala 32:46]
  assign _GEN_3624 = 11'h6a3 == RADDR ? 11'h6a3 : _GEN_3623; // @[RAM_ST.scala 32:46]
  assign _GEN_3625 = 11'h6a4 == RADDR ? 11'h6a4 : _GEN_3624; // @[RAM_ST.scala 32:46]
  assign _GEN_3626 = 11'h6a5 == RADDR ? 11'h6a5 : _GEN_3625; // @[RAM_ST.scala 32:46]
  assign _GEN_3627 = 11'h6a6 == RADDR ? 11'h6a6 : _GEN_3626; // @[RAM_ST.scala 32:46]
  assign _GEN_3628 = 11'h6a7 == RADDR ? 11'h6a7 : _GEN_3627; // @[RAM_ST.scala 32:46]
  assign _GEN_3629 = 11'h6a8 == RADDR ? 11'h6a8 : _GEN_3628; // @[RAM_ST.scala 32:46]
  assign _GEN_3630 = 11'h6a9 == RADDR ? 11'h6a9 : _GEN_3629; // @[RAM_ST.scala 32:46]
  assign _GEN_3631 = 11'h6aa == RADDR ? 11'h6aa : _GEN_3630; // @[RAM_ST.scala 32:46]
  assign _GEN_3632 = 11'h6ab == RADDR ? 11'h6ab : _GEN_3631; // @[RAM_ST.scala 32:46]
  assign _GEN_3633 = 11'h6ac == RADDR ? 11'h6ac : _GEN_3632; // @[RAM_ST.scala 32:46]
  assign _GEN_3634 = 11'h6ad == RADDR ? 11'h6ad : _GEN_3633; // @[RAM_ST.scala 32:46]
  assign _GEN_3635 = 11'h6ae == RADDR ? 11'h6ae : _GEN_3634; // @[RAM_ST.scala 32:46]
  assign _GEN_3636 = 11'h6af == RADDR ? 11'h6af : _GEN_3635; // @[RAM_ST.scala 32:46]
  assign _GEN_3637 = 11'h6b0 == RADDR ? 11'h6b0 : _GEN_3636; // @[RAM_ST.scala 32:46]
  assign _GEN_3638 = 11'h6b1 == RADDR ? 11'h6b1 : _GEN_3637; // @[RAM_ST.scala 32:46]
  assign _GEN_3639 = 11'h6b2 == RADDR ? 11'h6b2 : _GEN_3638; // @[RAM_ST.scala 32:46]
  assign _GEN_3640 = 11'h6b3 == RADDR ? 11'h6b3 : _GEN_3639; // @[RAM_ST.scala 32:46]
  assign _GEN_3641 = 11'h6b4 == RADDR ? 11'h6b4 : _GEN_3640; // @[RAM_ST.scala 32:46]
  assign _GEN_3642 = 11'h6b5 == RADDR ? 11'h6b5 : _GEN_3641; // @[RAM_ST.scala 32:46]
  assign _GEN_3643 = 11'h6b6 == RADDR ? 11'h6b6 : _GEN_3642; // @[RAM_ST.scala 32:46]
  assign _GEN_3644 = 11'h6b7 == RADDR ? 11'h6b7 : _GEN_3643; // @[RAM_ST.scala 32:46]
  assign _GEN_3645 = 11'h6b8 == RADDR ? 11'h6b8 : _GEN_3644; // @[RAM_ST.scala 32:46]
  assign _GEN_3646 = 11'h6b9 == RADDR ? 11'h6b9 : _GEN_3645; // @[RAM_ST.scala 32:46]
  assign _GEN_3647 = 11'h6ba == RADDR ? 11'h6ba : _GEN_3646; // @[RAM_ST.scala 32:46]
  assign _GEN_3648 = 11'h6bb == RADDR ? 11'h6bb : _GEN_3647; // @[RAM_ST.scala 32:46]
  assign _GEN_3649 = 11'h6bc == RADDR ? 11'h6bc : _GEN_3648; // @[RAM_ST.scala 32:46]
  assign _GEN_3650 = 11'h6bd == RADDR ? 11'h6bd : _GEN_3649; // @[RAM_ST.scala 32:46]
  assign _GEN_3651 = 11'h6be == RADDR ? 11'h6be : _GEN_3650; // @[RAM_ST.scala 32:46]
  assign _GEN_3652 = 11'h6bf == RADDR ? 11'h6bf : _GEN_3651; // @[RAM_ST.scala 32:46]
  assign _GEN_3653 = 11'h6c0 == RADDR ? 11'h6c0 : _GEN_3652; // @[RAM_ST.scala 32:46]
  assign _GEN_3654 = 11'h6c1 == RADDR ? 11'h6c1 : _GEN_3653; // @[RAM_ST.scala 32:46]
  assign _GEN_3655 = 11'h6c2 == RADDR ? 11'h6c2 : _GEN_3654; // @[RAM_ST.scala 32:46]
  assign _GEN_3656 = 11'h6c3 == RADDR ? 11'h6c3 : _GEN_3655; // @[RAM_ST.scala 32:46]
  assign _GEN_3657 = 11'h6c4 == RADDR ? 11'h6c4 : _GEN_3656; // @[RAM_ST.scala 32:46]
  assign _GEN_3658 = 11'h6c5 == RADDR ? 11'h6c5 : _GEN_3657; // @[RAM_ST.scala 32:46]
  assign _GEN_3659 = 11'h6c6 == RADDR ? 11'h6c6 : _GEN_3658; // @[RAM_ST.scala 32:46]
  assign _GEN_3660 = 11'h6c7 == RADDR ? 11'h6c7 : _GEN_3659; // @[RAM_ST.scala 32:46]
  assign _GEN_3661 = 11'h6c8 == RADDR ? 11'h6c8 : _GEN_3660; // @[RAM_ST.scala 32:46]
  assign _GEN_3662 = 11'h6c9 == RADDR ? 11'h6c9 : _GEN_3661; // @[RAM_ST.scala 32:46]
  assign _GEN_3663 = 11'h6ca == RADDR ? 11'h6ca : _GEN_3662; // @[RAM_ST.scala 32:46]
  assign _GEN_3664 = 11'h6cb == RADDR ? 11'h6cb : _GEN_3663; // @[RAM_ST.scala 32:46]
  assign _GEN_3665 = 11'h6cc == RADDR ? 11'h6cc : _GEN_3664; // @[RAM_ST.scala 32:46]
  assign _GEN_3666 = 11'h6cd == RADDR ? 11'h6cd : _GEN_3665; // @[RAM_ST.scala 32:46]
  assign _GEN_3667 = 11'h6ce == RADDR ? 11'h6ce : _GEN_3666; // @[RAM_ST.scala 32:46]
  assign _GEN_3668 = 11'h6cf == RADDR ? 11'h6cf : _GEN_3667; // @[RAM_ST.scala 32:46]
  assign _GEN_3669 = 11'h6d0 == RADDR ? 11'h6d0 : _GEN_3668; // @[RAM_ST.scala 32:46]
  assign _GEN_3670 = 11'h6d1 == RADDR ? 11'h6d1 : _GEN_3669; // @[RAM_ST.scala 32:46]
  assign _GEN_3671 = 11'h6d2 == RADDR ? 11'h6d2 : _GEN_3670; // @[RAM_ST.scala 32:46]
  assign _GEN_3672 = 11'h6d3 == RADDR ? 11'h6d3 : _GEN_3671; // @[RAM_ST.scala 32:46]
  assign _GEN_3673 = 11'h6d4 == RADDR ? 11'h6d4 : _GEN_3672; // @[RAM_ST.scala 32:46]
  assign _GEN_3674 = 11'h6d5 == RADDR ? 11'h6d5 : _GEN_3673; // @[RAM_ST.scala 32:46]
  assign _GEN_3675 = 11'h6d6 == RADDR ? 11'h6d6 : _GEN_3674; // @[RAM_ST.scala 32:46]
  assign _GEN_3676 = 11'h6d7 == RADDR ? 11'h6d7 : _GEN_3675; // @[RAM_ST.scala 32:46]
  assign _GEN_3677 = 11'h6d8 == RADDR ? 11'h6d8 : _GEN_3676; // @[RAM_ST.scala 32:46]
  assign _GEN_3678 = 11'h6d9 == RADDR ? 11'h6d9 : _GEN_3677; // @[RAM_ST.scala 32:46]
  assign _GEN_3679 = 11'h6da == RADDR ? 11'h6da : _GEN_3678; // @[RAM_ST.scala 32:46]
  assign _GEN_3680 = 11'h6db == RADDR ? 11'h6db : _GEN_3679; // @[RAM_ST.scala 32:46]
  assign _GEN_3681 = 11'h6dc == RADDR ? 11'h6dc : _GEN_3680; // @[RAM_ST.scala 32:46]
  assign _GEN_3682 = 11'h6dd == RADDR ? 11'h6dd : _GEN_3681; // @[RAM_ST.scala 32:46]
  assign _GEN_3683 = 11'h6de == RADDR ? 11'h6de : _GEN_3682; // @[RAM_ST.scala 32:46]
  assign _GEN_3684 = 11'h6df == RADDR ? 11'h6df : _GEN_3683; // @[RAM_ST.scala 32:46]
  assign _GEN_3685 = 11'h6e0 == RADDR ? 11'h6e0 : _GEN_3684; // @[RAM_ST.scala 32:46]
  assign _GEN_3686 = 11'h6e1 == RADDR ? 11'h6e1 : _GEN_3685; // @[RAM_ST.scala 32:46]
  assign _GEN_3687 = 11'h6e2 == RADDR ? 11'h6e2 : _GEN_3686; // @[RAM_ST.scala 32:46]
  assign _GEN_3688 = 11'h6e3 == RADDR ? 11'h6e3 : _GEN_3687; // @[RAM_ST.scala 32:46]
  assign _GEN_3689 = 11'h6e4 == RADDR ? 11'h6e4 : _GEN_3688; // @[RAM_ST.scala 32:46]
  assign _GEN_3690 = 11'h6e5 == RADDR ? 11'h6e5 : _GEN_3689; // @[RAM_ST.scala 32:46]
  assign _GEN_3691 = 11'h6e6 == RADDR ? 11'h6e6 : _GEN_3690; // @[RAM_ST.scala 32:46]
  assign _GEN_3692 = 11'h6e7 == RADDR ? 11'h6e7 : _GEN_3691; // @[RAM_ST.scala 32:46]
  assign _GEN_3693 = 11'h6e8 == RADDR ? 11'h6e8 : _GEN_3692; // @[RAM_ST.scala 32:46]
  assign _GEN_3694 = 11'h6e9 == RADDR ? 11'h6e9 : _GEN_3693; // @[RAM_ST.scala 32:46]
  assign _GEN_3695 = 11'h6ea == RADDR ? 11'h6ea : _GEN_3694; // @[RAM_ST.scala 32:46]
  assign _GEN_3696 = 11'h6eb == RADDR ? 11'h6eb : _GEN_3695; // @[RAM_ST.scala 32:46]
  assign _GEN_3697 = 11'h6ec == RADDR ? 11'h6ec : _GEN_3696; // @[RAM_ST.scala 32:46]
  assign _GEN_3698 = 11'h6ed == RADDR ? 11'h6ed : _GEN_3697; // @[RAM_ST.scala 32:46]
  assign _GEN_3699 = 11'h6ee == RADDR ? 11'h6ee : _GEN_3698; // @[RAM_ST.scala 32:46]
  assign _GEN_3700 = 11'h6ef == RADDR ? 11'h6ef : _GEN_3699; // @[RAM_ST.scala 32:46]
  assign _GEN_3701 = 11'h6f0 == RADDR ? 11'h6f0 : _GEN_3700; // @[RAM_ST.scala 32:46]
  assign _GEN_3702 = 11'h6f1 == RADDR ? 11'h6f1 : _GEN_3701; // @[RAM_ST.scala 32:46]
  assign _GEN_3703 = 11'h6f2 == RADDR ? 11'h6f2 : _GEN_3702; // @[RAM_ST.scala 32:46]
  assign _GEN_3704 = 11'h6f3 == RADDR ? 11'h6f3 : _GEN_3703; // @[RAM_ST.scala 32:46]
  assign _GEN_3705 = 11'h6f4 == RADDR ? 11'h6f4 : _GEN_3704; // @[RAM_ST.scala 32:46]
  assign _GEN_3706 = 11'h6f5 == RADDR ? 11'h6f5 : _GEN_3705; // @[RAM_ST.scala 32:46]
  assign _GEN_3707 = 11'h6f6 == RADDR ? 11'h6f6 : _GEN_3706; // @[RAM_ST.scala 32:46]
  assign _GEN_3708 = 11'h6f7 == RADDR ? 11'h6f7 : _GEN_3707; // @[RAM_ST.scala 32:46]
  assign _GEN_3709 = 11'h6f8 == RADDR ? 11'h6f8 : _GEN_3708; // @[RAM_ST.scala 32:46]
  assign _GEN_3710 = 11'h6f9 == RADDR ? 11'h6f9 : _GEN_3709; // @[RAM_ST.scala 32:46]
  assign _GEN_3711 = 11'h6fa == RADDR ? 11'h6fa : _GEN_3710; // @[RAM_ST.scala 32:46]
  assign _GEN_3712 = 11'h6fb == RADDR ? 11'h6fb : _GEN_3711; // @[RAM_ST.scala 32:46]
  assign _GEN_3713 = 11'h6fc == RADDR ? 11'h6fc : _GEN_3712; // @[RAM_ST.scala 32:46]
  assign _GEN_3714 = 11'h6fd == RADDR ? 11'h6fd : _GEN_3713; // @[RAM_ST.scala 32:46]
  assign _GEN_3715 = 11'h6fe == RADDR ? 11'h6fe : _GEN_3714; // @[RAM_ST.scala 32:46]
  assign _GEN_3716 = 11'h6ff == RADDR ? 11'h6ff : _GEN_3715; // @[RAM_ST.scala 32:46]
  assign _GEN_3717 = 11'h700 == RADDR ? 11'h700 : _GEN_3716; // @[RAM_ST.scala 32:46]
  assign _GEN_3718 = 11'h701 == RADDR ? 11'h701 : _GEN_3717; // @[RAM_ST.scala 32:46]
  assign _GEN_3719 = 11'h702 == RADDR ? 11'h702 : _GEN_3718; // @[RAM_ST.scala 32:46]
  assign _GEN_3720 = 11'h703 == RADDR ? 11'h703 : _GEN_3719; // @[RAM_ST.scala 32:46]
  assign _GEN_3721 = 11'h704 == RADDR ? 11'h704 : _GEN_3720; // @[RAM_ST.scala 32:46]
  assign _GEN_3722 = 11'h705 == RADDR ? 11'h705 : _GEN_3721; // @[RAM_ST.scala 32:46]
  assign _GEN_3723 = 11'h706 == RADDR ? 11'h706 : _GEN_3722; // @[RAM_ST.scala 32:46]
  assign _GEN_3724 = 11'h707 == RADDR ? 11'h707 : _GEN_3723; // @[RAM_ST.scala 32:46]
  assign _GEN_3725 = 11'h708 == RADDR ? 11'h708 : _GEN_3724; // @[RAM_ST.scala 32:46]
  assign _GEN_3726 = 11'h709 == RADDR ? 11'h709 : _GEN_3725; // @[RAM_ST.scala 32:46]
  assign _GEN_3727 = 11'h70a == RADDR ? 11'h70a : _GEN_3726; // @[RAM_ST.scala 32:46]
  assign _GEN_3728 = 11'h70b == RADDR ? 11'h70b : _GEN_3727; // @[RAM_ST.scala 32:46]
  assign _GEN_3729 = 11'h70c == RADDR ? 11'h70c : _GEN_3728; // @[RAM_ST.scala 32:46]
  assign _GEN_3730 = 11'h70d == RADDR ? 11'h70d : _GEN_3729; // @[RAM_ST.scala 32:46]
  assign _GEN_3731 = 11'h70e == RADDR ? 11'h70e : _GEN_3730; // @[RAM_ST.scala 32:46]
  assign _GEN_3732 = 11'h70f == RADDR ? 11'h70f : _GEN_3731; // @[RAM_ST.scala 32:46]
  assign _GEN_3733 = 11'h710 == RADDR ? 11'h710 : _GEN_3732; // @[RAM_ST.scala 32:46]
  assign _GEN_3734 = 11'h711 == RADDR ? 11'h711 : _GEN_3733; // @[RAM_ST.scala 32:46]
  assign _GEN_3735 = 11'h712 == RADDR ? 11'h712 : _GEN_3734; // @[RAM_ST.scala 32:46]
  assign _GEN_3736 = 11'h713 == RADDR ? 11'h713 : _GEN_3735; // @[RAM_ST.scala 32:46]
  assign _GEN_3737 = 11'h714 == RADDR ? 11'h714 : _GEN_3736; // @[RAM_ST.scala 32:46]
  assign _GEN_3738 = 11'h715 == RADDR ? 11'h715 : _GEN_3737; // @[RAM_ST.scala 32:46]
  assign _GEN_3739 = 11'h716 == RADDR ? 11'h716 : _GEN_3738; // @[RAM_ST.scala 32:46]
  assign _GEN_3740 = 11'h717 == RADDR ? 11'h717 : _GEN_3739; // @[RAM_ST.scala 32:46]
  assign _GEN_3741 = 11'h718 == RADDR ? 11'h718 : _GEN_3740; // @[RAM_ST.scala 32:46]
  assign _GEN_3742 = 11'h719 == RADDR ? 11'h719 : _GEN_3741; // @[RAM_ST.scala 32:46]
  assign _GEN_3743 = 11'h71a == RADDR ? 11'h71a : _GEN_3742; // @[RAM_ST.scala 32:46]
  assign _GEN_3744 = 11'h71b == RADDR ? 11'h71b : _GEN_3743; // @[RAM_ST.scala 32:46]
  assign _GEN_3745 = 11'h71c == RADDR ? 11'h71c : _GEN_3744; // @[RAM_ST.scala 32:46]
  assign _GEN_3746 = 11'h71d == RADDR ? 11'h71d : _GEN_3745; // @[RAM_ST.scala 32:46]
  assign _GEN_3747 = 11'h71e == RADDR ? 11'h71e : _GEN_3746; // @[RAM_ST.scala 32:46]
  assign _GEN_3748 = 11'h71f == RADDR ? 11'h71f : _GEN_3747; // @[RAM_ST.scala 32:46]
  assign _GEN_3749 = 11'h720 == RADDR ? 11'h720 : _GEN_3748; // @[RAM_ST.scala 32:46]
  assign _GEN_3750 = 11'h721 == RADDR ? 11'h721 : _GEN_3749; // @[RAM_ST.scala 32:46]
  assign _GEN_3751 = 11'h722 == RADDR ? 11'h722 : _GEN_3750; // @[RAM_ST.scala 32:46]
  assign _GEN_3752 = 11'h723 == RADDR ? 11'h723 : _GEN_3751; // @[RAM_ST.scala 32:46]
  assign _GEN_3753 = 11'h724 == RADDR ? 11'h724 : _GEN_3752; // @[RAM_ST.scala 32:46]
  assign _GEN_3754 = 11'h725 == RADDR ? 11'h725 : _GEN_3753; // @[RAM_ST.scala 32:46]
  assign _GEN_3755 = 11'h726 == RADDR ? 11'h726 : _GEN_3754; // @[RAM_ST.scala 32:46]
  assign _GEN_3756 = 11'h727 == RADDR ? 11'h727 : _GEN_3755; // @[RAM_ST.scala 32:46]
  assign _GEN_3757 = 11'h728 == RADDR ? 11'h728 : _GEN_3756; // @[RAM_ST.scala 32:46]
  assign _GEN_3758 = 11'h729 == RADDR ? 11'h729 : _GEN_3757; // @[RAM_ST.scala 32:46]
  assign _GEN_3759 = 11'h72a == RADDR ? 11'h72a : _GEN_3758; // @[RAM_ST.scala 32:46]
  assign _GEN_3760 = 11'h72b == RADDR ? 11'h72b : _GEN_3759; // @[RAM_ST.scala 32:46]
  assign _GEN_3761 = 11'h72c == RADDR ? 11'h72c : _GEN_3760; // @[RAM_ST.scala 32:46]
  assign _GEN_3762 = 11'h72d == RADDR ? 11'h72d : _GEN_3761; // @[RAM_ST.scala 32:46]
  assign _GEN_3763 = 11'h72e == RADDR ? 11'h72e : _GEN_3762; // @[RAM_ST.scala 32:46]
  assign _GEN_3764 = 11'h72f == RADDR ? 11'h72f : _GEN_3763; // @[RAM_ST.scala 32:46]
  assign _GEN_3765 = 11'h730 == RADDR ? 11'h730 : _GEN_3764; // @[RAM_ST.scala 32:46]
  assign _GEN_3766 = 11'h731 == RADDR ? 11'h731 : _GEN_3765; // @[RAM_ST.scala 32:46]
  assign _GEN_3767 = 11'h732 == RADDR ? 11'h732 : _GEN_3766; // @[RAM_ST.scala 32:46]
  assign _GEN_3768 = 11'h733 == RADDR ? 11'h733 : _GEN_3767; // @[RAM_ST.scala 32:46]
  assign _GEN_3769 = 11'h734 == RADDR ? 11'h734 : _GEN_3768; // @[RAM_ST.scala 32:46]
  assign _GEN_3770 = 11'h735 == RADDR ? 11'h735 : _GEN_3769; // @[RAM_ST.scala 32:46]
  assign _GEN_3771 = 11'h736 == RADDR ? 11'h736 : _GEN_3770; // @[RAM_ST.scala 32:46]
  assign _GEN_3772 = 11'h737 == RADDR ? 11'h737 : _GEN_3771; // @[RAM_ST.scala 32:46]
  assign _GEN_3773 = 11'h738 == RADDR ? 11'h738 : _GEN_3772; // @[RAM_ST.scala 32:46]
  assign _GEN_3774 = 11'h739 == RADDR ? 11'h739 : _GEN_3773; // @[RAM_ST.scala 32:46]
  assign _GEN_3775 = 11'h73a == RADDR ? 11'h73a : _GEN_3774; // @[RAM_ST.scala 32:46]
  assign _GEN_3776 = 11'h73b == RADDR ? 11'h73b : _GEN_3775; // @[RAM_ST.scala 32:46]
  assign _GEN_3777 = 11'h73c == RADDR ? 11'h73c : _GEN_3776; // @[RAM_ST.scala 32:46]
  assign _GEN_3778 = 11'h73d == RADDR ? 11'h73d : _GEN_3777; // @[RAM_ST.scala 32:46]
  assign _GEN_3779 = 11'h73e == RADDR ? 11'h73e : _GEN_3778; // @[RAM_ST.scala 32:46]
  assign _GEN_3780 = 11'h73f == RADDR ? 11'h73f : _GEN_3779; // @[RAM_ST.scala 32:46]
  assign _GEN_3781 = 11'h740 == RADDR ? 11'h740 : _GEN_3780; // @[RAM_ST.scala 32:46]
  assign _GEN_3782 = 11'h741 == RADDR ? 11'h741 : _GEN_3781; // @[RAM_ST.scala 32:46]
  assign _GEN_3783 = 11'h742 == RADDR ? 11'h742 : _GEN_3782; // @[RAM_ST.scala 32:46]
  assign _GEN_3784 = 11'h743 == RADDR ? 11'h743 : _GEN_3783; // @[RAM_ST.scala 32:46]
  assign _GEN_3785 = 11'h744 == RADDR ? 11'h744 : _GEN_3784; // @[RAM_ST.scala 32:46]
  assign _GEN_3786 = 11'h745 == RADDR ? 11'h745 : _GEN_3785; // @[RAM_ST.scala 32:46]
  assign _GEN_3787 = 11'h746 == RADDR ? 11'h746 : _GEN_3786; // @[RAM_ST.scala 32:46]
  assign _GEN_3788 = 11'h747 == RADDR ? 11'h747 : _GEN_3787; // @[RAM_ST.scala 32:46]
  assign _GEN_3789 = 11'h748 == RADDR ? 11'h748 : _GEN_3788; // @[RAM_ST.scala 32:46]
  assign _GEN_3790 = 11'h749 == RADDR ? 11'h749 : _GEN_3789; // @[RAM_ST.scala 32:46]
  assign _GEN_3791 = 11'h74a == RADDR ? 11'h74a : _GEN_3790; // @[RAM_ST.scala 32:46]
  assign _GEN_3792 = 11'h74b == RADDR ? 11'h74b : _GEN_3791; // @[RAM_ST.scala 32:46]
  assign _GEN_3793 = 11'h74c == RADDR ? 11'h74c : _GEN_3792; // @[RAM_ST.scala 32:46]
  assign _GEN_3794 = 11'h74d == RADDR ? 11'h74d : _GEN_3793; // @[RAM_ST.scala 32:46]
  assign _GEN_3795 = 11'h74e == RADDR ? 11'h74e : _GEN_3794; // @[RAM_ST.scala 32:46]
  assign _GEN_3796 = 11'h74f == RADDR ? 11'h74f : _GEN_3795; // @[RAM_ST.scala 32:46]
  assign _GEN_3797 = 11'h750 == RADDR ? 11'h750 : _GEN_3796; // @[RAM_ST.scala 32:46]
  assign _GEN_3798 = 11'h751 == RADDR ? 11'h751 : _GEN_3797; // @[RAM_ST.scala 32:46]
  assign _GEN_3799 = 11'h752 == RADDR ? 11'h752 : _GEN_3798; // @[RAM_ST.scala 32:46]
  assign _GEN_3800 = 11'h753 == RADDR ? 11'h753 : _GEN_3799; // @[RAM_ST.scala 32:46]
  assign _GEN_3801 = 11'h754 == RADDR ? 11'h754 : _GEN_3800; // @[RAM_ST.scala 32:46]
  assign _GEN_3802 = 11'h755 == RADDR ? 11'h755 : _GEN_3801; // @[RAM_ST.scala 32:46]
  assign _GEN_3803 = 11'h756 == RADDR ? 11'h756 : _GEN_3802; // @[RAM_ST.scala 32:46]
  assign _GEN_3804 = 11'h757 == RADDR ? 11'h757 : _GEN_3803; // @[RAM_ST.scala 32:46]
  assign _GEN_3805 = 11'h758 == RADDR ? 11'h758 : _GEN_3804; // @[RAM_ST.scala 32:46]
  assign _GEN_3806 = 11'h759 == RADDR ? 11'h759 : _GEN_3805; // @[RAM_ST.scala 32:46]
  assign _GEN_3807 = 11'h75a == RADDR ? 11'h75a : _GEN_3806; // @[RAM_ST.scala 32:46]
  assign _GEN_3808 = 11'h75b == RADDR ? 11'h75b : _GEN_3807; // @[RAM_ST.scala 32:46]
  assign _GEN_3809 = 11'h75c == RADDR ? 11'h75c : _GEN_3808; // @[RAM_ST.scala 32:46]
  assign _GEN_3810 = 11'h75d == RADDR ? 11'h75d : _GEN_3809; // @[RAM_ST.scala 32:46]
  assign _GEN_3811 = 11'h75e == RADDR ? 11'h75e : _GEN_3810; // @[RAM_ST.scala 32:46]
  assign _GEN_3812 = 11'h75f == RADDR ? 11'h75f : _GEN_3811; // @[RAM_ST.scala 32:46]
  assign _GEN_3813 = 11'h760 == RADDR ? 11'h760 : _GEN_3812; // @[RAM_ST.scala 32:46]
  assign _GEN_3814 = 11'h761 == RADDR ? 11'h761 : _GEN_3813; // @[RAM_ST.scala 32:46]
  assign _GEN_3815 = 11'h762 == RADDR ? 11'h762 : _GEN_3814; // @[RAM_ST.scala 32:46]
  assign _GEN_3816 = 11'h763 == RADDR ? 11'h763 : _GEN_3815; // @[RAM_ST.scala 32:46]
  assign _GEN_3817 = 11'h764 == RADDR ? 11'h764 : _GEN_3816; // @[RAM_ST.scala 32:46]
  assign _GEN_3818 = 11'h765 == RADDR ? 11'h765 : _GEN_3817; // @[RAM_ST.scala 32:46]
  assign _GEN_3819 = 11'h766 == RADDR ? 11'h766 : _GEN_3818; // @[RAM_ST.scala 32:46]
  assign _GEN_3820 = 11'h767 == RADDR ? 11'h767 : _GEN_3819; // @[RAM_ST.scala 32:46]
  assign _GEN_3821 = 11'h768 == RADDR ? 11'h768 : _GEN_3820; // @[RAM_ST.scala 32:46]
  assign _GEN_3822 = 11'h769 == RADDR ? 11'h769 : _GEN_3821; // @[RAM_ST.scala 32:46]
  assign _GEN_3823 = 11'h76a == RADDR ? 11'h76a : _GEN_3822; // @[RAM_ST.scala 32:46]
  assign _GEN_3824 = 11'h76b == RADDR ? 11'h76b : _GEN_3823; // @[RAM_ST.scala 32:46]
  assign _GEN_3825 = 11'h76c == RADDR ? 11'h76c : _GEN_3824; // @[RAM_ST.scala 32:46]
  assign _GEN_3826 = 11'h76d == RADDR ? 11'h76d : _GEN_3825; // @[RAM_ST.scala 32:46]
  assign _GEN_3827 = 11'h76e == RADDR ? 11'h76e : _GEN_3826; // @[RAM_ST.scala 32:46]
  assign _GEN_3828 = 11'h76f == RADDR ? 11'h76f : _GEN_3827; // @[RAM_ST.scala 32:46]
  assign _GEN_3829 = 11'h770 == RADDR ? 11'h770 : _GEN_3828; // @[RAM_ST.scala 32:46]
  assign _GEN_3830 = 11'h771 == RADDR ? 11'h771 : _GEN_3829; // @[RAM_ST.scala 32:46]
  assign _GEN_3831 = 11'h772 == RADDR ? 11'h772 : _GEN_3830; // @[RAM_ST.scala 32:46]
  assign _GEN_3832 = 11'h773 == RADDR ? 11'h773 : _GEN_3831; // @[RAM_ST.scala 32:46]
  assign _GEN_3833 = 11'h774 == RADDR ? 11'h774 : _GEN_3832; // @[RAM_ST.scala 32:46]
  assign _GEN_3834 = 11'h775 == RADDR ? 11'h775 : _GEN_3833; // @[RAM_ST.scala 32:46]
  assign _GEN_3835 = 11'h776 == RADDR ? 11'h776 : _GEN_3834; // @[RAM_ST.scala 32:46]
  assign _GEN_3836 = 11'h777 == RADDR ? 11'h777 : _GEN_3835; // @[RAM_ST.scala 32:46]
  assign _GEN_3837 = 11'h778 == RADDR ? 11'h778 : _GEN_3836; // @[RAM_ST.scala 32:46]
  assign _GEN_3838 = 11'h779 == RADDR ? 11'h779 : _GEN_3837; // @[RAM_ST.scala 32:46]
  assign _GEN_3839 = 11'h77a == RADDR ? 11'h77a : _GEN_3838; // @[RAM_ST.scala 32:46]
  assign _GEN_3840 = 11'h77b == RADDR ? 11'h77b : _GEN_3839; // @[RAM_ST.scala 32:46]
  assign _GEN_3841 = 11'h77c == RADDR ? 11'h77c : _GEN_3840; // @[RAM_ST.scala 32:46]
  assign _GEN_3842 = 11'h77d == RADDR ? 11'h77d : _GEN_3841; // @[RAM_ST.scala 32:46]
  assign _GEN_3843 = 11'h77e == RADDR ? 11'h77e : _GEN_3842; // @[RAM_ST.scala 32:46]
  assign _GEN_3844 = 11'h77f == RADDR ? 11'h77f : _GEN_3843; // @[RAM_ST.scala 32:46]
  assign _T_3 = {{1'd0}, _GEN_3844}; // @[RAM_ST.scala 32:46]
  assign RDATA = ram__T_8_data; // @[RAM_ST.scala 32:9]
  assign write_elem_counter_CE = WE; // @[RAM_ST.scala 23:25]
  assign read_elem_counter_CE = RE; // @[RAM_ST.scala 24:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1920; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram__T_8_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ram__T_8_addr_pipe_0 = _RAND_3[10:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_2_en & ram__T_2_mask) begin
      ram[ram__T_2_addr] <= ram__T_2_data; // @[RAM_ST.scala 29:24]
    end
    ram__T_8_en_pipe_0 <= read_elem_counter_valid;
    if (read_elem_counter_valid) begin
      ram__T_8_addr_pipe_0 <= _T_3[10:0];
    end
  end
endmodule
module NestedCounters_4(
  input   clock,
  input   reset,
  input   CE,
  output  valid
);
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[Counter.scala 37:24]
  wire [1:0] _T_3; // @[Counter.scala 38:22]
  assign _T_1 = value == 2'h2; // @[Counter.scala 37:24]
  assign _T_3 = value + 2'h1; // @[Counter.scala 38:22]
  assign valid = value < 2'h1; // @[NestedCounters.scala 48:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 2'h0;
    end else if (CE) begin
      if (_T_1) begin
        value <= 2'h0;
      end else begin
        value <= _T_3;
      end
    end
  end
endmodule
module ShiftTN(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I,
  output [7:0] O
);
  wire  value_store_clock; // @[ShiftTN.scala 42:27]
  wire  value_store_RE; // @[ShiftTN.scala 42:27]
  wire [10:0] value_store_RADDR; // @[ShiftTN.scala 42:27]
  wire [7:0] value_store_RDATA; // @[ShiftTN.scala 42:27]
  wire  value_store_WE; // @[ShiftTN.scala 42:27]
  wire [10:0] value_store_WADDR; // @[ShiftTN.scala 42:27]
  wire [7:0] value_store_WDATA; // @[ShiftTN.scala 42:27]
  wire  next_ram_addr_CE; // @[ShiftTN.scala 44:29]
  wire  next_ram_addr_valid; // @[ShiftTN.scala 44:29]
  wire  inner_valid_clock; // @[ShiftTN.scala 56:27]
  wire  inner_valid_reset; // @[ShiftTN.scala 56:27]
  wire  inner_valid_CE; // @[ShiftTN.scala 56:27]
  wire  inner_valid_valid; // @[ShiftTN.scala 56:27]
  wire  _T_2; // @[ShiftTN.scala 58:74]
  reg [10:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_3; // @[Counter.scala 37:24]
  wire [10:0] _T_5; // @[Counter.scala 38:22]
  RAM_ST value_store ( // @[ShiftTN.scala 42:27]
    .clock(value_store_clock),
    .RE(value_store_RE),
    .RADDR(value_store_RADDR),
    .RDATA(value_store_RDATA),
    .WE(value_store_WE),
    .WADDR(value_store_WADDR),
    .WDATA(value_store_WDATA)
  );
  NestedCounters next_ram_addr ( // @[ShiftTN.scala 44:29]
    .CE(next_ram_addr_CE),
    .valid(next_ram_addr_valid)
  );
  NestedCounters_4 inner_valid ( // @[ShiftTN.scala 56:27]
    .clock(inner_valid_clock),
    .reset(inner_valid_reset),
    .CE(inner_valid_CE),
    .valid(inner_valid_valid)
  );
  assign _T_2 = valid_up & inner_valid_valid; // @[ShiftTN.scala 58:74]
  assign _T_3 = value == 11'h77f; // @[Counter.scala 37:24]
  assign _T_5 = value + 11'h1; // @[Counter.scala 38:22]
  assign valid_down = valid_up; // @[ShiftTN.scala 69:14]
  assign O = value_store_RDATA; // @[ShiftTN.scala 66:5]
  assign value_store_clock = clock;
  assign value_store_RE = valid_up & inner_valid_valid; // @[ShiftTN.scala 64:18]
  assign value_store_RADDR = _T_3 ? 11'h0 : _T_5; // @[ShiftTN.scala 61:74 ShiftTN.scala 62:36]
  assign value_store_WE = valid_up & inner_valid_valid; // @[ShiftTN.scala 63:18]
  assign value_store_WADDR = value; // @[ShiftTN.scala 60:21]
  assign value_store_WDATA = I; // @[ShiftTN.scala 65:21]
  assign next_ram_addr_CE = valid_up; // @[ShiftTN.scala 45:20]
  assign inner_valid_clock = clock;
  assign inner_valid_reset = reset;
  assign inner_valid_CE = valid_up; // @[ShiftTN.scala 57:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[10:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 11'h0;
    end else if (_T_2) begin
      if (_T_3) begin
        value <= 11'h0;
      end else begin
        value <= _T_5;
      end
    end
  end
endmodule
module RAM_ST_2(
  input        clock,
  input        RE,
  output [7:0] RDATA,
  input        WE,
  input  [7:0] WDATA
);
  wire  write_elem_counter_CE; // @[RAM_ST.scala 20:34]
  wire  write_elem_counter_valid; // @[RAM_ST.scala 20:34]
  wire  read_elem_counter_CE; // @[RAM_ST.scala 21:33]
  wire  read_elem_counter_valid; // @[RAM_ST.scala 21:33]
  reg [7:0] ram [0:0]; // @[RAM_ST.scala 29:24]
  reg [31:0] _RAND_0;
  wire [7:0] ram__T_6_data; // @[RAM_ST.scala 29:24]
  wire  ram__T_6_addr; // @[RAM_ST.scala 29:24]
  wire [7:0] ram__T_2_data; // @[RAM_ST.scala 29:24]
  wire  ram__T_2_addr; // @[RAM_ST.scala 29:24]
  wire  ram__T_2_mask; // @[RAM_ST.scala 29:24]
  wire  ram__T_2_en; // @[RAM_ST.scala 29:24]
  reg  ram__T_6_en_pipe_0;
  reg [31:0] _RAND_1;
  reg  ram__T_6_addr_pipe_0;
  reg [31:0] _RAND_2;
  NestedCountersWithNumValid write_elem_counter ( // @[RAM_ST.scala 20:34]
    .CE(write_elem_counter_CE),
    .valid(write_elem_counter_valid)
  );
  NestedCountersWithNumValid read_elem_counter ( // @[RAM_ST.scala 21:33]
    .CE(read_elem_counter_CE),
    .valid(read_elem_counter_valid)
  );
  assign ram__T_6_addr = ram__T_6_addr_pipe_0;
  assign ram__T_6_data = ram[ram__T_6_addr]; // @[RAM_ST.scala 29:24]
  assign ram__T_2_data = WDATA;
  assign ram__T_2_addr = 1'h0;
  assign ram__T_2_mask = 1'h1;
  assign ram__T_2_en = write_elem_counter_valid;
  assign RDATA = ram__T_6_data; // @[RAM_ST.scala 32:9]
  assign write_elem_counter_CE = WE; // @[RAM_ST.scala 23:25]
  assign read_elem_counter_CE = RE; // @[RAM_ST.scala 24:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram__T_6_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram__T_6_addr_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_2_en & ram__T_2_mask) begin
      ram[ram__T_2_addr] <= ram__T_2_data; // @[RAM_ST.scala 29:24]
    end
    ram__T_6_en_pipe_0 <= read_elem_counter_valid;
    if (read_elem_counter_valid) begin
      ram__T_6_addr_pipe_0 <= 1'h0;
    end
  end
endmodule
module ShiftTN_2(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I,
  output [7:0] O
);
  wire  value_store_clock; // @[ShiftTN.scala 42:27]
  wire  value_store_RE; // @[ShiftTN.scala 42:27]
  wire [7:0] value_store_RDATA; // @[ShiftTN.scala 42:27]
  wire  value_store_WE; // @[ShiftTN.scala 42:27]
  wire [7:0] value_store_WDATA; // @[ShiftTN.scala 42:27]
  wire  next_ram_addr_CE; // @[ShiftTN.scala 44:29]
  wire  next_ram_addr_valid; // @[ShiftTN.scala 44:29]
  wire  inner_valid_clock; // @[ShiftTN.scala 56:27]
  wire  inner_valid_reset; // @[ShiftTN.scala 56:27]
  wire  inner_valid_CE; // @[ShiftTN.scala 56:27]
  wire  inner_valid_valid; // @[ShiftTN.scala 56:27]
  RAM_ST_2 value_store ( // @[ShiftTN.scala 42:27]
    .clock(value_store_clock),
    .RE(value_store_RE),
    .RDATA(value_store_RDATA),
    .WE(value_store_WE),
    .WDATA(value_store_WDATA)
  );
  NestedCounters next_ram_addr ( // @[ShiftTN.scala 44:29]
    .CE(next_ram_addr_CE),
    .valid(next_ram_addr_valid)
  );
  NestedCounters_4 inner_valid ( // @[ShiftTN.scala 56:27]
    .clock(inner_valid_clock),
    .reset(inner_valid_reset),
    .CE(inner_valid_CE),
    .valid(inner_valid_valid)
  );
  assign valid_down = valid_up; // @[ShiftTN.scala 69:14]
  assign O = value_store_RDATA; // @[ShiftTN.scala 66:5]
  assign value_store_clock = clock;
  assign value_store_RE = valid_up & inner_valid_valid; // @[ShiftTN.scala 64:18]
  assign value_store_WE = valid_up & inner_valid_valid; // @[ShiftTN.scala 63:18]
  assign value_store_WDATA = I; // @[ShiftTN.scala 65:21]
  assign next_ram_addr_CE = valid_up; // @[ShiftTN.scala 45:20]
  assign inner_valid_clock = clock;
  assign inner_valid_reset = reset;
  assign inner_valid_CE = valid_up; // @[ShiftTN.scala 57:18]
endmodule
module SSeqTupleCreator(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0 = I0; // @[Tuple.scala 12:32]
  assign O_1 = I1; // @[Tuple.scala 13:32]
endmodule
module Map2T(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1; // @[Map2T.scala 8:20]
  SSeqTupleCreator op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0(op_I0),
    .I1(op_I1),
    .O_0(op_O_0),
    .O_1(op_O_1)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0 = op_O_0; // @[Map2T.scala 17:7]
  assign O_1 = op_O_1; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0 = I0; // @[Map2T.scala 15:11]
  assign op_I1 = I1; // @[Map2T.scala 16:11]
endmodule
module Map2T_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1; // @[Map2T.scala 8:20]
  Map2T op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0(op_I0),
    .I1(op_I1),
    .O_0(op_O_0),
    .O_1(op_O_1)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0 = op_O_0; // @[Map2T.scala 17:7]
  assign O_1 = op_O_1; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0 = I0; // @[Map2T.scala 15:11]
  assign op_I1 = I1; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0 = I0_0; // @[Tuple.scala 24:34]
  assign O_1 = I0_1; // @[Tuple.scala 24:34]
  assign O_2 = I1; // @[Tuple.scala 26:32]
endmodule
module Map2T_2(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2; // @[Map2T.scala 8:20]
  SSeqTupleAppender op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I1(op_I1),
    .O_0(op_O_0),
    .O_1(op_O_1),
    .O_2(op_O_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0 = op_O_0; // @[Map2T.scala 17:7]
  assign O_1 = op_O_1; // @[Map2T.scala 17:7]
  assign O_2 = op_O_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I1 = I1; // @[Map2T.scala 16:11]
endmodule
module Map2T_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2; // @[Map2T.scala 8:20]
  Map2T_2 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I1(op_I1),
    .O_0(op_O_0),
    .O_1(op_O_1),
    .O_2(op_O_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0 = op_O_0; // @[Map2T.scala 17:7]
  assign O_1 = op_O_1; // @[Map2T.scala 17:7]
  assign O_2 = op_O_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I1 = I1; // @[Map2T.scala 16:11]
endmodule
module Passthrough(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0 = I_0; // @[Passthrough.scala 17:68]
  assign O_0_1 = I_1; // @[Passthrough.scala 17:68]
  assign O_0_2 = I_2; // @[Passthrough.scala 17:68]
endmodule
module Serialize(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O
);
  wire  elem_counter_CE; // @[Serialize.scala 14:28]
  wire  elem_counter_valid; // @[Serialize.scala 14:28]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[Counter.scala 37:24]
  wire [1:0] _T_3; // @[Counter.scala 38:22]
  reg [7:0] mux_input_wire_1; // @[Serialize.scala 39:47]
  reg [31:0] _RAND_1;
  reg [7:0] mux_input_wire_2; // @[Serialize.scala 39:47]
  reg [31:0] _RAND_2;
  wire  _T_7; // @[Serialize.scala 42:34]
  wire  _T_8; // @[Serialize.scala 42:42]
  wire  _T_11; // @[Mux.scala 68:19]
  wire  _T_13; // @[Mux.scala 68:19]
  wire  _T_15; // @[Mux.scala 68:19]
  reg [7:0] _T_17; // @[Serialize.scala 53:15]
  reg [31:0] _RAND_3;
  reg  _T_18; // @[Serialize.scala 54:24]
  reg [31:0] _RAND_4;
  NestedCountersWithNumValid elem_counter ( // @[Serialize.scala 14:28]
    .CE(elem_counter_CE),
    .valid(elem_counter_valid)
  );
  assign _T_1 = value == 2'h2; // @[Counter.scala 37:24]
  assign _T_3 = value + 2'h1; // @[Counter.scala 38:22]
  assign _T_7 = value == 2'h0; // @[Serialize.scala 42:34]
  assign _T_8 = _T_7 & valid_up; // @[Serialize.scala 42:42]
  assign _T_11 = 2'h2 == value; // @[Mux.scala 68:19]
  assign _T_13 = 2'h1 == value; // @[Mux.scala 68:19]
  assign _T_15 = 2'h0 == value; // @[Mux.scala 68:19]
  assign valid_down = _T_18; // @[Serialize.scala 54:14]
  assign O = _T_17; // @[Serialize.scala 53:5]
  assign elem_counter_CE = valid_up; // @[Serialize.scala 16:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mux_input_wire_1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mux_input_wire_2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_17 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_18 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 2'h0;
    end else if (valid_up) begin
      if (_T_1) begin
        value <= 2'h0;
      end else begin
        value <= _T_3;
      end
    end
    if (_T_8) begin
      mux_input_wire_1 <= I_1;
    end
    if (_T_8) begin
      mux_input_wire_2 <= I_2;
    end
    if (_T_15) begin
      _T_17 <= I_0;
    end else if (_T_13) begin
      _T_17 <= mux_input_wire_1;
    end else if (_T_11) begin
      _T_17 <= mux_input_wire_2;
    end else begin
      _T_17 <= I_0;
    end
    if (reset) begin
      _T_18 <= 1'h0;
    end else begin
      _T_18 <= valid_up;
    end
  end
endmodule
module MapS(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  output [7:0] O_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  Serialize fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
endmodule
module MapT(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  output [7:0] O_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0; // @[MapT.scala 8:20]
  MapS op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0(op_I_0_0),
    .I_0_1(op_I_0_1),
    .I_0_2(op_I_0_2),
    .O_0(op_O_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0 = I_0_0; // @[MapT.scala 14:10]
  assign op_I_0_1 = I_0_1; // @[MapT.scala 14:10]
  assign op_I_0_2 = I_0_2; // @[MapT.scala 14:10]
endmodule
module Map2S(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I1_0,
  output [7:0] O_0_0,
  output [7:0] O_0_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1; // @[Map2S.scala 9:22]
  SSeqTupleCreator fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2T_8(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I1_0,
  output [7:0] O_0_0,
  output [7:0] O_0_1
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1; // @[Map2T.scala 8:20]
  Map2S op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I1_0(op_I1_0),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
endmodule
module Map2S_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I1_0,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2; // @[Map2S.scala 9:22]
  SSeqTupleAppender fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_0_2 = fst_op_O_2; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2T_13(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I1_0,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_2; // @[Map2T.scala 8:20]
  Map2S_1 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I1_0(op_I1_0),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_0_2(op_O_0_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign O_0_2 = op_O_0_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
endmodule
module Passthrough_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0 = I_0_0; // @[Passthrough.scala 17:68]
  assign O_0_1 = I_0_1; // @[Passthrough.scala 17:68]
  assign O_0_2 = I_0_2; // @[Passthrough.scala 17:68]
endmodule
module Passthrough_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0 = I_0_0; // @[Passthrough.scala 17:68]
  assign O_1 = I_0_1; // @[Passthrough.scala 17:68]
  assign O_2 = I_0_2; // @[Passthrough.scala 17:68]
endmodule
module MapT_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2; // @[MapT.scala 8:20]
  Passthrough_4 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0(op_I_0_0),
    .I_0_1(op_I_0_1),
    .I_0_2(op_I_0_2),
    .O_0(op_O_0),
    .O_1(op_O_1),
    .O_2(op_O_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign O_1 = op_O_1; // @[MapT.scala 15:7]
  assign O_2 = op_O_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0 = I_0_0; // @[MapT.scala 14:10]
  assign op_I_0_1 = I_0_1; // @[MapT.scala 14:10]
  assign op_I_0_2 = I_0_2; // @[MapT.scala 14:10]
endmodule
module InitialDelayCounter(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [1:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [1:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 2'h2; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 2'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 2'h2; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 2'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module AtomTuple(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_t0b,
  output [7:0] O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Map2T_14(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_t0b,
  output [7:0] O_t1b
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_t0b; // @[Map2T.scala 8:20]
  wire [7:0] op_O_t1b; // @[Map2T.scala 8:20]
  AtomTuple op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0(op_I0),
    .I1(op_I1),
    .O_t0b(op_O_t0b),
    .O_t1b(op_O_t1b)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_t0b = op_O_t0b; // @[Map2T.scala 17:7]
  assign O_t1b = op_O_t1b; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0 = I0; // @[Map2T.scala 15:11]
  assign op_I1 = I1; // @[Map2T.scala 16:11]
endmodule
module Map2S_2(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_t0b,
  output [7:0] O_0_t1b,
  output [7:0] O_1_t0b,
  output [7:0] O_1_t1b,
  output [7:0] O_2_t0b,
  output [7:0] O_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  Map2T_14 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  Map2T_14 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  Map2T_14 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_t0b(other_ops_1_O_t0b),
    .O_t1b(other_ops_1_O_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign O_2_t0b = other_ops_1_O_t0b; // @[Map2S.scala 24:12]
  assign O_2_t1b = other_ops_1_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_15(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_t0b,
  output [7:0] O_0_t1b,
  output [7:0] O_1_t0b,
  output [7:0] O_1_t1b,
  output [7:0] O_2_t0b,
  output [7:0] O_2_t1b
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_t0b; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_t1b; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_t0b; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_t1b; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_t0b; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_t1b; // @[Map2T.scala 8:20]
  Map2S_2 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I0_2(op_I0_2),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .O_0_t0b(op_O_0_t0b),
    .O_0_t1b(op_O_0_t1b),
    .O_1_t0b(op_O_1_t0b),
    .O_1_t1b(op_O_1_t1b),
    .O_2_t0b(op_O_2_t0b),
    .O_2_t1b(op_O_2_t1b)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_t0b = op_O_0_t0b; // @[Map2T.scala 17:7]
  assign O_0_t1b = op_O_0_t1b; // @[Map2T.scala 17:7]
  assign O_1_t0b = op_O_1_t0b; // @[Map2T.scala 17:7]
  assign O_1_t1b = op_O_1_t1b; // @[Map2T.scala 17:7]
  assign O_2_t0b = op_O_2_t0b; // @[Map2T.scala 17:7]
  assign O_2_t1b = op_O_2_t1b; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I0_2 = I0_2; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
endmodule
module LShift(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  wire [262:0] _GEN_0; // @[Arithmetic.scala 301:25]
  wire [262:0] _T; // @[Arithmetic.scala 301:25]
  assign _GEN_0 = {{255'd0}, I_t0b}; // @[Arithmetic.scala 301:25]
  assign _T = _GEN_0 << I_t1b; // @[Arithmetic.scala 301:25]
  assign valid_down = valid_up; // @[Arithmetic.scala 303:14]
  assign O = _T[7:0]; // @[Arithmetic.scala 301:7]
endmodule
module MapT_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_t0b; // @[MapT.scala 8:20]
  wire [7:0] op_I_t1b; // @[MapT.scala 8:20]
  wire [7:0] op_O; // @[MapT.scala 8:20]
  LShift op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_t0b(op_I_t0b),
    .I_t1b(op_I_t1b),
    .O(op_O)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O = op_O; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_t0b = I_t0b; // @[MapT.scala 14:10]
  assign op_I_t1b = I_t1b; // @[MapT.scala 14:10]
endmodule
module MapS_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  input  [7:0] I_1_t0b,
  input  [7:0] I_1_t1b,
  input  [7:0] I_2_t0b,
  input  [7:0] I_2_t1b,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  MapT_4 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  MapT_4 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t0b(other_ops_0_I_t0b),
    .I_t1b(other_ops_0_I_t1b),
    .O(other_ops_0_O)
  );
  MapT_4 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_t0b(other_ops_1_I_t0b),
    .I_t1b(other_ops_1_I_t1b),
    .O(other_ops_1_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t0b = I_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_t1b = I_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_t0b = I_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_t1b = I_2_t1b; // @[MapS.scala 20:41]
endmodule
module MapT_5(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  input  [7:0] I_1_t0b,
  input  [7:0] I_1_t1b,
  input  [7:0] I_2_t0b,
  input  [7:0] I_2_t1b,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_t0b; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_t1b; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_t0b; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_t1b; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_t0b; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_t1b; // @[MapT.scala 8:20]
  wire [7:0] op_O_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2; // @[MapT.scala 8:20]
  MapS_3 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_t0b(op_I_0_t0b),
    .I_0_t1b(op_I_0_t1b),
    .I_1_t0b(op_I_1_t0b),
    .I_1_t1b(op_I_1_t1b),
    .I_2_t0b(op_I_2_t0b),
    .I_2_t1b(op_I_2_t1b),
    .O_0(op_O_0),
    .O_1(op_O_1),
    .O_2(op_O_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign O_1 = op_O_1; // @[MapT.scala 15:7]
  assign O_2 = op_O_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_t0b = I_0_t0b; // @[MapT.scala 14:10]
  assign op_I_0_t1b = I_0_t1b; // @[MapT.scala 14:10]
  assign op_I_1_t0b = I_1_t0b; // @[MapT.scala 14:10]
  assign op_I_1_t1b = I_1_t1b; // @[MapT.scala 14:10]
  assign op_I_2_t0b = I_2_t0b; // @[MapT.scala 14:10]
  assign op_I_2_t1b = I_2_t1b; // @[MapT.scala 14:10]
endmodule
module AddNoValid(
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  assign O = I_t0b + I_t1b; // @[Arithmetic.scala 122:7]
endmodule
module ReduceT(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I,
  output [7:0] O
);
  wire  NestedCountersWithNumValid_CE; // @[ReduceT.scala 22:34]
  wire  NestedCountersWithNumValid_valid; // @[ReduceT.scala 22:34]
  wire [7:0] AddNoValid_I_t0b; // @[ReduceT.scala 25:25]
  wire [7:0] AddNoValid_I_t1b; // @[ReduceT.scala 25:25]
  wire [7:0] AddNoValid_O; // @[ReduceT.scala 25:25]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[Counter.scala 37:24]
  wire [1:0] _T_3; // @[Counter.scala 38:22]
  wire  _T_5; // @[ReduceT.scala 34:60]
  reg [7:0] _T_7; // @[ReduceT.scala 35:24]
  reg [31:0] _RAND_1;
  reg  _T_8; // @[ReduceT.scala 50:28]
  reg [31:0] _RAND_2;
  wire  _T_10; // @[ReduceT.scala 51:28]
  reg [7:0] _T_11; // @[ReduceT.scala 55:15]
  reg [31:0] _RAND_3;
  NestedCountersWithNumValid NestedCountersWithNumValid ( // @[ReduceT.scala 22:34]
    .CE(NestedCountersWithNumValid_CE),
    .valid(NestedCountersWithNumValid_valid)
  );
  AddNoValid AddNoValid ( // @[ReduceT.scala 25:25]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  assign _T_1 = value == 2'h2; // @[Counter.scala 37:24]
  assign _T_3 = value + 2'h1; // @[Counter.scala 38:22]
  assign _T_5 = value == 2'h0; // @[ReduceT.scala 34:60]
  assign _T_10 = _T_8 | _T_1; // @[ReduceT.scala 51:28]
  assign valid_down = _T_8; // @[ReduceT.scala 52:16]
  assign O = _T_11; // @[ReduceT.scala 55:5]
  assign NestedCountersWithNumValid_CE = valid_up; // @[ReduceT.scala 37:25]
  assign AddNoValid_I_t0b = I; // @[ReduceT.scala 43:55]
  assign AddNoValid_I_t1b = _T_7; // @[ReduceT.scala 44:55]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_7 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_8 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_11 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 2'h0;
    end else if (valid_up) begin
      if (_T_1) begin
        value <= 2'h0;
      end else begin
        value <= _T_3;
      end
    end
    if (NestedCountersWithNumValid_valid) begin
      if (_T_5) begin
        _T_7 <= I;
      end else begin
        _T_7 <= AddNoValid_O;
      end
    end
    if (reset) begin
      _T_8 <= 1'h0;
    end else begin
      _T_8 <= _T_10;
    end
    _T_11 <= AddNoValid_O;
  end
endmodule
module MapS_4(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  ReduceT fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I(fst_op_I),
    .O(fst_op_O)
  );
  ReduceT other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I(other_ops_0_I),
    .O(other_ops_0_O)
  );
  ReduceT other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I(other_ops_1_I),
    .O(other_ops_1_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I = I_0; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I = I_1; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I = I_2; // @[MapS.scala 20:41]
endmodule
module MapT_6(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2; // @[MapT.scala 8:20]
  MapS_4 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0(op_I_0),
    .I_1(op_I_1),
    .I_2(op_I_2),
    .O_0(op_O_0),
    .O_1(op_O_1),
    .O_2(op_O_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign O_1 = op_O_1; // @[MapT.scala 15:7]
  assign O_2 = op_O_2; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0 = I_0; // @[MapT.scala 14:10]
  assign op_I_1 = I_1; // @[MapT.scala 14:10]
  assign op_I_2 = I_2; // @[MapT.scala 14:10]
endmodule
module MapTNoValid(
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  wire [7:0] op_I_t0b; // @[MapT.scala 21:20]
  wire [7:0] op_I_t1b; // @[MapT.scala 21:20]
  wire [7:0] op_O; // @[MapT.scala 21:20]
  AddNoValid op ( // @[MapT.scala 21:20]
    .I_t0b(op_I_t0b),
    .I_t1b(op_I_t1b),
    .O(op_O)
  );
  assign O = op_O; // @[MapT.scala 27:7]
  assign op_I_t0b = I_t0b; // @[MapT.scala 26:10]
  assign op_I_t1b = I_t1b; // @[MapT.scala 26:10]
endmodule
module ReduceS(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O_0
);
  wire [7:0] MapTNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] MapTNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] MapTNoValid_O; // @[ReduceS.scala 20:43]
  wire [7:0] MapTNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] MapTNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] MapTNoValid_1_O; // @[ReduceS.scala 20:43]
  reg [7:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_1;
  MapTNoValid MapTNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(MapTNoValid_I_t0b),
    .I_t1b(MapTNoValid_I_t1b),
    .O(MapTNoValid_O)
  );
  MapTNoValid MapTNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(MapTNoValid_1_I_t0b),
    .I_t1b(MapTNoValid_1_I_t1b),
    .O(MapTNoValid_1_O)
  );
  assign valid_down = _T_1; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign MapTNoValid_I_t0b = I_2; // @[ReduceS.scala 43:18]
  assign MapTNoValid_I_t1b = MapTNoValid_1_O; // @[ReduceS.scala 36:18]
  assign MapTNoValid_1_I_t0b = I_1; // @[ReduceS.scala 43:18]
  assign MapTNoValid_1_I_t1b = I_0; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= MapTNoValid_O;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module MapT_7(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0; // @[MapT.scala 8:20]
  ReduceS op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0(op_I_0),
    .I_1(op_I_1),
    .I_2(op_I_2),
    .O_0(op_O_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0 = I_0; // @[MapT.scala 14:10]
  assign op_I_1 = I_1; // @[MapT.scala 14:10]
  assign op_I_2 = I_2; // @[MapT.scala 14:10]
endmodule
module ReduceT_1(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  output [7:0] O_0
);
  reg  _T; // @[ReduceT.scala 18:26]
  reg [31:0] _RAND_0;
  reg [7:0] _T_1_0; // @[ReduceT.scala 55:15]
  reg [31:0] _RAND_1;
  assign valid_down = _T; // @[ReduceT.scala 18:16]
  assign O_0 = _T_1_0; // @[ReduceT.scala 55:5]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1_0 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T <= 1'h0;
    end else begin
      _T <= valid_up;
    end
    _T_1_0 <= I_0;
  end
endmodule
module Passthrough_5(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  output [7:0] O
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O = I_0; // @[Passthrough.scala 17:68]
endmodule
module InitialDelayCounter_1(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [2:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [2:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 3'h7; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 3'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 3'h7; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 3'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Map2T_17(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_t0b,
  output [7:0] O_t1b
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_t0b; // @[Map2T.scala 8:20]
  wire [7:0] op_O_t1b; // @[Map2T.scala 8:20]
  Map2T_14 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0(op_I0),
    .I1(op_I1),
    .O_t0b(op_O_t0b),
    .O_t1b(op_O_t1b)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_t0b = op_O_t0b; // @[Map2T.scala 17:7]
  assign O_t1b = op_O_t1b; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0 = I0; // @[Map2T.scala 15:11]
  assign op_I1 = I1; // @[Map2T.scala 16:11]
endmodule
module RShift(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 272:14]
  assign O = I_t0b >> I_t1b; // @[Arithmetic.scala 270:7]
endmodule
module MapT_8(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_t0b; // @[MapT.scala 8:20]
  wire [7:0] op_I_t1b; // @[MapT.scala 8:20]
  wire [7:0] op_O; // @[MapT.scala 8:20]
  RShift op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_t0b(op_I_t0b),
    .I_t1b(op_I_t1b),
    .O(op_O)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O = op_O; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_t0b = I_t0b; // @[MapT.scala 14:10]
  assign op_I_t1b = I_t1b; // @[MapT.scala 14:10]
endmodule
module MapT_9(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_t0b; // @[MapT.scala 8:20]
  wire [7:0] op_I_t1b; // @[MapT.scala 8:20]
  wire [7:0] op_O; // @[MapT.scala 8:20]
  MapT_8 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_t0b(op_I_t0b),
    .I_t1b(op_I_t1b),
    .O(op_O)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O = op_O; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_t0b = I_t0b; // @[MapT.scala 14:10]
  assign op_I_t1b = I_t1b; // @[MapT.scala 14:10]
endmodule
module Module_0(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n91_valid_up; // @[Top.scala 17:21]
  wire  n91_valid_down; // @[Top.scala 17:21]
  wire [7:0] n91_I0_0; // @[Top.scala 17:21]
  wire [7:0] n91_I0_1; // @[Top.scala 17:21]
  wire [7:0] n91_I0_2; // @[Top.scala 17:21]
  wire [7:0] n91_I1_0; // @[Top.scala 17:21]
  wire [7:0] n91_I1_1; // @[Top.scala 17:21]
  wire [7:0] n91_I1_2; // @[Top.scala 17:21]
  wire [7:0] n91_O_0_t0b; // @[Top.scala 17:21]
  wire [7:0] n91_O_0_t1b; // @[Top.scala 17:21]
  wire [7:0] n91_O_1_t0b; // @[Top.scala 17:21]
  wire [7:0] n91_O_1_t1b; // @[Top.scala 17:21]
  wire [7:0] n91_O_2_t0b; // @[Top.scala 17:21]
  wire [7:0] n91_O_2_t1b; // @[Top.scala 17:21]
  wire  n107_valid_up; // @[Top.scala 21:22]
  wire  n107_valid_down; // @[Top.scala 21:22]
  wire [7:0] n107_I_0_t0b; // @[Top.scala 21:22]
  wire [7:0] n107_I_0_t1b; // @[Top.scala 21:22]
  wire [7:0] n107_I_1_t0b; // @[Top.scala 21:22]
  wire [7:0] n107_I_1_t1b; // @[Top.scala 21:22]
  wire [7:0] n107_I_2_t0b; // @[Top.scala 21:22]
  wire [7:0] n107_I_2_t1b; // @[Top.scala 21:22]
  wire [7:0] n107_O_0; // @[Top.scala 21:22]
  wire [7:0] n107_O_1; // @[Top.scala 21:22]
  wire [7:0] n107_O_2; // @[Top.scala 21:22]
  wire  n114_clock; // @[Top.scala 24:22]
  wire  n114_reset; // @[Top.scala 24:22]
  wire  n114_valid_up; // @[Top.scala 24:22]
  wire  n114_valid_down; // @[Top.scala 24:22]
  wire [7:0] n114_I_0; // @[Top.scala 24:22]
  wire [7:0] n114_I_1; // @[Top.scala 24:22]
  wire [7:0] n114_I_2; // @[Top.scala 24:22]
  wire [7:0] n114_O_0; // @[Top.scala 24:22]
  wire [7:0] n114_O_1; // @[Top.scala 24:22]
  wire [7:0] n114_O_2; // @[Top.scala 24:22]
  wire  n121_clock; // @[Top.scala 27:22]
  wire  n121_reset; // @[Top.scala 27:22]
  wire  n121_valid_up; // @[Top.scala 27:22]
  wire  n121_valid_down; // @[Top.scala 27:22]
  wire [7:0] n121_I_0; // @[Top.scala 27:22]
  wire [7:0] n121_I_1; // @[Top.scala 27:22]
  wire [7:0] n121_I_2; // @[Top.scala 27:22]
  wire [7:0] n121_O_0; // @[Top.scala 27:22]
  wire  n124_clock; // @[Top.scala 30:22]
  wire  n124_reset; // @[Top.scala 30:22]
  wire  n124_valid_up; // @[Top.scala 30:22]
  wire  n124_valid_down; // @[Top.scala 30:22]
  wire [7:0] n124_I_0; // @[Top.scala 30:22]
  wire [7:0] n124_O_0; // @[Top.scala 30:22]
  wire  n125_valid_up; // @[Top.scala 33:22]
  wire  n125_valid_down; // @[Top.scala 33:22]
  wire [7:0] n125_I_0; // @[Top.scala 33:22]
  wire [7:0] n125_O; // @[Top.scala 33:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n128_valid_up; // @[Top.scala 37:22]
  wire  n128_valid_down; // @[Top.scala 37:22]
  wire [7:0] n128_I0; // @[Top.scala 37:22]
  wire [7:0] n128_I1; // @[Top.scala 37:22]
  wire [7:0] n128_O_t0b; // @[Top.scala 37:22]
  wire [7:0] n128_O_t1b; // @[Top.scala 37:22]
  wire  n139_valid_up; // @[Top.scala 41:22]
  wire  n139_valid_down; // @[Top.scala 41:22]
  wire [7:0] n139_I_t0b; // @[Top.scala 41:22]
  wire [7:0] n139_I_t1b; // @[Top.scala 41:22]
  wire [7:0] n139_O; // @[Top.scala 41:22]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_4; // @[Counter.scala 37:24]
  wire [1:0] _T_6; // @[Counter.scala 38:22]
  wire [7:0] _GEN_5; // @[Const.scala 25:72]
  wire [7:0] _GEN_6; // @[Const.scala 25:72]
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  wire  _T_10; // @[Counter.scala 37:24]
  wire [1:0] _T_12; // @[Counter.scala 38:22]
  wire [7:0] _GEN_14; // @[Const.scala 25:72]
  InitialDelayCounter InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  Map2T_15 n91 ( // @[Top.scala 17:21]
    .valid_up(n91_valid_up),
    .valid_down(n91_valid_down),
    .I0_0(n91_I0_0),
    .I0_1(n91_I0_1),
    .I0_2(n91_I0_2),
    .I1_0(n91_I1_0),
    .I1_1(n91_I1_1),
    .I1_2(n91_I1_2),
    .O_0_t0b(n91_O_0_t0b),
    .O_0_t1b(n91_O_0_t1b),
    .O_1_t0b(n91_O_1_t0b),
    .O_1_t1b(n91_O_1_t1b),
    .O_2_t0b(n91_O_2_t0b),
    .O_2_t1b(n91_O_2_t1b)
  );
  MapT_5 n107 ( // @[Top.scala 21:22]
    .valid_up(n107_valid_up),
    .valid_down(n107_valid_down),
    .I_0_t0b(n107_I_0_t0b),
    .I_0_t1b(n107_I_0_t1b),
    .I_1_t0b(n107_I_1_t0b),
    .I_1_t1b(n107_I_1_t1b),
    .I_2_t0b(n107_I_2_t0b),
    .I_2_t1b(n107_I_2_t1b),
    .O_0(n107_O_0),
    .O_1(n107_O_1),
    .O_2(n107_O_2)
  );
  MapT_6 n114 ( // @[Top.scala 24:22]
    .clock(n114_clock),
    .reset(n114_reset),
    .valid_up(n114_valid_up),
    .valid_down(n114_valid_down),
    .I_0(n114_I_0),
    .I_1(n114_I_1),
    .I_2(n114_I_2),
    .O_0(n114_O_0),
    .O_1(n114_O_1),
    .O_2(n114_O_2)
  );
  MapT_7 n121 ( // @[Top.scala 27:22]
    .clock(n121_clock),
    .reset(n121_reset),
    .valid_up(n121_valid_up),
    .valid_down(n121_valid_down),
    .I_0(n121_I_0),
    .I_1(n121_I_1),
    .I_2(n121_I_2),
    .O_0(n121_O_0)
  );
  ReduceT_1 n124 ( // @[Top.scala 30:22]
    .clock(n124_clock),
    .reset(n124_reset),
    .valid_up(n124_valid_up),
    .valid_down(n124_valid_down),
    .I_0(n124_I_0),
    .O_0(n124_O_0)
  );
  Passthrough_5 n125 ( // @[Top.scala 33:22]
    .valid_up(n125_valid_up),
    .valid_down(n125_valid_down),
    .I_0(n125_I_0),
    .O(n125_O)
  );
  InitialDelayCounter_1 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  Map2T_17 n128 ( // @[Top.scala 37:22]
    .valid_up(n128_valid_up),
    .valid_down(n128_valid_down),
    .I0(n128_I0),
    .I1(n128_I1),
    .O_t0b(n128_O_t0b),
    .O_t1b(n128_O_t1b)
  );
  MapT_9 n139 ( // @[Top.scala 41:22]
    .valid_up(n139_valid_up),
    .valid_down(n139_valid_down),
    .I_t0b(n139_I_t0b),
    .I_t1b(n139_I_t1b),
    .O(n139_O)
  );
  assign _T_4 = value == 2'h2; // @[Counter.scala 37:24]
  assign _T_6 = value + 2'h1; // @[Counter.scala 38:22]
  assign _GEN_5 = 2'h1 == value ? 8'h1 : 8'h0; // @[Const.scala 25:72]
  assign _GEN_6 = 2'h1 == value ? 8'h2 : 8'h1; // @[Const.scala 25:72]
  assign _T_10 = value_1 == 2'h2; // @[Counter.scala 37:24]
  assign _T_12 = value_1 + 2'h1; // @[Counter.scala 38:22]
  assign _GEN_14 = 2'h1 == value_1 ? 8'h0 : 8'h4; // @[Const.scala 25:72]
  assign valid_down = n139_valid_down; // @[Top.scala 45:16]
  assign O = n139_O; // @[Top.scala 44:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n91_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 20:18]
  assign n91_I0_0 = I_0; // @[Top.scala 18:12]
  assign n91_I0_1 = I_1; // @[Top.scala 18:12]
  assign n91_I0_2 = I_2; // @[Top.scala 18:12]
  assign n91_I1_0 = 2'h2 == value ? 8'h0 : _GEN_5; // @[Top.scala 19:12]
  assign n91_I1_1 = 2'h2 == value ? 8'h1 : _GEN_6; // @[Top.scala 19:12]
  assign n91_I1_2 = 2'h2 == value ? 8'h0 : _GEN_5; // @[Top.scala 19:12]
  assign n107_valid_up = n91_valid_down; // @[Top.scala 23:19]
  assign n107_I_0_t0b = n91_O_0_t0b; // @[Top.scala 22:12]
  assign n107_I_0_t1b = n91_O_0_t1b; // @[Top.scala 22:12]
  assign n107_I_1_t0b = n91_O_1_t0b; // @[Top.scala 22:12]
  assign n107_I_1_t1b = n91_O_1_t1b; // @[Top.scala 22:12]
  assign n107_I_2_t0b = n91_O_2_t0b; // @[Top.scala 22:12]
  assign n107_I_2_t1b = n91_O_2_t1b; // @[Top.scala 22:12]
  assign n114_clock = clock;
  assign n114_reset = reset;
  assign n114_valid_up = n107_valid_down; // @[Top.scala 26:19]
  assign n114_I_0 = n107_O_0; // @[Top.scala 25:12]
  assign n114_I_1 = n107_O_1; // @[Top.scala 25:12]
  assign n114_I_2 = n107_O_2; // @[Top.scala 25:12]
  assign n121_clock = clock;
  assign n121_reset = reset;
  assign n121_valid_up = n114_valid_down; // @[Top.scala 29:19]
  assign n121_I_0 = n114_O_0; // @[Top.scala 28:12]
  assign n121_I_1 = n114_O_1; // @[Top.scala 28:12]
  assign n121_I_2 = n114_O_2; // @[Top.scala 28:12]
  assign n124_clock = clock;
  assign n124_reset = reset;
  assign n124_valid_up = n121_valid_down; // @[Top.scala 32:19]
  assign n124_I_0 = n121_O_0; // @[Top.scala 31:12]
  assign n125_valid_up = n124_valid_down; // @[Top.scala 35:19]
  assign n125_I_0 = n124_O_0; // @[Top.scala 34:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n128_valid_up = n125_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 40:19]
  assign n128_I0 = n125_O; // @[Top.scala 38:13]
  assign n128_I1 = 2'h2 == value_1 ? 8'h0 : _GEN_14; // @[Top.scala 39:13]
  assign n139_valid_up = n128_valid_down; // @[Top.scala 43:19]
  assign n139_I_t0b = n128_O_t0b; // @[Top.scala 42:12]
  assign n139_I_t1b = n128_O_t1b; // @[Top.scala 42:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value_1 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 2'h0;
    end else if (InitialDelayCounter_valid_down) begin
      if (_T_4) begin
        value <= 2'h0;
      end else begin
        value <= _T_6;
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (InitialDelayCounter_1_valid_down) begin
      if (_T_10) begin
        value_1 <= 2'h0;
      end else begin
        value_1 <= _T_12;
      end
    end
  end
endmodule
module MapT_10(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2; // @[MapT.scala 8:20]
  wire [7:0] op_O; // @[MapT.scala 8:20]
  Module_0 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0(op_I_0),
    .I_1(op_I_1),
    .I_2(op_I_2),
    .O(op_O)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O = op_O; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0 = I_0; // @[MapT.scala 14:10]
  assign op_I_1 = I_1; // @[MapT.scala 14:10]
  assign op_I_2 = I_2; // @[MapT.scala 14:10]
endmodule
module Passthrough_6(
  input        valid_up,
  output       valid_down,
  input  [7:0] I,
  output [7:0] O
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O = I; // @[Passthrough.scala 17:68]
endmodule
module Passthrough_7(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O_0_0,
  output [7:0] O_0_1
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0 = I_0; // @[Passthrough.scala 17:68]
  assign O_0_1 = I_1; // @[Passthrough.scala 17:68]
endmodule
module Serialize_3(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O
);
  wire  elem_counter_CE; // @[Serialize.scala 14:28]
  wire  elem_counter_valid; // @[Serialize.scala 14:28]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[Counter.scala 37:24]
  wire [1:0] _T_3; // @[Counter.scala 38:22]
  reg [7:0] mux_input_wire_1; // @[Serialize.scala 39:47]
  reg [31:0] _RAND_1;
  wire  _T_6; // @[Serialize.scala 42:34]
  wire  _T_7; // @[Serialize.scala 42:42]
  wire  _T_8; // @[Mux.scala 68:19]
  wire  _T_10; // @[Mux.scala 68:19]
  reg [7:0] _T_12; // @[Serialize.scala 53:15]
  reg [31:0] _RAND_2;
  reg  _T_13; // @[Serialize.scala 54:24]
  reg [31:0] _RAND_3;
  NestedCountersWithNumValid elem_counter ( // @[Serialize.scala 14:28]
    .CE(elem_counter_CE),
    .valid(elem_counter_valid)
  );
  assign _T_1 = value == 2'h2; // @[Counter.scala 37:24]
  assign _T_3 = value + 2'h1; // @[Counter.scala 38:22]
  assign _T_6 = value == 2'h0; // @[Serialize.scala 42:34]
  assign _T_7 = _T_6 & valid_up; // @[Serialize.scala 42:42]
  assign _T_8 = 2'h1 == value; // @[Mux.scala 68:19]
  assign _T_10 = 2'h0 == value; // @[Mux.scala 68:19]
  assign valid_down = _T_13; // @[Serialize.scala 54:14]
  assign O = _T_12; // @[Serialize.scala 53:5]
  assign elem_counter_CE = valid_up; // @[Serialize.scala 16:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mux_input_wire_1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_12 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_13 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 2'h0;
    end else if (valid_up) begin
      if (_T_1) begin
        value <= 2'h0;
      end else begin
        value <= _T_3;
      end
    end
    if (_T_7) begin
      mux_input_wire_1 <= I_1;
    end
    if (_T_10) begin
      _T_12 <= I_0;
    end else if (_T_8) begin
      _T_12 <= mux_input_wire_1;
    end else begin
      _T_12 <= I_0;
    end
    if (reset) begin
      _T_13 <= 1'h0;
    end else begin
      _T_13 <= valid_up;
    end
  end
endmodule
module MapS_5(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  output [7:0] O_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  Serialize_3 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
endmodule
module MapT_11(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  output [7:0] O_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0; // @[MapT.scala 8:20]
  MapS_5 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0(op_I_0_0),
    .I_0_1(op_I_0_1),
    .O_0(op_O_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0 = I_0_0; // @[MapT.scala 14:10]
  assign op_I_0_1 = I_0_1; // @[MapT.scala 14:10]
endmodule
module Passthrough_9(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  output [7:0] O_0_0,
  output [7:0] O_0_1
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0 = I_0_0; // @[Passthrough.scala 17:68]
  assign O_0_1 = I_0_1; // @[Passthrough.scala 17:68]
endmodule
module Passthrough_10(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  output [7:0] O_0,
  output [7:0] O_1
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0 = I_0_0; // @[Passthrough.scala 17:68]
  assign O_1 = I_0_1; // @[Passthrough.scala 17:68]
endmodule
module MapT_13(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  output [7:0] O_0,
  output [7:0] O_1
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1; // @[MapT.scala 8:20]
  Passthrough_10 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0(op_I_0_0),
    .I_0_1(op_I_0_1),
    .O_0(op_O_0),
    .O_1(op_O_1)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign O_1 = op_O_1; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0 = I_0_0; // @[MapT.scala 14:10]
  assign op_I_0_1 = I_0_1; // @[MapT.scala 14:10]
endmodule
module InitialDelayCounter_2(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [3:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [3:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 4'h8; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 4'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 4'h8; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 4'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Map2S_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  output [7:0] O_0_t0b,
  output [7:0] O_0_t1b,
  output [7:0] O_1_t0b,
  output [7:0] O_1_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  Map2T_14 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  Map2T_14 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
endmodule
module Map2T_24(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  output [7:0] O_0_t0b,
  output [7:0] O_0_t1b,
  output [7:0] O_1_t0b,
  output [7:0] O_1_t1b
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_t0b; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_t1b; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_t0b; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_t1b; // @[Map2T.scala 8:20]
  Map2S_4 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .O_0_t0b(op_O_0_t0b),
    .O_0_t1b(op_O_0_t1b),
    .O_1_t0b(op_O_1_t0b),
    .O_1_t1b(op_O_1_t1b)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_t0b = op_O_0_t0b; // @[Map2T.scala 17:7]
  assign O_0_t1b = op_O_0_t1b; // @[Map2T.scala 17:7]
  assign O_1_t0b = op_O_1_t0b; // @[Map2T.scala 17:7]
  assign O_1_t1b = op_O_1_t1b; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
endmodule
module MapS_7(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  input  [7:0] I_1_t0b,
  input  [7:0] I_1_t1b,
  output [7:0] O_0,
  output [7:0] O_1
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O; // @[MapS.scala 10:86]
  MapT_4 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  MapT_4 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t0b(other_ops_0_I_t0b),
    .I_t1b(other_ops_0_I_t1b),
    .O(other_ops_0_O)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t0b = I_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_t1b = I_1_t1b; // @[MapS.scala 20:41]
endmodule
module MapT_15(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  input  [7:0] I_1_t0b,
  input  [7:0] I_1_t1b,
  output [7:0] O_0,
  output [7:0] O_1
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_t0b; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_t1b; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_t0b; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_t1b; // @[MapT.scala 8:20]
  wire [7:0] op_O_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1; // @[MapT.scala 8:20]
  MapS_7 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_t0b(op_I_0_t0b),
    .I_0_t1b(op_I_0_t1b),
    .I_1_t0b(op_I_1_t0b),
    .I_1_t1b(op_I_1_t1b),
    .O_0(op_O_0),
    .O_1(op_O_1)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign O_1 = op_O_1; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_t0b = I_0_t0b; // @[MapT.scala 14:10]
  assign op_I_0_t1b = I_0_t1b; // @[MapT.scala 14:10]
  assign op_I_1_t0b = I_1_t0b; // @[MapT.scala 14:10]
  assign op_I_1_t1b = I_1_t1b; // @[MapT.scala 14:10]
endmodule
module ReduceT_2(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I,
  output [7:0] O
);
  wire  NestedCountersWithNumValid_CE; // @[ReduceT.scala 22:34]
  wire  NestedCountersWithNumValid_valid; // @[ReduceT.scala 22:34]
  wire [7:0] AddNoValid_I_t0b; // @[ReduceT.scala 25:25]
  wire [7:0] AddNoValid_I_t1b; // @[ReduceT.scala 25:25]
  wire [7:0] AddNoValid_O; // @[ReduceT.scala 25:25]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[Counter.scala 37:24]
  wire [1:0] _T_3; // @[Counter.scala 38:22]
  wire  _T_5; // @[ReduceT.scala 34:60]
  reg [7:0] _T_7; // @[ReduceT.scala 35:24]
  reg [31:0] _RAND_1;
  reg  _T_8; // @[ReduceT.scala 50:28]
  reg [31:0] _RAND_2;
  wire  _T_9; // @[ReduceT.scala 51:51]
  wire  _T_10; // @[ReduceT.scala 51:28]
  reg [7:0] _T_11; // @[ReduceT.scala 55:15]
  reg [31:0] _RAND_3;
  NestedCountersWithNumValid NestedCountersWithNumValid ( // @[ReduceT.scala 22:34]
    .CE(NestedCountersWithNumValid_CE),
    .valid(NestedCountersWithNumValid_valid)
  );
  AddNoValid AddNoValid ( // @[ReduceT.scala 25:25]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  assign _T_1 = value == 2'h2; // @[Counter.scala 37:24]
  assign _T_3 = value + 2'h1; // @[Counter.scala 38:22]
  assign _T_5 = value == 2'h0; // @[ReduceT.scala 34:60]
  assign _T_9 = value == 2'h1; // @[ReduceT.scala 51:51]
  assign _T_10 = _T_8 | _T_9; // @[ReduceT.scala 51:28]
  assign valid_down = _T_8; // @[ReduceT.scala 52:16]
  assign O = _T_11; // @[ReduceT.scala 55:5]
  assign NestedCountersWithNumValid_CE = valid_up; // @[ReduceT.scala 37:25]
  assign AddNoValid_I_t0b = I; // @[ReduceT.scala 43:55]
  assign AddNoValid_I_t1b = _T_7; // @[ReduceT.scala 44:55]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_7 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_8 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_11 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 2'h0;
    end else if (valid_up) begin
      if (_T_1) begin
        value <= 2'h0;
      end else begin
        value <= _T_3;
      end
    end
    if (NestedCountersWithNumValid_valid) begin
      if (_T_5) begin
        _T_7 <= I;
      end else begin
        _T_7 <= AddNoValid_O;
      end
    end
    if (reset) begin
      _T_8 <= 1'h0;
    end else begin
      _T_8 <= _T_10;
    end
    _T_11 <= AddNoValid_O;
  end
endmodule
module MapS_8(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O_0,
  output [7:0] O_1
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O; // @[MapS.scala 10:86]
  ReduceT_2 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I(fst_op_I),
    .O(fst_op_O)
  );
  ReduceT_2 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I(other_ops_0_I),
    .O(other_ops_0_O)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I = I_0; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I = I_1; // @[MapS.scala 20:41]
endmodule
module MapT_16(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O_0,
  output [7:0] O_1
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1; // @[MapT.scala 8:20]
  MapS_8 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0(op_I_0),
    .I_1(op_I_1),
    .O_0(op_O_0),
    .O_1(op_O_1)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign O_1 = op_O_1; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0 = I_0; // @[MapT.scala 14:10]
  assign op_I_1 = I_1; // @[MapT.scala 14:10]
endmodule
module ReduceS_1(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O_0
);
  wire [7:0] MapTNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] MapTNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] MapTNoValid_O; // @[ReduceS.scala 20:43]
  reg [7:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_1;
  MapTNoValid MapTNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(MapTNoValid_I_t0b),
    .I_t1b(MapTNoValid_I_t1b),
    .O(MapTNoValid_O)
  );
  assign valid_down = _T_1; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign MapTNoValid_I_t0b = I_0; // @[ReduceS.scala 43:18]
  assign MapTNoValid_I_t1b = I_1; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= MapTNoValid_O;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module MapT_17(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0; // @[MapT.scala 8:20]
  ReduceS_1 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0(op_I_0),
    .I_1(op_I_1),
    .O_0(op_O_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0 = I_0; // @[MapT.scala 14:10]
  assign op_I_1 = I_1; // @[MapT.scala 14:10]
endmodule
module InitialDelayCounter_3(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [3:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [3:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 4'hc; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 4'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 4'hc; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 4'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Module_1(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n185_valid_up; // @[Top.scala 52:22]
  wire  n185_valid_down; // @[Top.scala 52:22]
  wire [7:0] n185_I0_0; // @[Top.scala 52:22]
  wire [7:0] n185_I0_1; // @[Top.scala 52:22]
  wire [7:0] n185_I1_0; // @[Top.scala 52:22]
  wire [7:0] n185_I1_1; // @[Top.scala 52:22]
  wire [7:0] n185_O_0_t0b; // @[Top.scala 52:22]
  wire [7:0] n185_O_0_t1b; // @[Top.scala 52:22]
  wire [7:0] n185_O_1_t0b; // @[Top.scala 52:22]
  wire [7:0] n185_O_1_t1b; // @[Top.scala 52:22]
  wire  n201_valid_up; // @[Top.scala 56:22]
  wire  n201_valid_down; // @[Top.scala 56:22]
  wire [7:0] n201_I_0_t0b; // @[Top.scala 56:22]
  wire [7:0] n201_I_0_t1b; // @[Top.scala 56:22]
  wire [7:0] n201_I_1_t0b; // @[Top.scala 56:22]
  wire [7:0] n201_I_1_t1b; // @[Top.scala 56:22]
  wire [7:0] n201_O_0; // @[Top.scala 56:22]
  wire [7:0] n201_O_1; // @[Top.scala 56:22]
  wire  n208_clock; // @[Top.scala 59:22]
  wire  n208_reset; // @[Top.scala 59:22]
  wire  n208_valid_up; // @[Top.scala 59:22]
  wire  n208_valid_down; // @[Top.scala 59:22]
  wire [7:0] n208_I_0; // @[Top.scala 59:22]
  wire [7:0] n208_I_1; // @[Top.scala 59:22]
  wire [7:0] n208_O_0; // @[Top.scala 59:22]
  wire [7:0] n208_O_1; // @[Top.scala 59:22]
  wire  n215_clock; // @[Top.scala 62:22]
  wire  n215_reset; // @[Top.scala 62:22]
  wire  n215_valid_up; // @[Top.scala 62:22]
  wire  n215_valid_down; // @[Top.scala 62:22]
  wire [7:0] n215_I_0; // @[Top.scala 62:22]
  wire [7:0] n215_I_1; // @[Top.scala 62:22]
  wire [7:0] n215_O_0; // @[Top.scala 62:22]
  wire  n218_clock; // @[Top.scala 65:22]
  wire  n218_reset; // @[Top.scala 65:22]
  wire  n218_valid_up; // @[Top.scala 65:22]
  wire  n218_valid_down; // @[Top.scala 65:22]
  wire [7:0] n218_I_0; // @[Top.scala 65:22]
  wire [7:0] n218_O_0; // @[Top.scala 65:22]
  wire  n219_valid_up; // @[Top.scala 68:22]
  wire  n219_valid_down; // @[Top.scala 68:22]
  wire [7:0] n219_I_0; // @[Top.scala 68:22]
  wire [7:0] n219_O; // @[Top.scala 68:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n222_valid_up; // @[Top.scala 72:22]
  wire  n222_valid_down; // @[Top.scala 72:22]
  wire [7:0] n222_I0; // @[Top.scala 72:22]
  wire [7:0] n222_I1; // @[Top.scala 72:22]
  wire [7:0] n222_O_t0b; // @[Top.scala 72:22]
  wire [7:0] n222_O_t1b; // @[Top.scala 72:22]
  wire  n233_valid_up; // @[Top.scala 76:22]
  wire  n233_valid_down; // @[Top.scala 76:22]
  wire [7:0] n233_I_t0b; // @[Top.scala 76:22]
  wire [7:0] n233_I_t1b; // @[Top.scala 76:22]
  wire [7:0] n233_O; // @[Top.scala 76:22]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_4; // @[Counter.scala 37:24]
  wire [1:0] _T_6; // @[Counter.scala 38:22]
  wire [7:0] _GEN_4; // @[Const.scala 25:72]
  wire [7:0] _GEN_5; // @[Const.scala 25:72]
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  wire  _T_10; // @[Counter.scala 37:24]
  wire [1:0] _T_12; // @[Counter.scala 38:22]
  wire [7:0] _GEN_11; // @[Const.scala 25:72]
  InitialDelayCounter_2 InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  Map2T_24 n185 ( // @[Top.scala 52:22]
    .valid_up(n185_valid_up),
    .valid_down(n185_valid_down),
    .I0_0(n185_I0_0),
    .I0_1(n185_I0_1),
    .I1_0(n185_I1_0),
    .I1_1(n185_I1_1),
    .O_0_t0b(n185_O_0_t0b),
    .O_0_t1b(n185_O_0_t1b),
    .O_1_t0b(n185_O_1_t0b),
    .O_1_t1b(n185_O_1_t1b)
  );
  MapT_15 n201 ( // @[Top.scala 56:22]
    .valid_up(n201_valid_up),
    .valid_down(n201_valid_down),
    .I_0_t0b(n201_I_0_t0b),
    .I_0_t1b(n201_I_0_t1b),
    .I_1_t0b(n201_I_1_t0b),
    .I_1_t1b(n201_I_1_t1b),
    .O_0(n201_O_0),
    .O_1(n201_O_1)
  );
  MapT_16 n208 ( // @[Top.scala 59:22]
    .clock(n208_clock),
    .reset(n208_reset),
    .valid_up(n208_valid_up),
    .valid_down(n208_valid_down),
    .I_0(n208_I_0),
    .I_1(n208_I_1),
    .O_0(n208_O_0),
    .O_1(n208_O_1)
  );
  MapT_17 n215 ( // @[Top.scala 62:22]
    .clock(n215_clock),
    .reset(n215_reset),
    .valid_up(n215_valid_up),
    .valid_down(n215_valid_down),
    .I_0(n215_I_0),
    .I_1(n215_I_1),
    .O_0(n215_O_0)
  );
  ReduceT_1 n218 ( // @[Top.scala 65:22]
    .clock(n218_clock),
    .reset(n218_reset),
    .valid_up(n218_valid_up),
    .valid_down(n218_valid_down),
    .I_0(n218_I_0),
    .O_0(n218_O_0)
  );
  Passthrough_5 n219 ( // @[Top.scala 68:22]
    .valid_up(n219_valid_up),
    .valid_down(n219_valid_down),
    .I_0(n219_I_0),
    .O(n219_O)
  );
  InitialDelayCounter_3 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  Map2T_17 n222 ( // @[Top.scala 72:22]
    .valid_up(n222_valid_up),
    .valid_down(n222_valid_down),
    .I0(n222_I0),
    .I1(n222_I1),
    .O_t0b(n222_O_t0b),
    .O_t1b(n222_O_t1b)
  );
  MapT_9 n233 ( // @[Top.scala 76:22]
    .valid_up(n233_valid_up),
    .valid_down(n233_valid_down),
    .I_t0b(n233_I_t0b),
    .I_t1b(n233_I_t1b),
    .O(n233_O)
  );
  assign _T_4 = value == 2'h2; // @[Counter.scala 37:24]
  assign _T_6 = value + 2'h1; // @[Counter.scala 38:22]
  assign _GEN_4 = 2'h1 == value ? 8'h2 : 8'h0; // @[Const.scala 25:72]
  assign _GEN_5 = 2'h1 == value ? 8'h0 : 8'h1; // @[Const.scala 25:72]
  assign _T_10 = value_1 == 2'h2; // @[Counter.scala 37:24]
  assign _T_12 = value_1 + 2'h1; // @[Counter.scala 38:22]
  assign _GEN_11 = 2'h1 == value_1 ? 8'h0 : 8'h3; // @[Const.scala 25:72]
  assign valid_down = n233_valid_down; // @[Top.scala 80:16]
  assign O = n233_O; // @[Top.scala 79:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n185_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 55:19]
  assign n185_I0_0 = I_0; // @[Top.scala 53:13]
  assign n185_I0_1 = I_1; // @[Top.scala 53:13]
  assign n185_I1_0 = 2'h2 == value ? 8'h1 : _GEN_4; // @[Top.scala 54:13]
  assign n185_I1_1 = 2'h2 == value ? 8'h0 : _GEN_5; // @[Top.scala 54:13]
  assign n201_valid_up = n185_valid_down; // @[Top.scala 58:19]
  assign n201_I_0_t0b = n185_O_0_t0b; // @[Top.scala 57:12]
  assign n201_I_0_t1b = n185_O_0_t1b; // @[Top.scala 57:12]
  assign n201_I_1_t0b = n185_O_1_t0b; // @[Top.scala 57:12]
  assign n201_I_1_t1b = n185_O_1_t1b; // @[Top.scala 57:12]
  assign n208_clock = clock;
  assign n208_reset = reset;
  assign n208_valid_up = n201_valid_down; // @[Top.scala 61:19]
  assign n208_I_0 = n201_O_0; // @[Top.scala 60:12]
  assign n208_I_1 = n201_O_1; // @[Top.scala 60:12]
  assign n215_clock = clock;
  assign n215_reset = reset;
  assign n215_valid_up = n208_valid_down; // @[Top.scala 64:19]
  assign n215_I_0 = n208_O_0; // @[Top.scala 63:12]
  assign n215_I_1 = n208_O_1; // @[Top.scala 63:12]
  assign n218_clock = clock;
  assign n218_reset = reset;
  assign n218_valid_up = n215_valid_down; // @[Top.scala 67:19]
  assign n218_I_0 = n215_O_0; // @[Top.scala 66:12]
  assign n219_valid_up = n218_valid_down; // @[Top.scala 70:19]
  assign n219_I_0 = n218_O_0; // @[Top.scala 69:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n222_valid_up = n219_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 75:19]
  assign n222_I0 = n219_O; // @[Top.scala 73:13]
  assign n222_I1 = 2'h2 == value_1 ? 8'h0 : _GEN_11; // @[Top.scala 74:13]
  assign n233_valid_up = n222_valid_down; // @[Top.scala 78:19]
  assign n233_I_t0b = n222_O_t0b; // @[Top.scala 77:12]
  assign n233_I_t1b = n222_O_t1b; // @[Top.scala 77:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value_1 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 2'h0;
    end else if (InitialDelayCounter_valid_down) begin
      if (_T_4) begin
        value <= 2'h0;
      end else begin
        value <= _T_6;
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (InitialDelayCounter_1_valid_down) begin
      if (_T_10) begin
        value_1 <= 2'h0;
      end else begin
        value_1 <= _T_12;
      end
    end
  end
endmodule
module MapT_20(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1; // @[MapT.scala 8:20]
  wire [7:0] op_O; // @[MapT.scala 8:20]
  Module_1 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0(op_I_0),
    .I_1(op_I_1),
    .O(op_O)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O = op_O; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0 = I_0; // @[MapT.scala 14:10]
  assign op_I_1 = I_1; // @[MapT.scala 14:10]
endmodule
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I,
  output [7:0] O
);
  wire  n1_clock; // @[Top.scala 86:20]
  wire  n1_reset; // @[Top.scala 86:20]
  wire  n1_valid_up; // @[Top.scala 86:20]
  wire  n1_valid_down; // @[Top.scala 86:20]
  wire [7:0] n1_I; // @[Top.scala 86:20]
  wire [7:0] n1_O; // @[Top.scala 86:20]
  wire  n2_clock; // @[Top.scala 89:20]
  wire  n2_reset; // @[Top.scala 89:20]
  wire  n2_valid_up; // @[Top.scala 89:20]
  wire  n2_valid_down; // @[Top.scala 89:20]
  wire [7:0] n2_I; // @[Top.scala 89:20]
  wire [7:0] n2_O; // @[Top.scala 89:20]
  wire  n3_clock; // @[Top.scala 92:20]
  wire  n3_reset; // @[Top.scala 92:20]
  wire  n3_valid_up; // @[Top.scala 92:20]
  wire  n3_valid_down; // @[Top.scala 92:20]
  wire [7:0] n3_I; // @[Top.scala 92:20]
  wire [7:0] n3_O; // @[Top.scala 92:20]
  wire  n4_clock; // @[Top.scala 95:20]
  wire  n4_reset; // @[Top.scala 95:20]
  wire  n4_valid_up; // @[Top.scala 95:20]
  wire  n4_valid_down; // @[Top.scala 95:20]
  wire [7:0] n4_I; // @[Top.scala 95:20]
  wire [7:0] n4_O; // @[Top.scala 95:20]
  wire  n5_clock; // @[Top.scala 98:20]
  wire  n5_reset; // @[Top.scala 98:20]
  wire  n5_valid_up; // @[Top.scala 98:20]
  wire  n5_valid_down; // @[Top.scala 98:20]
  wire [7:0] n5_I; // @[Top.scala 98:20]
  wire [7:0] n5_O; // @[Top.scala 98:20]
  wire  n6_valid_up; // @[Top.scala 101:20]
  wire  n6_valid_down; // @[Top.scala 101:20]
  wire [7:0] n6_I0; // @[Top.scala 101:20]
  wire [7:0] n6_I1; // @[Top.scala 101:20]
  wire [7:0] n6_O_0; // @[Top.scala 101:20]
  wire [7:0] n6_O_1; // @[Top.scala 101:20]
  wire  n13_valid_up; // @[Top.scala 105:21]
  wire  n13_valid_down; // @[Top.scala 105:21]
  wire [7:0] n13_I0_0; // @[Top.scala 105:21]
  wire [7:0] n13_I0_1; // @[Top.scala 105:21]
  wire [7:0] n13_I1; // @[Top.scala 105:21]
  wire [7:0] n13_O_0; // @[Top.scala 105:21]
  wire [7:0] n13_O_1; // @[Top.scala 105:21]
  wire [7:0] n13_O_2; // @[Top.scala 105:21]
  wire  n20_valid_up; // @[Top.scala 109:21]
  wire  n20_valid_down; // @[Top.scala 109:21]
  wire [7:0] n20_I_0; // @[Top.scala 109:21]
  wire [7:0] n20_I_1; // @[Top.scala 109:21]
  wire [7:0] n20_I_2; // @[Top.scala 109:21]
  wire [7:0] n20_O_0_0; // @[Top.scala 109:21]
  wire [7:0] n20_O_0_1; // @[Top.scala 109:21]
  wire [7:0] n20_O_0_2; // @[Top.scala 109:21]
  wire  n25_clock; // @[Top.scala 112:21]
  wire  n25_reset; // @[Top.scala 112:21]
  wire  n25_valid_up; // @[Top.scala 112:21]
  wire  n25_valid_down; // @[Top.scala 112:21]
  wire [7:0] n25_I_0_0; // @[Top.scala 112:21]
  wire [7:0] n25_I_0_1; // @[Top.scala 112:21]
  wire [7:0] n25_I_0_2; // @[Top.scala 112:21]
  wire [7:0] n25_O_0; // @[Top.scala 112:21]
  wire  n26_clock; // @[Top.scala 115:21]
  wire  n26_reset; // @[Top.scala 115:21]
  wire  n26_valid_up; // @[Top.scala 115:21]
  wire  n26_valid_down; // @[Top.scala 115:21]
  wire [7:0] n26_I; // @[Top.scala 115:21]
  wire [7:0] n26_O; // @[Top.scala 115:21]
  wire  n27_clock; // @[Top.scala 118:21]
  wire  n27_reset; // @[Top.scala 118:21]
  wire  n27_valid_up; // @[Top.scala 118:21]
  wire  n27_valid_down; // @[Top.scala 118:21]
  wire [7:0] n27_I; // @[Top.scala 118:21]
  wire [7:0] n27_O; // @[Top.scala 118:21]
  wire  n28_valid_up; // @[Top.scala 121:21]
  wire  n28_valid_down; // @[Top.scala 121:21]
  wire [7:0] n28_I0; // @[Top.scala 121:21]
  wire [7:0] n28_I1; // @[Top.scala 121:21]
  wire [7:0] n28_O_0; // @[Top.scala 121:21]
  wire [7:0] n28_O_1; // @[Top.scala 121:21]
  wire  n35_valid_up; // @[Top.scala 125:21]
  wire  n35_valid_down; // @[Top.scala 125:21]
  wire [7:0] n35_I0_0; // @[Top.scala 125:21]
  wire [7:0] n35_I0_1; // @[Top.scala 125:21]
  wire [7:0] n35_I1; // @[Top.scala 125:21]
  wire [7:0] n35_O_0; // @[Top.scala 125:21]
  wire [7:0] n35_O_1; // @[Top.scala 125:21]
  wire [7:0] n35_O_2; // @[Top.scala 125:21]
  wire  n42_valid_up; // @[Top.scala 129:21]
  wire  n42_valid_down; // @[Top.scala 129:21]
  wire [7:0] n42_I_0; // @[Top.scala 129:21]
  wire [7:0] n42_I_1; // @[Top.scala 129:21]
  wire [7:0] n42_I_2; // @[Top.scala 129:21]
  wire [7:0] n42_O_0_0; // @[Top.scala 129:21]
  wire [7:0] n42_O_0_1; // @[Top.scala 129:21]
  wire [7:0] n42_O_0_2; // @[Top.scala 129:21]
  wire  n47_clock; // @[Top.scala 132:21]
  wire  n47_reset; // @[Top.scala 132:21]
  wire  n47_valid_up; // @[Top.scala 132:21]
  wire  n47_valid_down; // @[Top.scala 132:21]
  wire [7:0] n47_I_0_0; // @[Top.scala 132:21]
  wire [7:0] n47_I_0_1; // @[Top.scala 132:21]
  wire [7:0] n47_I_0_2; // @[Top.scala 132:21]
  wire [7:0] n47_O_0; // @[Top.scala 132:21]
  wire  n48_valid_up; // @[Top.scala 135:21]
  wire  n48_valid_down; // @[Top.scala 135:21]
  wire [7:0] n48_I0_0; // @[Top.scala 135:21]
  wire [7:0] n48_I1_0; // @[Top.scala 135:21]
  wire [7:0] n48_O_0_0; // @[Top.scala 135:21]
  wire [7:0] n48_O_0_1; // @[Top.scala 135:21]
  wire  n55_clock; // @[Top.scala 139:21]
  wire  n55_reset; // @[Top.scala 139:21]
  wire  n55_valid_up; // @[Top.scala 139:21]
  wire  n55_valid_down; // @[Top.scala 139:21]
  wire [7:0] n55_I; // @[Top.scala 139:21]
  wire [7:0] n55_O; // @[Top.scala 139:21]
  wire  n56_clock; // @[Top.scala 142:21]
  wire  n56_reset; // @[Top.scala 142:21]
  wire  n56_valid_up; // @[Top.scala 142:21]
  wire  n56_valid_down; // @[Top.scala 142:21]
  wire [7:0] n56_I; // @[Top.scala 142:21]
  wire [7:0] n56_O; // @[Top.scala 142:21]
  wire  n57_valid_up; // @[Top.scala 145:21]
  wire  n57_valid_down; // @[Top.scala 145:21]
  wire [7:0] n57_I0; // @[Top.scala 145:21]
  wire [7:0] n57_I1; // @[Top.scala 145:21]
  wire [7:0] n57_O_0; // @[Top.scala 145:21]
  wire [7:0] n57_O_1; // @[Top.scala 145:21]
  wire  n64_valid_up; // @[Top.scala 149:21]
  wire  n64_valid_down; // @[Top.scala 149:21]
  wire [7:0] n64_I0_0; // @[Top.scala 149:21]
  wire [7:0] n64_I0_1; // @[Top.scala 149:21]
  wire [7:0] n64_I1; // @[Top.scala 149:21]
  wire [7:0] n64_O_0; // @[Top.scala 149:21]
  wire [7:0] n64_O_1; // @[Top.scala 149:21]
  wire [7:0] n64_O_2; // @[Top.scala 149:21]
  wire  n71_valid_up; // @[Top.scala 153:21]
  wire  n71_valid_down; // @[Top.scala 153:21]
  wire [7:0] n71_I_0; // @[Top.scala 153:21]
  wire [7:0] n71_I_1; // @[Top.scala 153:21]
  wire [7:0] n71_I_2; // @[Top.scala 153:21]
  wire [7:0] n71_O_0_0; // @[Top.scala 153:21]
  wire [7:0] n71_O_0_1; // @[Top.scala 153:21]
  wire [7:0] n71_O_0_2; // @[Top.scala 153:21]
  wire  n76_clock; // @[Top.scala 156:21]
  wire  n76_reset; // @[Top.scala 156:21]
  wire  n76_valid_up; // @[Top.scala 156:21]
  wire  n76_valid_down; // @[Top.scala 156:21]
  wire [7:0] n76_I_0_0; // @[Top.scala 156:21]
  wire [7:0] n76_I_0_1; // @[Top.scala 156:21]
  wire [7:0] n76_I_0_2; // @[Top.scala 156:21]
  wire [7:0] n76_O_0; // @[Top.scala 156:21]
  wire  n77_valid_up; // @[Top.scala 159:21]
  wire  n77_valid_down; // @[Top.scala 159:21]
  wire [7:0] n77_I0_0_0; // @[Top.scala 159:21]
  wire [7:0] n77_I0_0_1; // @[Top.scala 159:21]
  wire [7:0] n77_I1_0; // @[Top.scala 159:21]
  wire [7:0] n77_O_0_0; // @[Top.scala 159:21]
  wire [7:0] n77_O_0_1; // @[Top.scala 159:21]
  wire [7:0] n77_O_0_2; // @[Top.scala 159:21]
  wire  n84_valid_up; // @[Top.scala 163:21]
  wire  n84_valid_down; // @[Top.scala 163:21]
  wire [7:0] n84_I_0_0; // @[Top.scala 163:21]
  wire [7:0] n84_I_0_1; // @[Top.scala 163:21]
  wire [7:0] n84_I_0_2; // @[Top.scala 163:21]
  wire [7:0] n84_O_0_0; // @[Top.scala 163:21]
  wire [7:0] n84_O_0_1; // @[Top.scala 163:21]
  wire [7:0] n84_O_0_2; // @[Top.scala 163:21]
  wire  n87_valid_up; // @[Top.scala 166:21]
  wire  n87_valid_down; // @[Top.scala 166:21]
  wire [7:0] n87_I_0_0; // @[Top.scala 166:21]
  wire [7:0] n87_I_0_1; // @[Top.scala 166:21]
  wire [7:0] n87_I_0_2; // @[Top.scala 166:21]
  wire [7:0] n87_O_0; // @[Top.scala 166:21]
  wire [7:0] n87_O_1; // @[Top.scala 166:21]
  wire [7:0] n87_O_2; // @[Top.scala 166:21]
  wire  n140_clock; // @[Top.scala 169:22]
  wire  n140_reset; // @[Top.scala 169:22]
  wire  n140_valid_up; // @[Top.scala 169:22]
  wire  n140_valid_down; // @[Top.scala 169:22]
  wire [7:0] n140_I_0; // @[Top.scala 169:22]
  wire [7:0] n140_I_1; // @[Top.scala 169:22]
  wire [7:0] n140_I_2; // @[Top.scala 169:22]
  wire [7:0] n140_O; // @[Top.scala 169:22]
  wire  n141_valid_up; // @[Top.scala 172:22]
  wire  n141_valid_down; // @[Top.scala 172:22]
  wire [7:0] n141_I; // @[Top.scala 172:22]
  wire [7:0] n141_O; // @[Top.scala 172:22]
  wire  n142_clock; // @[Top.scala 175:22]
  wire  n142_reset; // @[Top.scala 175:22]
  wire  n142_valid_up; // @[Top.scala 175:22]
  wire  n142_valid_down; // @[Top.scala 175:22]
  wire [7:0] n142_I; // @[Top.scala 175:22]
  wire [7:0] n142_O; // @[Top.scala 175:22]
  wire  n143_clock; // @[Top.scala 178:22]
  wire  n143_reset; // @[Top.scala 178:22]
  wire  n143_valid_up; // @[Top.scala 178:22]
  wire  n143_valid_down; // @[Top.scala 178:22]
  wire [7:0] n143_I; // @[Top.scala 178:22]
  wire [7:0] n143_O; // @[Top.scala 178:22]
  wire  n144_valid_up; // @[Top.scala 181:22]
  wire  n144_valid_down; // @[Top.scala 181:22]
  wire [7:0] n144_I0; // @[Top.scala 181:22]
  wire [7:0] n144_I1; // @[Top.scala 181:22]
  wire [7:0] n144_O_0; // @[Top.scala 181:22]
  wire [7:0] n144_O_1; // @[Top.scala 181:22]
  wire  n151_valid_up; // @[Top.scala 185:22]
  wire  n151_valid_down; // @[Top.scala 185:22]
  wire [7:0] n151_I_0; // @[Top.scala 185:22]
  wire [7:0] n151_I_1; // @[Top.scala 185:22]
  wire [7:0] n151_O_0_0; // @[Top.scala 185:22]
  wire [7:0] n151_O_0_1; // @[Top.scala 185:22]
  wire  n156_clock; // @[Top.scala 188:22]
  wire  n156_reset; // @[Top.scala 188:22]
  wire  n156_valid_up; // @[Top.scala 188:22]
  wire  n156_valid_down; // @[Top.scala 188:22]
  wire [7:0] n156_I_0_0; // @[Top.scala 188:22]
  wire [7:0] n156_I_0_1; // @[Top.scala 188:22]
  wire [7:0] n156_O_0; // @[Top.scala 188:22]
  wire  n157_clock; // @[Top.scala 191:22]
  wire  n157_reset; // @[Top.scala 191:22]
  wire  n157_valid_up; // @[Top.scala 191:22]
  wire  n157_valid_down; // @[Top.scala 191:22]
  wire [7:0] n157_I; // @[Top.scala 191:22]
  wire [7:0] n157_O; // @[Top.scala 191:22]
  wire  n158_valid_up; // @[Top.scala 194:22]
  wire  n158_valid_down; // @[Top.scala 194:22]
  wire [7:0] n158_I0; // @[Top.scala 194:22]
  wire [7:0] n158_I1; // @[Top.scala 194:22]
  wire [7:0] n158_O_0; // @[Top.scala 194:22]
  wire [7:0] n158_O_1; // @[Top.scala 194:22]
  wire  n165_valid_up; // @[Top.scala 198:22]
  wire  n165_valid_down; // @[Top.scala 198:22]
  wire [7:0] n165_I_0; // @[Top.scala 198:22]
  wire [7:0] n165_I_1; // @[Top.scala 198:22]
  wire [7:0] n165_O_0_0; // @[Top.scala 198:22]
  wire [7:0] n165_O_0_1; // @[Top.scala 198:22]
  wire  n170_clock; // @[Top.scala 201:22]
  wire  n170_reset; // @[Top.scala 201:22]
  wire  n170_valid_up; // @[Top.scala 201:22]
  wire  n170_valid_down; // @[Top.scala 201:22]
  wire [7:0] n170_I_0_0; // @[Top.scala 201:22]
  wire [7:0] n170_I_0_1; // @[Top.scala 201:22]
  wire [7:0] n170_O_0; // @[Top.scala 201:22]
  wire  n171_valid_up; // @[Top.scala 204:22]
  wire  n171_valid_down; // @[Top.scala 204:22]
  wire [7:0] n171_I0_0; // @[Top.scala 204:22]
  wire [7:0] n171_I1_0; // @[Top.scala 204:22]
  wire [7:0] n171_O_0_0; // @[Top.scala 204:22]
  wire [7:0] n171_O_0_1; // @[Top.scala 204:22]
  wire  n178_valid_up; // @[Top.scala 208:22]
  wire  n178_valid_down; // @[Top.scala 208:22]
  wire [7:0] n178_I_0_0; // @[Top.scala 208:22]
  wire [7:0] n178_I_0_1; // @[Top.scala 208:22]
  wire [7:0] n178_O_0_0; // @[Top.scala 208:22]
  wire [7:0] n178_O_0_1; // @[Top.scala 208:22]
  wire  n181_valid_up; // @[Top.scala 211:22]
  wire  n181_valid_down; // @[Top.scala 211:22]
  wire [7:0] n181_I_0_0; // @[Top.scala 211:22]
  wire [7:0] n181_I_0_1; // @[Top.scala 211:22]
  wire [7:0] n181_O_0; // @[Top.scala 211:22]
  wire [7:0] n181_O_1; // @[Top.scala 211:22]
  wire  n234_clock; // @[Top.scala 214:22]
  wire  n234_reset; // @[Top.scala 214:22]
  wire  n234_valid_up; // @[Top.scala 214:22]
  wire  n234_valid_down; // @[Top.scala 214:22]
  wire [7:0] n234_I_0; // @[Top.scala 214:22]
  wire [7:0] n234_I_1; // @[Top.scala 214:22]
  wire [7:0] n234_O; // @[Top.scala 214:22]
  wire  n235_valid_up; // @[Top.scala 217:22]
  wire  n235_valid_down; // @[Top.scala 217:22]
  wire [7:0] n235_I; // @[Top.scala 217:22]
  wire [7:0] n235_O; // @[Top.scala 217:22]
  wire  n236_clock; // @[Top.scala 220:22]
  wire  n236_reset; // @[Top.scala 220:22]
  wire  n236_valid_up; // @[Top.scala 220:22]
  wire  n236_valid_down; // @[Top.scala 220:22]
  wire [7:0] n236_I; // @[Top.scala 220:22]
  wire [7:0] n236_O; // @[Top.scala 220:22]
  wire  n237_clock; // @[Top.scala 223:22]
  wire  n237_reset; // @[Top.scala 223:22]
  wire  n237_valid_up; // @[Top.scala 223:22]
  wire  n237_valid_down; // @[Top.scala 223:22]
  wire [7:0] n237_I; // @[Top.scala 223:22]
  wire [7:0] n237_O; // @[Top.scala 223:22]
  wire  n238_clock; // @[Top.scala 226:22]
  wire  n238_reset; // @[Top.scala 226:22]
  wire  n238_valid_up; // @[Top.scala 226:22]
  wire  n238_valid_down; // @[Top.scala 226:22]
  wire [7:0] n238_I; // @[Top.scala 226:22]
  wire [7:0] n238_O; // @[Top.scala 226:22]
  FIFO n1 ( // @[Top.scala 86:20]
    .clock(n1_clock),
    .reset(n1_reset),
    .valid_up(n1_valid_up),
    .valid_down(n1_valid_down),
    .I(n1_I),
    .O(n1_O)
  );
  ShiftTN n2 ( // @[Top.scala 89:20]
    .clock(n2_clock),
    .reset(n2_reset),
    .valid_up(n2_valid_up),
    .valid_down(n2_valid_down),
    .I(n2_I),
    .O(n2_O)
  );
  ShiftTN n3 ( // @[Top.scala 92:20]
    .clock(n3_clock),
    .reset(n3_reset),
    .valid_up(n3_valid_up),
    .valid_down(n3_valid_down),
    .I(n3_I),
    .O(n3_O)
  );
  ShiftTN_2 n4 ( // @[Top.scala 95:20]
    .clock(n4_clock),
    .reset(n4_reset),
    .valid_up(n4_valid_up),
    .valid_down(n4_valid_down),
    .I(n4_I),
    .O(n4_O)
  );
  ShiftTN_2 n5 ( // @[Top.scala 98:20]
    .clock(n5_clock),
    .reset(n5_reset),
    .valid_up(n5_valid_up),
    .valid_down(n5_valid_down),
    .I(n5_I),
    .O(n5_O)
  );
  Map2T_1 n6 ( // @[Top.scala 101:20]
    .valid_up(n6_valid_up),
    .valid_down(n6_valid_down),
    .I0(n6_I0),
    .I1(n6_I1),
    .O_0(n6_O_0),
    .O_1(n6_O_1)
  );
  Map2T_3 n13 ( // @[Top.scala 105:21]
    .valid_up(n13_valid_up),
    .valid_down(n13_valid_down),
    .I0_0(n13_I0_0),
    .I0_1(n13_I0_1),
    .I1(n13_I1),
    .O_0(n13_O_0),
    .O_1(n13_O_1),
    .O_2(n13_O_2)
  );
  Passthrough n20 ( // @[Top.scala 109:21]
    .valid_up(n20_valid_up),
    .valid_down(n20_valid_down),
    .I_0(n20_I_0),
    .I_1(n20_I_1),
    .I_2(n20_I_2),
    .O_0_0(n20_O_0_0),
    .O_0_1(n20_O_0_1),
    .O_0_2(n20_O_0_2)
  );
  MapT n25 ( // @[Top.scala 112:21]
    .clock(n25_clock),
    .reset(n25_reset),
    .valid_up(n25_valid_up),
    .valid_down(n25_valid_down),
    .I_0_0(n25_I_0_0),
    .I_0_1(n25_I_0_1),
    .I_0_2(n25_I_0_2),
    .O_0(n25_O_0)
  );
  ShiftTN_2 n26 ( // @[Top.scala 115:21]
    .clock(n26_clock),
    .reset(n26_reset),
    .valid_up(n26_valid_up),
    .valid_down(n26_valid_down),
    .I(n26_I),
    .O(n26_O)
  );
  ShiftTN_2 n27 ( // @[Top.scala 118:21]
    .clock(n27_clock),
    .reset(n27_reset),
    .valid_up(n27_valid_up),
    .valid_down(n27_valid_down),
    .I(n27_I),
    .O(n27_O)
  );
  Map2T_1 n28 ( // @[Top.scala 121:21]
    .valid_up(n28_valid_up),
    .valid_down(n28_valid_down),
    .I0(n28_I0),
    .I1(n28_I1),
    .O_0(n28_O_0),
    .O_1(n28_O_1)
  );
  Map2T_3 n35 ( // @[Top.scala 125:21]
    .valid_up(n35_valid_up),
    .valid_down(n35_valid_down),
    .I0_0(n35_I0_0),
    .I0_1(n35_I0_1),
    .I1(n35_I1),
    .O_0(n35_O_0),
    .O_1(n35_O_1),
    .O_2(n35_O_2)
  );
  Passthrough n42 ( // @[Top.scala 129:21]
    .valid_up(n42_valid_up),
    .valid_down(n42_valid_down),
    .I_0(n42_I_0),
    .I_1(n42_I_1),
    .I_2(n42_I_2),
    .O_0_0(n42_O_0_0),
    .O_0_1(n42_O_0_1),
    .O_0_2(n42_O_0_2)
  );
  MapT n47 ( // @[Top.scala 132:21]
    .clock(n47_clock),
    .reset(n47_reset),
    .valid_up(n47_valid_up),
    .valid_down(n47_valid_down),
    .I_0_0(n47_I_0_0),
    .I_0_1(n47_I_0_1),
    .I_0_2(n47_I_0_2),
    .O_0(n47_O_0)
  );
  Map2T_8 n48 ( // @[Top.scala 135:21]
    .valid_up(n48_valid_up),
    .valid_down(n48_valid_down),
    .I0_0(n48_I0_0),
    .I1_0(n48_I1_0),
    .O_0_0(n48_O_0_0),
    .O_0_1(n48_O_0_1)
  );
  ShiftTN_2 n55 ( // @[Top.scala 139:21]
    .clock(n55_clock),
    .reset(n55_reset),
    .valid_up(n55_valid_up),
    .valid_down(n55_valid_down),
    .I(n55_I),
    .O(n55_O)
  );
  ShiftTN_2 n56 ( // @[Top.scala 142:21]
    .clock(n56_clock),
    .reset(n56_reset),
    .valid_up(n56_valid_up),
    .valid_down(n56_valid_down),
    .I(n56_I),
    .O(n56_O)
  );
  Map2T_1 n57 ( // @[Top.scala 145:21]
    .valid_up(n57_valid_up),
    .valid_down(n57_valid_down),
    .I0(n57_I0),
    .I1(n57_I1),
    .O_0(n57_O_0),
    .O_1(n57_O_1)
  );
  Map2T_3 n64 ( // @[Top.scala 149:21]
    .valid_up(n64_valid_up),
    .valid_down(n64_valid_down),
    .I0_0(n64_I0_0),
    .I0_1(n64_I0_1),
    .I1(n64_I1),
    .O_0(n64_O_0),
    .O_1(n64_O_1),
    .O_2(n64_O_2)
  );
  Passthrough n71 ( // @[Top.scala 153:21]
    .valid_up(n71_valid_up),
    .valid_down(n71_valid_down),
    .I_0(n71_I_0),
    .I_1(n71_I_1),
    .I_2(n71_I_2),
    .O_0_0(n71_O_0_0),
    .O_0_1(n71_O_0_1),
    .O_0_2(n71_O_0_2)
  );
  MapT n76 ( // @[Top.scala 156:21]
    .clock(n76_clock),
    .reset(n76_reset),
    .valid_up(n76_valid_up),
    .valid_down(n76_valid_down),
    .I_0_0(n76_I_0_0),
    .I_0_1(n76_I_0_1),
    .I_0_2(n76_I_0_2),
    .O_0(n76_O_0)
  );
  Map2T_13 n77 ( // @[Top.scala 159:21]
    .valid_up(n77_valid_up),
    .valid_down(n77_valid_down),
    .I0_0_0(n77_I0_0_0),
    .I0_0_1(n77_I0_0_1),
    .I1_0(n77_I1_0),
    .O_0_0(n77_O_0_0),
    .O_0_1(n77_O_0_1),
    .O_0_2(n77_O_0_2)
  );
  Passthrough_3 n84 ( // @[Top.scala 163:21]
    .valid_up(n84_valid_up),
    .valid_down(n84_valid_down),
    .I_0_0(n84_I_0_0),
    .I_0_1(n84_I_0_1),
    .I_0_2(n84_I_0_2),
    .O_0_0(n84_O_0_0),
    .O_0_1(n84_O_0_1),
    .O_0_2(n84_O_0_2)
  );
  MapT_3 n87 ( // @[Top.scala 166:21]
    .valid_up(n87_valid_up),
    .valid_down(n87_valid_down),
    .I_0_0(n87_I_0_0),
    .I_0_1(n87_I_0_1),
    .I_0_2(n87_I_0_2),
    .O_0(n87_O_0),
    .O_1(n87_O_1),
    .O_2(n87_O_2)
  );
  MapT_10 n140 ( // @[Top.scala 169:22]
    .clock(n140_clock),
    .reset(n140_reset),
    .valid_up(n140_valid_up),
    .valid_down(n140_valid_down),
    .I_0(n140_I_0),
    .I_1(n140_I_1),
    .I_2(n140_I_2),
    .O(n140_O)
  );
  Passthrough_6 n141 ( // @[Top.scala 172:22]
    .valid_up(n141_valid_up),
    .valid_down(n141_valid_down),
    .I(n141_I),
    .O(n141_O)
  );
  ShiftTN n142 ( // @[Top.scala 175:22]
    .clock(n142_clock),
    .reset(n142_reset),
    .valid_up(n142_valid_up),
    .valid_down(n142_valid_down),
    .I(n142_I),
    .O(n142_O)
  );
  ShiftTN_2 n143 ( // @[Top.scala 178:22]
    .clock(n143_clock),
    .reset(n143_reset),
    .valid_up(n143_valid_up),
    .valid_down(n143_valid_down),
    .I(n143_I),
    .O(n143_O)
  );
  Map2T_1 n144 ( // @[Top.scala 181:22]
    .valid_up(n144_valid_up),
    .valid_down(n144_valid_down),
    .I0(n144_I0),
    .I1(n144_I1),
    .O_0(n144_O_0),
    .O_1(n144_O_1)
  );
  Passthrough_7 n151 ( // @[Top.scala 185:22]
    .valid_up(n151_valid_up),
    .valid_down(n151_valid_down),
    .I_0(n151_I_0),
    .I_1(n151_I_1),
    .O_0_0(n151_O_0_0),
    .O_0_1(n151_O_0_1)
  );
  MapT_11 n156 ( // @[Top.scala 188:22]
    .clock(n156_clock),
    .reset(n156_reset),
    .valid_up(n156_valid_up),
    .valid_down(n156_valid_down),
    .I_0_0(n156_I_0_0),
    .I_0_1(n156_I_0_1),
    .O_0(n156_O_0)
  );
  ShiftTN_2 n157 ( // @[Top.scala 191:22]
    .clock(n157_clock),
    .reset(n157_reset),
    .valid_up(n157_valid_up),
    .valid_down(n157_valid_down),
    .I(n157_I),
    .O(n157_O)
  );
  Map2T_1 n158 ( // @[Top.scala 194:22]
    .valid_up(n158_valid_up),
    .valid_down(n158_valid_down),
    .I0(n158_I0),
    .I1(n158_I1),
    .O_0(n158_O_0),
    .O_1(n158_O_1)
  );
  Passthrough_7 n165 ( // @[Top.scala 198:22]
    .valid_up(n165_valid_up),
    .valid_down(n165_valid_down),
    .I_0(n165_I_0),
    .I_1(n165_I_1),
    .O_0_0(n165_O_0_0),
    .O_0_1(n165_O_0_1)
  );
  MapT_11 n170 ( // @[Top.scala 201:22]
    .clock(n170_clock),
    .reset(n170_reset),
    .valid_up(n170_valid_up),
    .valid_down(n170_valid_down),
    .I_0_0(n170_I_0_0),
    .I_0_1(n170_I_0_1),
    .O_0(n170_O_0)
  );
  Map2T_8 n171 ( // @[Top.scala 204:22]
    .valid_up(n171_valid_up),
    .valid_down(n171_valid_down),
    .I0_0(n171_I0_0),
    .I1_0(n171_I1_0),
    .O_0_0(n171_O_0_0),
    .O_0_1(n171_O_0_1)
  );
  Passthrough_9 n178 ( // @[Top.scala 208:22]
    .valid_up(n178_valid_up),
    .valid_down(n178_valid_down),
    .I_0_0(n178_I_0_0),
    .I_0_1(n178_I_0_1),
    .O_0_0(n178_O_0_0),
    .O_0_1(n178_O_0_1)
  );
  MapT_13 n181 ( // @[Top.scala 211:22]
    .valid_up(n181_valid_up),
    .valid_down(n181_valid_down),
    .I_0_0(n181_I_0_0),
    .I_0_1(n181_I_0_1),
    .O_0(n181_O_0),
    .O_1(n181_O_1)
  );
  MapT_20 n234 ( // @[Top.scala 214:22]
    .clock(n234_clock),
    .reset(n234_reset),
    .valid_up(n234_valid_up),
    .valid_down(n234_valid_down),
    .I_0(n234_I_0),
    .I_1(n234_I_1),
    .O(n234_O)
  );
  Passthrough_6 n235 ( // @[Top.scala 217:22]
    .valid_up(n235_valid_up),
    .valid_down(n235_valid_down),
    .I(n235_I),
    .O(n235_O)
  );
  FIFO n236 ( // @[Top.scala 220:22]
    .clock(n236_clock),
    .reset(n236_reset),
    .valid_up(n236_valid_up),
    .valid_down(n236_valid_down),
    .I(n236_I),
    .O(n236_O)
  );
  FIFO n237 ( // @[Top.scala 223:22]
    .clock(n237_clock),
    .reset(n237_reset),
    .valid_up(n237_valid_up),
    .valid_down(n237_valid_down),
    .I(n237_I),
    .O(n237_O)
  );
  FIFO n238 ( // @[Top.scala 226:22]
    .clock(n238_clock),
    .reset(n238_reset),
    .valid_up(n238_valid_up),
    .valid_down(n238_valid_down),
    .I(n238_I),
    .O(n238_O)
  );
  assign valid_down = n238_valid_down; // @[Top.scala 230:16]
  assign O = n238_O; // @[Top.scala 229:7]
  assign n1_clock = clock;
  assign n1_reset = reset;
  assign n1_valid_up = valid_up; // @[Top.scala 88:17]
  assign n1_I = I; // @[Top.scala 87:10]
  assign n2_clock = clock;
  assign n2_reset = reset;
  assign n2_valid_up = n1_valid_down; // @[Top.scala 91:17]
  assign n2_I = n1_O; // @[Top.scala 90:10]
  assign n3_clock = clock;
  assign n3_reset = reset;
  assign n3_valid_up = n2_valid_down; // @[Top.scala 94:17]
  assign n3_I = n2_O; // @[Top.scala 93:10]
  assign n4_clock = clock;
  assign n4_reset = reset;
  assign n4_valid_up = n3_valid_down; // @[Top.scala 97:17]
  assign n4_I = n3_O; // @[Top.scala 96:10]
  assign n5_clock = clock;
  assign n5_reset = reset;
  assign n5_valid_up = n4_valid_down; // @[Top.scala 100:17]
  assign n5_I = n4_O; // @[Top.scala 99:10]
  assign n6_valid_up = n5_valid_down & n4_valid_down; // @[Top.scala 104:17]
  assign n6_I0 = n5_O; // @[Top.scala 102:11]
  assign n6_I1 = n4_O; // @[Top.scala 103:11]
  assign n13_valid_up = n6_valid_down & n3_valid_down; // @[Top.scala 108:18]
  assign n13_I0_0 = n6_O_0; // @[Top.scala 106:12]
  assign n13_I0_1 = n6_O_1; // @[Top.scala 106:12]
  assign n13_I1 = n3_O; // @[Top.scala 107:12]
  assign n20_valid_up = n13_valid_down; // @[Top.scala 111:18]
  assign n20_I_0 = n13_O_0; // @[Top.scala 110:11]
  assign n20_I_1 = n13_O_1; // @[Top.scala 110:11]
  assign n20_I_2 = n13_O_2; // @[Top.scala 110:11]
  assign n25_clock = clock;
  assign n25_reset = reset;
  assign n25_valid_up = n20_valid_down; // @[Top.scala 114:18]
  assign n25_I_0_0 = n20_O_0_0; // @[Top.scala 113:11]
  assign n25_I_0_1 = n20_O_0_1; // @[Top.scala 113:11]
  assign n25_I_0_2 = n20_O_0_2; // @[Top.scala 113:11]
  assign n26_clock = clock;
  assign n26_reset = reset;
  assign n26_valid_up = n2_valid_down; // @[Top.scala 117:18]
  assign n26_I = n2_O; // @[Top.scala 116:11]
  assign n27_clock = clock;
  assign n27_reset = reset;
  assign n27_valid_up = n26_valid_down; // @[Top.scala 120:18]
  assign n27_I = n26_O; // @[Top.scala 119:11]
  assign n28_valid_up = n27_valid_down & n26_valid_down; // @[Top.scala 124:18]
  assign n28_I0 = n27_O; // @[Top.scala 122:12]
  assign n28_I1 = n26_O; // @[Top.scala 123:12]
  assign n35_valid_up = n28_valid_down & n2_valid_down; // @[Top.scala 128:18]
  assign n35_I0_0 = n28_O_0; // @[Top.scala 126:12]
  assign n35_I0_1 = n28_O_1; // @[Top.scala 126:12]
  assign n35_I1 = n2_O; // @[Top.scala 127:12]
  assign n42_valid_up = n35_valid_down; // @[Top.scala 131:18]
  assign n42_I_0 = n35_O_0; // @[Top.scala 130:11]
  assign n42_I_1 = n35_O_1; // @[Top.scala 130:11]
  assign n42_I_2 = n35_O_2; // @[Top.scala 130:11]
  assign n47_clock = clock;
  assign n47_reset = reset;
  assign n47_valid_up = n42_valid_down; // @[Top.scala 134:18]
  assign n47_I_0_0 = n42_O_0_0; // @[Top.scala 133:11]
  assign n47_I_0_1 = n42_O_0_1; // @[Top.scala 133:11]
  assign n47_I_0_2 = n42_O_0_2; // @[Top.scala 133:11]
  assign n48_valid_up = n25_valid_down & n47_valid_down; // @[Top.scala 138:18]
  assign n48_I0_0 = n25_O_0; // @[Top.scala 136:12]
  assign n48_I1_0 = n47_O_0; // @[Top.scala 137:12]
  assign n55_clock = clock;
  assign n55_reset = reset;
  assign n55_valid_up = n1_valid_down; // @[Top.scala 141:18]
  assign n55_I = n1_O; // @[Top.scala 140:11]
  assign n56_clock = clock;
  assign n56_reset = reset;
  assign n56_valid_up = n55_valid_down; // @[Top.scala 144:18]
  assign n56_I = n55_O; // @[Top.scala 143:11]
  assign n57_valid_up = n56_valid_down & n55_valid_down; // @[Top.scala 148:18]
  assign n57_I0 = n56_O; // @[Top.scala 146:12]
  assign n57_I1 = n55_O; // @[Top.scala 147:12]
  assign n64_valid_up = n57_valid_down & n1_valid_down; // @[Top.scala 152:18]
  assign n64_I0_0 = n57_O_0; // @[Top.scala 150:12]
  assign n64_I0_1 = n57_O_1; // @[Top.scala 150:12]
  assign n64_I1 = n1_O; // @[Top.scala 151:12]
  assign n71_valid_up = n64_valid_down; // @[Top.scala 155:18]
  assign n71_I_0 = n64_O_0; // @[Top.scala 154:11]
  assign n71_I_1 = n64_O_1; // @[Top.scala 154:11]
  assign n71_I_2 = n64_O_2; // @[Top.scala 154:11]
  assign n76_clock = clock;
  assign n76_reset = reset;
  assign n76_valid_up = n71_valid_down; // @[Top.scala 158:18]
  assign n76_I_0_0 = n71_O_0_0; // @[Top.scala 157:11]
  assign n76_I_0_1 = n71_O_0_1; // @[Top.scala 157:11]
  assign n76_I_0_2 = n71_O_0_2; // @[Top.scala 157:11]
  assign n77_valid_up = n48_valid_down & n76_valid_down; // @[Top.scala 162:18]
  assign n77_I0_0_0 = n48_O_0_0; // @[Top.scala 160:12]
  assign n77_I0_0_1 = n48_O_0_1; // @[Top.scala 160:12]
  assign n77_I1_0 = n76_O_0; // @[Top.scala 161:12]
  assign n84_valid_up = n77_valid_down; // @[Top.scala 165:18]
  assign n84_I_0_0 = n77_O_0_0; // @[Top.scala 164:11]
  assign n84_I_0_1 = n77_O_0_1; // @[Top.scala 164:11]
  assign n84_I_0_2 = n77_O_0_2; // @[Top.scala 164:11]
  assign n87_valid_up = n84_valid_down; // @[Top.scala 168:18]
  assign n87_I_0_0 = n84_O_0_0; // @[Top.scala 167:11]
  assign n87_I_0_1 = n84_O_0_1; // @[Top.scala 167:11]
  assign n87_I_0_2 = n84_O_0_2; // @[Top.scala 167:11]
  assign n140_clock = clock;
  assign n140_reset = reset;
  assign n140_valid_up = n87_valid_down; // @[Top.scala 171:19]
  assign n140_I_0 = n87_O_0; // @[Top.scala 170:12]
  assign n140_I_1 = n87_O_1; // @[Top.scala 170:12]
  assign n140_I_2 = n87_O_2; // @[Top.scala 170:12]
  assign n141_valid_up = n140_valid_down; // @[Top.scala 174:19]
  assign n141_I = n140_O; // @[Top.scala 173:12]
  assign n142_clock = clock;
  assign n142_reset = reset;
  assign n142_valid_up = n141_valid_down; // @[Top.scala 177:19]
  assign n142_I = n141_O; // @[Top.scala 176:12]
  assign n143_clock = clock;
  assign n143_reset = reset;
  assign n143_valid_up = n142_valid_down; // @[Top.scala 180:19]
  assign n143_I = n142_O; // @[Top.scala 179:12]
  assign n144_valid_up = n143_valid_down & n142_valid_down; // @[Top.scala 184:19]
  assign n144_I0 = n143_O; // @[Top.scala 182:13]
  assign n144_I1 = n142_O; // @[Top.scala 183:13]
  assign n151_valid_up = n144_valid_down; // @[Top.scala 187:19]
  assign n151_I_0 = n144_O_0; // @[Top.scala 186:12]
  assign n151_I_1 = n144_O_1; // @[Top.scala 186:12]
  assign n156_clock = clock;
  assign n156_reset = reset;
  assign n156_valid_up = n151_valid_down; // @[Top.scala 190:19]
  assign n156_I_0_0 = n151_O_0_0; // @[Top.scala 189:12]
  assign n156_I_0_1 = n151_O_0_1; // @[Top.scala 189:12]
  assign n157_clock = clock;
  assign n157_reset = reset;
  assign n157_valid_up = n141_valid_down; // @[Top.scala 193:19]
  assign n157_I = n141_O; // @[Top.scala 192:12]
  assign n158_valid_up = n157_valid_down & n141_valid_down; // @[Top.scala 197:19]
  assign n158_I0 = n157_O; // @[Top.scala 195:13]
  assign n158_I1 = n141_O; // @[Top.scala 196:13]
  assign n165_valid_up = n158_valid_down; // @[Top.scala 200:19]
  assign n165_I_0 = n158_O_0; // @[Top.scala 199:12]
  assign n165_I_1 = n158_O_1; // @[Top.scala 199:12]
  assign n170_clock = clock;
  assign n170_reset = reset;
  assign n170_valid_up = n165_valid_down; // @[Top.scala 203:19]
  assign n170_I_0_0 = n165_O_0_0; // @[Top.scala 202:12]
  assign n170_I_0_1 = n165_O_0_1; // @[Top.scala 202:12]
  assign n171_valid_up = n156_valid_down & n170_valid_down; // @[Top.scala 207:19]
  assign n171_I0_0 = n156_O_0; // @[Top.scala 205:13]
  assign n171_I1_0 = n170_O_0; // @[Top.scala 206:13]
  assign n178_valid_up = n171_valid_down; // @[Top.scala 210:19]
  assign n178_I_0_0 = n171_O_0_0; // @[Top.scala 209:12]
  assign n178_I_0_1 = n171_O_0_1; // @[Top.scala 209:12]
  assign n181_valid_up = n178_valid_down; // @[Top.scala 213:19]
  assign n181_I_0_0 = n178_O_0_0; // @[Top.scala 212:12]
  assign n181_I_0_1 = n178_O_0_1; // @[Top.scala 212:12]
  assign n234_clock = clock;
  assign n234_reset = reset;
  assign n234_valid_up = n181_valid_down; // @[Top.scala 216:19]
  assign n234_I_0 = n181_O_0; // @[Top.scala 215:12]
  assign n234_I_1 = n181_O_1; // @[Top.scala 215:12]
  assign n235_valid_up = n234_valid_down; // @[Top.scala 219:19]
  assign n235_I = n234_O; // @[Top.scala 218:12]
  assign n236_clock = clock;
  assign n236_reset = reset;
  assign n236_valid_up = n235_valid_down; // @[Top.scala 222:19]
  assign n236_I = n235_O; // @[Top.scala 221:12]
  assign n237_clock = clock;
  assign n237_reset = reset;
  assign n237_valid_up = n236_valid_down; // @[Top.scala 225:19]
  assign n237_I = n236_O; // @[Top.scala 224:12]
  assign n238_clock = clock;
  assign n238_reset = reset;
  assign n238_valid_up = n237_valid_down; // @[Top.scala 228:19]
  assign n238_I = n237_O; // @[Top.scala 227:12]
endmodule
