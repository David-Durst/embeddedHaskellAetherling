module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [31:0] I_0,
  output [31:0] O_0
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset(reset), // @[:@1297.4]
    .io_in_x209_TREADY(dontcare), // @[:@1298.4]
    .io_in_x209_TDATA(I_0), // @[:@1298.4]
    .io_in_x209_TID(8'h0),
    .io_in_x209_TDEST(8'h0),
    .io_in_x210_TVALID(valid_down), // @[:@1298.4]
    .io_in_x210_TDATA(O_0), // @[:@1298.4]
    .io_in_x210_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x217_ctrchain cchain ( // @[:@2879.2]
    .clock(CLK), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule


module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule



module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 325:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh49); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh49); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [31:0] io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@512.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@512.4]
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@512.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign io_rdata = SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@539.4]
  assign SRAMVerilogAWS_wdata = 32'h0; // @[SRAM.scala 175:20:@526.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@527.4]
  assign SRAMVerilogAWS_wen = 1'h0; // @[SRAM.scala 173:18:@524.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@529.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@528.4]
  assign SRAMVerilogAWS_waddr = 21'h0; // @[SRAM.scala 174:20:@525.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@523.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@553.2]
  input         clock, // @[:@554.4]
  input         reset, // @[:@555.4]
  input         io_flow, // @[:@556.4]
  input  [20:0] io_in, // @[:@556.4]
  output [20:0] io_out // @[:@556.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@558.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@558.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@571.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@570.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@569.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@568.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@567.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@565.4]
endmodule
module Mem1D( // @[:@573.2]
  input         clock, // @[:@574.4]
  input         reset, // @[:@575.4]
  input  [20:0] io_r_ofs_0, // @[:@576.4]
  input         io_r_backpressure, // @[:@576.4]
  output [31:0] io_output // @[:@576.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@580.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@580.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@580.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@580.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@583.4]
  SRAM SRAM ( // @[MemPrimitives.scala 715:21:@580.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@583.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@596.4]
  assign SRAM_clock = clock; // @[:@581.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@590.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@595.4]
  assign RetimeWrapper_clock = clock; // @[:@584.4]
  assign RetimeWrapper_reset = reset; // @[:@585.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@587.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@586.4]
endmodule
module StickySelects( // @[:@598.2]
  input   io_ins_0, // @[:@601.4]
  output  io_outs_0 // @[:@601.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@603.4]
endmodule
module RetimeWrapper_6( // @[:@617.2]
  input   clock, // @[:@618.4]
  input   reset, // @[:@619.4]
  input   io_flow, // @[:@620.4]
  input   io_in, // @[:@620.4]
  output  io_out // @[:@620.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@622.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@622.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@635.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@634.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@633.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@632.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@631.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@629.4]
endmodule
module x211_outbuf_0( // @[:@637.2]
  input         clock, // @[:@638.4]
  input         reset, // @[:@639.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@640.4]
  input         io_rPort_0_en_0, // @[:@640.4]
  input         io_rPort_0_backpressure, // @[:@640.4]
  output [31:0] io_rPort_0_output_0 // @[:@640.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@655.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@655.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@655.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@695.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@685.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@687.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@655.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@681.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@695.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@685.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@687.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@702.4]
  assign Mem1D_clock = clock; // @[:@656.4]
  assign Mem1D_reset = reset; // @[:@657.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 131:28:@691.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 132:32:@692.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@684.4]
  assign RetimeWrapper_clock = clock; // @[:@696.4]
  assign RetimeWrapper_reset = reset; // @[:@697.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@699.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@698.4]
endmodule
module x493_sm( // @[:@846.2]
  input   clock, // @[:@847.4]
  input   reset, // @[:@848.4]
  input   io_enable, // @[:@849.4]
  output  io_done, // @[:@849.4]
  input   io_ctrDone, // @[:@849.4]
  output  io_ctrInc, // @[:@849.4]
  input   io_parentAck, // @[:@849.4]
  input   io_doneIn_0, // @[:@849.4]
  input   io_doneIn_1, // @[:@849.4]
  output  io_enableOut_0, // @[:@849.4]
  output  io_enableOut_1, // @[:@849.4]
  output  io_childAck_0, // @[:@849.4]
  output  io_childAck_1 // @[:@849.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@852.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@855.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@858.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@861.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@893.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1011.4]
  wire  allDone; // @[Controllers.scala 80:47:@864.4]
  wire  synchronize; // @[Controllers.scala 146:56:@918.4]
  wire  _T_127; // @[Controllers.scala 150:35:@920.4]
  wire  _T_129; // @[Controllers.scala 150:60:@921.4]
  wire  _T_130; // @[Controllers.scala 150:58:@922.4]
  wire  _T_132; // @[Controllers.scala 150:76:@923.4]
  wire  _T_133; // @[Controllers.scala 150:74:@924.4]
  wire  _T_135; // @[Controllers.scala 150:97:@925.4]
  wire  _T_136; // @[Controllers.scala 150:95:@926.4]
  wire  _T_152; // @[Controllers.scala 150:35:@944.4]
  wire  _T_154; // @[Controllers.scala 150:60:@945.4]
  wire  _T_155; // @[Controllers.scala 150:58:@946.4]
  wire  _T_157; // @[Controllers.scala 150:76:@947.4]
  wire  _T_158; // @[Controllers.scala 150:74:@948.4]
  wire  _T_161; // @[Controllers.scala 150:95:@950.4]
  wire  _T_179; // @[Controllers.scala 213:68:@972.4]
  wire  _T_181; // @[Controllers.scala 213:90:@974.4]
  wire  _T_183; // @[Controllers.scala 213:132:@976.4]
  wire  _T_184; // @[Controllers.scala 213:130:@977.4]
  wire  _T_185; // @[Controllers.scala 213:156:@978.4]
  wire  _T_187; // @[Controllers.scala 213:68:@981.4]
  wire  _T_189; // @[Controllers.scala 213:90:@983.4]
  wire  _T_196; // @[package.scala 100:49:@989.4]
  reg  _T_199; // @[package.scala 48:56:@990.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@992.4]
  reg  _T_213; // @[package.scala 48:56:@1008.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@852.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@855.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@858.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@861.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@890.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@893.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@994.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1011.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@864.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@918.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@920.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@921.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@922.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@923.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@924.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@925.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@926.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@944.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@945.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@946.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@947.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@948.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@950.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@972.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@974.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@976.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@977.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@978.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@981.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@983.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@989.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@992.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1018.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@917.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@980.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@988.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@969.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@971.4]
  assign active_0_clock = clock; // @[:@853.4]
  assign active_0_reset = reset; // @[:@854.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@929.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@933.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@867.4]
  assign active_1_clock = clock; // @[:@856.4]
  assign active_1_reset = reset; // @[:@857.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@953.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@957.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@868.4]
  assign done_0_clock = clock; // @[:@859.4]
  assign done_0_reset = reset; // @[:@860.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@943.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@879.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@869.4]
  assign done_1_clock = clock; // @[:@862.4]
  assign done_1_reset = reset; // @[:@863.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@967.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@888.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@870.4]
  assign iterDone_0_clock = clock; // @[:@891.4]
  assign iterDone_0_reset = reset; // @[:@892.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@939.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@906.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@896.4]
  assign iterDone_1_clock = clock; // @[:@894.4]
  assign iterDone_1_reset = reset; // @[:@895.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@963.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@915.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@897.4]
  assign RetimeWrapper_clock = clock; // @[:@995.4]
  assign RetimeWrapper_reset = reset; // @[:@996.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@998.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@997.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1012.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1013.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1015.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1014.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x361_outr_UnitPipe_sm( // @[:@1435.2]
  input   clock, // @[:@1436.4]
  input   reset, // @[:@1437.4]
  input   io_enable, // @[:@1438.4]
  output  io_done, // @[:@1438.4]
  input   io_parentAck, // @[:@1438.4]
  input   io_doneIn_0, // @[:@1438.4]
  input   io_doneIn_1, // @[:@1438.4]
  output  io_enableOut_0, // @[:@1438.4]
  output  io_enableOut_1, // @[:@1438.4]
  output  io_childAck_0, // @[:@1438.4]
  output  io_childAck_1, // @[:@1438.4]
  input   io_ctrCopyDone_0, // @[:@1438.4]
  input   io_ctrCopyDone_1 // @[:@1438.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1441.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1444.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1447.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1450.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1482.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1688.4]
  wire  allDone; // @[Controllers.scala 80:47:@1453.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1507.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1508.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1509.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1510.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1511.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1514.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1516.4]
  wire  _T_148; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1531.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1532.4]
  wire  _T_160; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  wire  _T_178; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1563.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1564.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1576.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1577.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1578.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1579.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1580.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1583.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1585.4]
  wire  _T_216; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1600.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1601.4]
  wire  _T_228; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  wire  _T_246; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1632.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1633.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1649.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1651.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1653.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1658.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1660.4]
  wire  _T_282; // @[package.scala 100:49:@1666.4]
  reg  _T_285; // @[package.scala 48:56:@1667.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1669.4]
  reg  _T_299; // @[package.scala 48:56:@1685.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1441.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1444.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1447.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1450.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1479.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1482.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1523.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1537.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1555.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1592.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1606.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1624.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1671.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1688.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1453.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1507.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1508.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1509.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1510.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1511.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1514.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1516.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1531.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1532.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1563.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1564.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1576.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1577.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1578.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1579.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1580.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1583.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1585.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1600.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1601.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1632.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1633.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1649.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1651.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1653.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1658.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1660.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1666.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1669.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1695.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1657.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1665.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1646.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1648.4]
  assign active_0_clock = clock; // @[:@1442.4]
  assign active_0_reset = reset; // @[:@1443.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1518.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1522.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1456.4]
  assign active_1_clock = clock; // @[:@1445.4]
  assign active_1_reset = reset; // @[:@1446.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1587.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1591.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1457.4]
  assign done_0_clock = clock; // @[:@1448.4]
  assign done_0_reset = reset; // @[:@1449.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1568.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1468.4 Controllers.scala 170:32:@1575.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1458.4]
  assign done_1_clock = clock; // @[:@1451.4]
  assign done_1_reset = reset; // @[:@1452.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1637.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1477.4 Controllers.scala 170:32:@1644.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1459.4]
  assign iterDone_0_clock = clock; // @[:@1480.4]
  assign iterDone_0_reset = reset; // @[:@1481.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1536.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1495.4 Controllers.scala 168:36:@1552.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1485.4]
  assign iterDone_1_clock = clock; // @[:@1483.4]
  assign iterDone_1_reset = reset; // @[:@1484.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1605.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1504.4 Controllers.scala 168:36:@1621.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1486.4]
  assign RetimeWrapper_clock = clock; // @[:@1524.4]
  assign RetimeWrapper_reset = reset; // @[:@1525.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1527.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1526.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1538.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1539.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1541.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1540.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1556.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1557.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1559.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1558.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1593.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1594.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1596.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1595.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1607.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1608.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1610.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1609.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1625.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1626.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1628.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1627.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1672.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1673.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1675.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1674.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1689.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1690.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1692.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1691.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1924.2]
  input   clock, // @[:@1925.4]
  input   reset, // @[:@1926.4]
  input   io_input_inc_en_0, // @[:@1927.4]
  input   io_input_dinc_en_0, // @[:@1927.4]
  output  io_output_full // @[:@1927.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1929.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1930.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1931.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1932.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1932.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1933.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1934.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1935.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1935.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1936.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1937.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1930.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1931.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1932.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1932.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1933.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1934.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1935.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1935.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1936.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1937.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1951.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x212_fifoinraw_0( // @[:@2074.2]
  input   clock, // @[:@2075.4]
  input   reset // @[:@2076.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2121.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2121.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2122.4]
  assign elements_reset = reset; // @[:@2123.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 394:79:@2133.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2134.4]
endmodule
module x213_fifoinpacked_0( // @[:@2497.2]
  input   clock, // @[:@2498.4]
  input   reset, // @[:@2499.4]
  input   io_wPort_0_en_0, // @[:@2500.4]
  output  io_full, // @[:@2500.4]
  input   io_active_0_in, // @[:@2500.4]
  output  io_active_0_out // @[:@2500.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2544.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2544.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 439:39:@2618.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 437:129:@2616.4]
  assign elements_clock = clock; // @[:@2545.4]
  assign elements_reset = reset; // @[:@2546.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 394:79:@2556.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2557.4]
endmodule
module FF_7( // @[:@3047.2]
  input         clock, // @[:@3048.4]
  input         reset, // @[:@3049.4]
  output [12:0] io_rPort_0_output_0, // @[:@3050.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3050.4]
  input         io_wPort_0_reset, // @[:@3050.4]
  input         io_wPort_0_en_0 // @[:@3050.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 321:19:@3065.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 325:32:@3067.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 325:12:@3068.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@3067.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 325:12:@3068.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@3070.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3085.2]
  input         clock, // @[:@3086.4]
  input         reset, // @[:@3087.4]
  input         io_setup_saturate, // @[:@3088.4]
  input         io_input_reset, // @[:@3088.4]
  input         io_input_enable, // @[:@3088.4]
  output [12:0] io_output_count_0, // @[:@3088.4]
  output        io_output_oobs_0, // @[:@3088.4]
  output        io_output_done, // @[:@3088.4]
  output        io_output_saturated // @[:@3088.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3101.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3117.4]
  wire  _T_36; // @[Counter.scala 264:45:@3120.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3145.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3146.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3147.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3148.4]
  wire  _T_57; // @[Counter.scala 293:18:@3150.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3158.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3160.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3161.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3162.4]
  wire  _T_75; // @[Counter.scala 322:102:@3166.4]
  wire  _T_77; // @[Counter.scala 322:130:@3167.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3101.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3117.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3120.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3145.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3146.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3147.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3148.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3150.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3158.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3160.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3161.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3162.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3166.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3167.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3165.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3169.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3171.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3174.4]
  assign bases_0_clock = clock; // @[:@3102.4]
  assign bases_0_reset = reset; // @[:@3103.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3164.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3143.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3144.4]
  assign SRFF_clock = clock; // @[:@3118.4]
  assign SRFF_reset = reset; // @[:@3119.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3122.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3124.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3125.4]
endmodule
module SingleCounter_2( // @[:@3214.2]
  input         clock, // @[:@3215.4]
  input         reset, // @[:@3216.4]
  input         io_setup_saturate, // @[:@3217.4]
  input         io_input_reset, // @[:@3217.4]
  input         io_input_enable, // @[:@3217.4]
  output [12:0] io_output_count_0, // @[:@3217.4]
  output        io_output_oobs_0, // @[:@3217.4]
  output        io_output_done // @[:@3217.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3230.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3246.4]
  wire  _T_36; // @[Counter.scala 264:45:@3249.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3274.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3275.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3276.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3277.4]
  wire  _T_57; // @[Counter.scala 293:18:@3279.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3287.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3289.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3290.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3291.4]
  wire  _T_75; // @[Counter.scala 322:102:@3295.4]
  wire  _T_77; // @[Counter.scala 322:130:@3296.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3230.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3246.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3249.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3274.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3275.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3276.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3277.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3279.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3287.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3289.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3290.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3291.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3295.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3296.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3294.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3298.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3300.4]
  assign bases_0_clock = clock; // @[:@3231.4]
  assign bases_0_reset = reset; // @[:@3232.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3293.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3272.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3273.4]
  assign SRFF_clock = clock; // @[:@3247.4]
  assign SRFF_reset = reset; // @[:@3248.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3251.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3253.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3254.4]
endmodule
module x217_ctrchain( // @[:@3305.2]
  input         clock, // @[:@3306.4]
  input         reset, // @[:@3307.4]
  input         io_input_reset, // @[:@3308.4]
  input         io_input_enable, // @[:@3308.4]
  output [12:0] io_output_counts_1, // @[:@3308.4]
  output [12:0] io_output_counts_0, // @[:@3308.4]
  output        io_output_oobs_0, // @[:@3308.4]
  output        io_output_oobs_1, // @[:@3308.4]
  output        io_output_done // @[:@3308.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3310.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3313.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3313.4]
  wire  isDone; // @[Counter.scala 541:51:@3330.4]
  reg  wasDone; // @[Counter.scala 542:24:@3331.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3339.4]
  wire  _T_66; // @[Counter.scala 546:80:@3340.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3345.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3346.4]
  wire  _T_74; // @[Counter.scala 551:19:@3347.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3310.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3313.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3330.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3339.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3340.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3346.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3347.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3352.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3349.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3351.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3354.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3342.4]
  assign ctrs_0_clock = clock; // @[:@3311.4]
  assign ctrs_0_reset = reset; // @[:@3312.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3327.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3319.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3326.4]
  assign ctrs_1_clock = clock; // @[:@3314.4]
  assign ctrs_1_reset = reset; // @[:@3315.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3329.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3323.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3324.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3394.2]
  input   clock, // @[:@3395.4]
  input   reset, // @[:@3396.4]
  input   io_flow, // @[:@3397.4]
  input   io_in, // @[:@3397.4]
  output  io_out // @[:@3397.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3399.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3412.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3411.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3410.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3409.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3408.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3406.4]
endmodule
module RetimeWrapper_25( // @[:@3522.2]
  input   clock, // @[:@3523.4]
  input   reset, // @[:@3524.4]
  input   io_flow, // @[:@3525.4]
  input   io_in, // @[:@3525.4]
  output  io_out // @[:@3525.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@3527.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3540.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3539.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3538.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3537.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3536.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3534.4]
endmodule
module x230_inr_Foreach_sm( // @[:@3542.2]
  input   clock, // @[:@3543.4]
  input   reset, // @[:@3544.4]
  input   io_enable, // @[:@3545.4]
  output  io_done, // @[:@3545.4]
  output  io_doneLatch, // @[:@3545.4]
  input   io_ctrDone, // @[:@3545.4]
  output  io_datapathEn, // @[:@3545.4]
  output  io_ctrInc, // @[:@3545.4]
  output  io_ctrRst, // @[:@3545.4]
  input   io_parentAck, // @[:@3545.4]
  input   io_backpressure, // @[:@3545.4]
  input   io_break // @[:@3545.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3547.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3547.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3550.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3550.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3642.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3555.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3556.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3557.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3558.4]
  wire  _T_100; // @[package.scala 100:49:@3575.4]
  reg  _T_103; // @[package.scala 48:56:@3576.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  wire  _T_110; // @[package.scala 100:49:@3591.4]
  reg  _T_113; // @[package.scala 48:56:@3592.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3594.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3599.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3600.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3603.4]
  wire  _T_124; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  wire  _T_126; // @[package.scala 100:49:@3613.4]
  reg  _T_129; // @[package.scala 48:56:@3614.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3636.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3638.4]
  reg  _T_153; // @[package.scala 48:56:@3639.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3649.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3650.4]
  SRFF active ( // @[Controllers.scala 261:22:@3547.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3550.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3584.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3606.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3618.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3626.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3642.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3555.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3556.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3557.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3558.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3575.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3591.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3594.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3599.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3600.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3603.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3613.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3638.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3649.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3650.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3617.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3652.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3602.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3605.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3597.4]
  assign active_clock = clock; // @[:@3548.4]
  assign active_reset = reset; // @[:@3549.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3560.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3564.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3565.4]
  assign done_clock = clock; // @[:@3551.4]
  assign done_reset = reset; // @[:@3552.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3580.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3573.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3574.4]
  assign RetimeWrapper_clock = clock; // @[:@3585.4]
  assign RetimeWrapper_reset = reset; // @[:@3586.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3588.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3587.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3607.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3608.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3610.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3609.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3619.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3620.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3622.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3621.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3627.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3628.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3630.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3629.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3643.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3644.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3646.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3645.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@3759.2]
  input  [31:0] io_a, // @[:@3762.4]
  output [31:0] io_b // @[:@3762.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@3775.4]
endmodule
module _( // @[:@3777.2]
  input  [31:0] io_b, // @[:@3780.4]
  output [31:0] io_result // @[:@3780.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3785.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3785.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@3785.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3793.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3788.4]
endmodule
module fix2fixBox_2( // @[:@3831.2]
  input  [31:0] io_a, // @[:@3834.4]
  output [32:0] io_b // @[:@3834.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3844.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3844.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@3849.4]
endmodule
module __2( // @[:@3851.2]
  input  [31:0] io_b, // @[:@3854.4]
  output [32:0] io_result // @[:@3854.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3859.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3859.4]
  fix2fixBox_2 fix2fixBox ( // @[BigIPZynq.scala 219:30:@3859.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3867.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3862.4]
endmodule
module RetimeWrapper_29( // @[:@3919.2]
  input         clock, // @[:@3920.4]
  input         reset, // @[:@3921.4]
  input         io_flow, // @[:@3922.4]
  input  [31:0] io_in, // @[:@3922.4]
  output [31:0] io_out // @[:@3922.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3924.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3937.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3936.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3935.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3934.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3933.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3931.4]
endmodule
module fix2fixBox_4( // @[:@3939.2]
  input         clock, // @[:@3940.4]
  input         reset, // @[:@3941.4]
  input  [32:0] io_a, // @[:@3942.4]
  input         io_flow, // @[:@3942.4]
  output [31:0] io_b // @[:@3942.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3955.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3955.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3962.4]
  assign RetimeWrapper_clock = clock; // @[:@3956.4]
  assign RetimeWrapper_reset = reset; // @[:@3957.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3959.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3958.4]
endmodule
module x410_sub( // @[:@3964.2]
  input         clock, // @[:@3965.4]
  input         reset, // @[:@3966.4]
  input  [31:0] io_a, // @[:@3967.4]
  input  [31:0] io_b, // @[:@3967.4]
  input         io_flow, // @[:@3967.4]
  output [31:0] io_result // @[:@3967.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3975.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3975.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3982.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3982.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4001.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4001.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4001.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@3989.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@3990.4]
  __2 _ ( // @[Math.scala 720:24:@3975.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@3982.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@4001.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@3989.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@3990.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4009.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3978.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3985.4]
  assign fix2fixBox_clock = clock; // @[:@4002.4]
  assign fix2fixBox_reset = reset; // @[:@4003.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4004.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4007.4]
endmodule
module x223_sum( // @[:@4176.2]
  input         clock, // @[:@4177.4]
  input         reset, // @[:@4178.4]
  input  [31:0] io_a, // @[:@4179.4]
  input  [31:0] io_b, // @[:@4179.4]
  input         io_flow, // @[:@4179.4]
  output [31:0] io_result // @[:@4179.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4187.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@4187.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4194.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@4194.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4212.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4212.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4212.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4201.4]
  __2 _ ( // @[Math.scala 720:24:@4187.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@4194.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@4212.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4201.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4220.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@4190.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@4197.4]
  assign fix2fixBox_clock = clock; // @[:@4213.4]
  assign fix2fixBox_reset = reset; // @[:@4214.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4215.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4218.4]
endmodule
module x230_inr_Foreach_kernelx230_inr_Foreach_concrete1( // @[:@4533.2]
  input         clock, // @[:@4534.4]
  input         reset, // @[:@4535.4]
  output        io_in_x213_fifoinpacked_0_wPort_0_en_0, // @[:@4536.4]
  input         io_in_x213_fifoinpacked_0_full, // @[:@4536.4]
  output        io_in_x213_fifoinpacked_0_active_0_in, // @[:@4536.4]
  input         io_in_x213_fifoinpacked_0_active_0_out, // @[:@4536.4]
  input         io_sigsIn_backpressure, // @[:@4536.4]
  input         io_sigsIn_datapathEn, // @[:@4536.4]
  input         io_sigsIn_break, // @[:@4536.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@4536.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@4536.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@4536.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@4536.4]
  input         io_rr // @[:@4536.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4570.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@4570.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4582.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@4582.4]
  wire  x410_sub_1_clock; // @[Math.scala 191:24:@4609.4]
  wire  x410_sub_1_reset; // @[Math.scala 191:24:@4609.4]
  wire [31:0] x410_sub_1_io_a; // @[Math.scala 191:24:@4609.4]
  wire [31:0] x410_sub_1_io_b; // @[Math.scala 191:24:@4609.4]
  wire  x410_sub_1_io_flow; // @[Math.scala 191:24:@4609.4]
  wire [31:0] x410_sub_1_io_result; // @[Math.scala 191:24:@4609.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4619.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4619.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4619.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@4619.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@4619.4]
  wire  x223_sum_1_clock; // @[Math.scala 150:24:@4628.4]
  wire  x223_sum_1_reset; // @[Math.scala 150:24:@4628.4]
  wire [31:0] x223_sum_1_io_a; // @[Math.scala 150:24:@4628.4]
  wire [31:0] x223_sum_1_io_b; // @[Math.scala 150:24:@4628.4]
  wire  x223_sum_1_io_flow; // @[Math.scala 150:24:@4628.4]
  wire [31:0] x223_sum_1_io_result; // @[Math.scala 150:24:@4628.4]
  wire  x224_sum_1_clock; // @[Math.scala 150:24:@4640.4]
  wire  x224_sum_1_reset; // @[Math.scala 150:24:@4640.4]
  wire [31:0] x224_sum_1_io_a; // @[Math.scala 150:24:@4640.4]
  wire [31:0] x224_sum_1_io_b; // @[Math.scala 150:24:@4640.4]
  wire  x224_sum_1_io_flow; // @[Math.scala 150:24:@4640.4]
  wire [31:0] x224_sum_1_io_result; // @[Math.scala 150:24:@4640.4]
  wire [31:0] x226_1_io_b; // @[Math.scala 720:24:@4661.4]
  wire [31:0] x226_1_io_result; // @[Math.scala 720:24:@4661.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4674.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4674.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@4674.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4674.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4674.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@4683.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@4683.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@4683.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@4683.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@4683.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@4694.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@4694.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@4694.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@4694.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@4694.4]
  wire  _T_327; // @[sm_x230_inr_Foreach.scala 62:18:@4595.4]
  wire  _T_328; // @[sm_x230_inr_Foreach.scala 62:55:@4596.4]
  wire [31:0] b218_number; // @[Math.scala 723:22:@4575.4 Math.scala 724:14:@4576.4]
  wire [42:0] _GEN_0; // @[Math.scala 461:32:@4600.4]
  wire [42:0] _T_331; // @[Math.scala 461:32:@4600.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@4605.4]
  wire [38:0] _T_334; // @[Math.scala 461:32:@4605.4]
  wire [31:0] x224_sum_number; // @[Math.scala 154:22:@4646.4 Math.scala 155:14:@4647.4]
  wire [31:0] _T_358; // @[Math.scala 406:49:@4653.4]
  wire [31:0] _T_360; // @[Math.scala 406:56:@4655.4]
  wire [31:0] _T_361; // @[Math.scala 406:56:@4656.4]
  wire  _T_379; // @[sm_x230_inr_Foreach.scala 89:131:@4691.4]
  wire  _T_383; // @[package.scala 96:25:@4699.4 package.scala 96:25:@4700.4]
  wire  _T_385; // @[implicits.scala 55:10:@4701.4]
  wire  _T_386; // @[sm_x230_inr_Foreach.scala 89:148:@4702.4]
  wire  _T_388; // @[sm_x230_inr_Foreach.scala 89:236:@4704.4]
  wire  _T_389; // @[sm_x230_inr_Foreach.scala 89:255:@4705.4]
  wire  x496_b220_D3; // @[package.scala 96:25:@4679.4 package.scala 96:25:@4680.4]
  wire  _T_392; // @[sm_x230_inr_Foreach.scala 89:291:@4707.4]
  wire  x497_b221_D3; // @[package.scala 96:25:@4688.4 package.scala 96:25:@4689.4]
  _ _ ( // @[Math.scala 720:24:@4570.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@4582.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x410_sub x410_sub_1 ( // @[Math.scala 191:24:@4609.4]
    .clock(x410_sub_1_clock),
    .reset(x410_sub_1_reset),
    .io_a(x410_sub_1_io_a),
    .io_b(x410_sub_1_io_b),
    .io_flow(x410_sub_1_io_flow),
    .io_result(x410_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@4619.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x223_sum x223_sum_1 ( // @[Math.scala 150:24:@4628.4]
    .clock(x223_sum_1_clock),
    .reset(x223_sum_1_reset),
    .io_a(x223_sum_1_io_a),
    .io_b(x223_sum_1_io_b),
    .io_flow(x223_sum_1_io_flow),
    .io_result(x223_sum_1_io_result)
  );
  x223_sum x224_sum_1 ( // @[Math.scala 150:24:@4640.4]
    .clock(x224_sum_1_clock),
    .reset(x224_sum_1_reset),
    .io_a(x224_sum_1_io_a),
    .io_b(x224_sum_1_io_b),
    .io_flow(x224_sum_1_io_flow),
    .io_result(x224_sum_1_io_result)
  );
  _ x226_1 ( // @[Math.scala 720:24:@4661.4]
    .io_b(x226_1_io_b),
    .io_result(x226_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@4674.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@4683.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@4694.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_327 = ~ io_in_x213_fifoinpacked_0_full; // @[sm_x230_inr_Foreach.scala 62:18:@4595.4]
  assign _T_328 = ~ io_in_x213_fifoinpacked_0_active_0_out; // @[sm_x230_inr_Foreach.scala 62:55:@4596.4]
  assign b218_number = __io_result; // @[Math.scala 723:22:@4575.4 Math.scala 724:14:@4576.4]
  assign _GEN_0 = {{11'd0}, b218_number}; // @[Math.scala 461:32:@4600.4]
  assign _T_331 = _GEN_0 << 11; // @[Math.scala 461:32:@4600.4]
  assign _GEN_1 = {{7'd0}, b218_number}; // @[Math.scala 461:32:@4605.4]
  assign _T_334 = _GEN_1 << 7; // @[Math.scala 461:32:@4605.4]
  assign x224_sum_number = x224_sum_1_io_result; // @[Math.scala 154:22:@4646.4 Math.scala 155:14:@4647.4]
  assign _T_358 = $signed(x224_sum_number); // @[Math.scala 406:49:@4653.4]
  assign _T_360 = $signed(_T_358) & $signed(32'shff); // @[Math.scala 406:56:@4655.4]
  assign _T_361 = $signed(_T_360); // @[Math.scala 406:56:@4656.4]
  assign _T_379 = ~ io_sigsIn_break; // @[sm_x230_inr_Foreach.scala 89:131:@4691.4]
  assign _T_383 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@4699.4 package.scala 96:25:@4700.4]
  assign _T_385 = io_rr ? _T_383 : 1'h0; // @[implicits.scala 55:10:@4701.4]
  assign _T_386 = _T_379 & _T_385; // @[sm_x230_inr_Foreach.scala 89:148:@4702.4]
  assign _T_388 = _T_386 & _T_379; // @[sm_x230_inr_Foreach.scala 89:236:@4704.4]
  assign _T_389 = _T_388 & io_sigsIn_backpressure; // @[sm_x230_inr_Foreach.scala 89:255:@4705.4]
  assign x496_b220_D3 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4679.4 package.scala 96:25:@4680.4]
  assign _T_392 = _T_389 & x496_b220_D3; // @[sm_x230_inr_Foreach.scala 89:291:@4707.4]
  assign x497_b221_D3 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@4688.4 package.scala 96:25:@4689.4]
  assign io_in_x213_fifoinpacked_0_wPort_0_en_0 = _T_392 & x497_b221_D3; // @[MemInterfaceType.scala 93:57:@4711.4]
  assign io_in_x213_fifoinpacked_0_active_0_in = x496_b220_D3 & x497_b221_D3; // @[MemInterfaceType.scala 147:18:@4714.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@4573.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@4585.4]
  assign x410_sub_1_clock = clock; // @[:@4610.4]
  assign x410_sub_1_reset = reset; // @[:@4611.4]
  assign x410_sub_1_io_a = _T_331[31:0]; // @[Math.scala 192:17:@4612.4]
  assign x410_sub_1_io_b = _T_334[31:0]; // @[Math.scala 193:17:@4613.4]
  assign x410_sub_1_io_flow = _T_327 | _T_328; // @[Math.scala 194:20:@4614.4]
  assign RetimeWrapper_clock = clock; // @[:@4620.4]
  assign RetimeWrapper_reset = reset; // @[:@4621.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4623.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@4622.4]
  assign x223_sum_1_clock = clock; // @[:@4629.4]
  assign x223_sum_1_reset = reset; // @[:@4630.4]
  assign x223_sum_1_io_a = x410_sub_1_io_result; // @[Math.scala 151:17:@4631.4]
  assign x223_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@4632.4]
  assign x223_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4633.4]
  assign x224_sum_1_clock = clock; // @[:@4641.4]
  assign x224_sum_1_reset = reset; // @[:@4642.4]
  assign x224_sum_1_io_a = x223_sum_1_io_result; // @[Math.scala 151:17:@4643.4]
  assign x224_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@4644.4]
  assign x224_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4645.4]
  assign x226_1_io_b = $unsigned(_T_361); // @[Math.scala 721:17:@4664.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4675.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4676.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4678.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@4677.4]
  assign RetimeWrapper_2_clock = clock; // @[:@4684.4]
  assign RetimeWrapper_2_reset = reset; // @[:@4685.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4687.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@4686.4]
  assign RetimeWrapper_3_clock = clock; // @[:@4695.4]
  assign RetimeWrapper_3_reset = reset; // @[:@4696.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4698.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@4697.4]
endmodule
module RetimeWrapper_41( // @[:@5832.2]
  input   clock, // @[:@5833.4]
  input   reset, // @[:@5834.4]
  input   io_flow, // @[:@5835.4]
  input   io_in, // @[:@5835.4]
  output  io_out // @[:@5835.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@5837.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@5837.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@5837.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@5837.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@5837.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@5837.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(145)) sr ( // @[RetimeShiftRegister.scala 15:20:@5837.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@5850.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@5849.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@5848.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@5847.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@5846.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@5844.4]
endmodule
module RetimeWrapper_45( // @[:@5960.2]
  input   clock, // @[:@5961.4]
  input   reset, // @[:@5962.4]
  input   io_flow, // @[:@5963.4]
  input   io_in, // @[:@5963.4]
  output  io_out // @[:@5963.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@5965.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@5965.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@5965.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@5965.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@5965.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@5965.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(144)) sr ( // @[RetimeShiftRegister.scala 15:20:@5965.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@5978.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@5977.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@5976.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@5975.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@5974.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@5972.4]
endmodule
module x359_inr_Foreach_SAMPLER_BOX_sm( // @[:@5980.2]
  input   clock, // @[:@5981.4]
  input   reset, // @[:@5982.4]
  input   io_enable, // @[:@5983.4]
  output  io_done, // @[:@5983.4]
  output  io_doneLatch, // @[:@5983.4]
  input   io_ctrDone, // @[:@5983.4]
  output  io_datapathEn, // @[:@5983.4]
  output  io_ctrInc, // @[:@5983.4]
  output  io_ctrRst, // @[:@5983.4]
  input   io_parentAck, // @[:@5983.4]
  input   io_backpressure, // @[:@5983.4]
  input   io_break // @[:@5983.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@5985.4]
  wire  active_reset; // @[Controllers.scala 261:22:@5985.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@5985.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@5985.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@5985.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@5985.4]
  wire  done_clock; // @[Controllers.scala 262:20:@5988.4]
  wire  done_reset; // @[Controllers.scala 262:20:@5988.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@5988.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@5988.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@5988.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@5988.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6022.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6022.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6022.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6022.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6022.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6044.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6044.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6044.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6044.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6044.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6056.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6056.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6056.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6056.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6056.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6064.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6064.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6064.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6064.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6064.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6080.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6080.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@6080.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6080.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6080.4]
  wire  _T_80; // @[Controllers.scala 264:48:@5993.4]
  wire  _T_81; // @[Controllers.scala 264:46:@5994.4]
  wire  _T_82; // @[Controllers.scala 264:62:@5995.4]
  wire  _T_83; // @[Controllers.scala 264:60:@5996.4]
  wire  _T_100; // @[package.scala 100:49:@6013.4]
  reg  _T_103; // @[package.scala 48:56:@6014.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@6027.4 package.scala 96:25:@6028.4]
  wire  _T_110; // @[package.scala 100:49:@6029.4]
  reg  _T_113; // @[package.scala 48:56:@6030.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@6032.4]
  wire  _T_118; // @[Controllers.scala 283:41:@6037.4]
  wire  _T_119; // @[Controllers.scala 283:59:@6038.4]
  wire  _T_121; // @[Controllers.scala 284:37:@6041.4]
  wire  _T_124; // @[package.scala 96:25:@6049.4 package.scala 96:25:@6050.4]
  wire  _T_126; // @[package.scala 100:49:@6051.4]
  reg  _T_129; // @[package.scala 48:56:@6052.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@6074.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@6076.4]
  reg  _T_153; // @[package.scala 48:56:@6077.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@6085.4 package.scala 96:25:@6086.4]
  wire  _T_158; // @[Controllers.scala 292:61:@6087.4]
  wire  _T_159; // @[Controllers.scala 292:24:@6088.4]
  SRFF active ( // @[Controllers.scala 261:22:@5985.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@5988.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_41 RetimeWrapper ( // @[package.scala 93:22:@6022.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_41 RetimeWrapper_1 ( // @[package.scala 93:22:@6044.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6056.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6064.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_45 RetimeWrapper_4 ( // @[package.scala 93:22:@6080.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@5993.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@5994.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@5995.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@5996.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@6013.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@6027.4 package.scala 96:25:@6028.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@6029.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@6032.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@6037.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@6038.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@6041.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6049.4 package.scala 96:25:@6050.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6051.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6076.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@6085.4 package.scala 96:25:@6086.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@6087.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@6088.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6055.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@6090.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@6040.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@6043.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@6035.4]
  assign active_clock = clock; // @[:@5986.4]
  assign active_reset = reset; // @[:@5987.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@5998.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@6002.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@6003.4]
  assign done_clock = clock; // @[:@5989.4]
  assign done_reset = reset; // @[:@5990.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@6018.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@6011.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@6012.4]
  assign RetimeWrapper_clock = clock; // @[:@6023.4]
  assign RetimeWrapper_reset = reset; // @[:@6024.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@6026.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@6025.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6045.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6046.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@6048.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6047.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6057.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6058.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6060.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6059.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6065.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6066.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6068.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6067.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6081.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6082.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@6084.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@6083.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SRAM_1( // @[:@6317.2]
  input         clock, // @[:@6318.4]
  input         reset, // @[:@6319.4]
  input  [9:0]  io_raddr, // @[:@6320.4]
  input         io_wen, // @[:@6320.4]
  input  [9:0]  io_waddr, // @[:@6320.4]
  input  [31:0] io_wdata, // @[:@6320.4]
  output [31:0] io_rdata, // @[:@6320.4]
  input         io_backpressure // @[:@6320.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@6322.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@6322.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@6322.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@6322.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@6322.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@6322.4]
  wire [9:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@6322.4]
  wire [9:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@6322.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@6322.4]
  wire  _T_19; // @[SRAM.scala 182:49:@6340.4]
  wire  _T_20; // @[SRAM.scala 182:37:@6341.4]
  reg  _T_23; // @[SRAM.scala 182:29:@6342.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@6344.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(640), .AWIDTH(10)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@6322.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@6340.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@6341.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@6349.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@6336.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@6337.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@6334.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@6339.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@6338.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@6335.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@6333.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@6332.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_50( // @[:@6363.2]
  input        clock, // @[:@6364.4]
  input        reset, // @[:@6365.4]
  input        io_flow, // @[:@6366.4]
  input  [9:0] io_in, // @[:@6366.4]
  output [9:0] io_out // @[:@6366.4]
);
  wire [9:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@6368.4]
  wire [9:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@6368.4]
  wire [9:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@6368.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6368.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6368.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6368.4]
  RetimeShiftRegister #(.WIDTH(10), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@6368.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6381.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6380.4]
  assign sr_init = 10'h0; // @[RetimeShiftRegister.scala 19:16:@6379.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6378.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6377.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6375.4]
endmodule
module Mem1D_5( // @[:@6383.2]
  input         clock, // @[:@6384.4]
  input         reset, // @[:@6385.4]
  input  [9:0]  io_r_ofs_0, // @[:@6386.4]
  input         io_r_backpressure, // @[:@6386.4]
  input  [9:0]  io_w_ofs_0, // @[:@6386.4]
  input  [31:0] io_w_data_0, // @[:@6386.4]
  input         io_w_en_0, // @[:@6386.4]
  output [31:0] io_output // @[:@6386.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@6390.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 715:21:@6390.4]
  wire [9:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@6390.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 715:21:@6390.4]
  wire [9:0] SRAM_io_waddr; // @[MemPrimitives.scala 715:21:@6390.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 715:21:@6390.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@6390.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@6390.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6393.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6393.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6393.4]
  wire [9:0] RetimeWrapper_io_in; // @[package.scala 93:22:@6393.4]
  wire [9:0] RetimeWrapper_io_out; // @[package.scala 93:22:@6393.4]
  wire  wInBound; // @[MemPrimitives.scala 702:32:@6388.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 715:21:@6390.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_50 RetimeWrapper ( // @[package.scala 93:22:@6393.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 10'h280; // @[MemPrimitives.scala 702:32:@6388.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@6406.4]
  assign SRAM_clock = clock; // @[:@6391.4]
  assign SRAM_reset = reset; // @[:@6392.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@6400.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 719:22:@6403.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 718:22:@6401.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 720:22:@6404.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@6405.4]
  assign RetimeWrapper_clock = clock; // @[:@6394.4]
  assign RetimeWrapper_reset = reset; // @[:@6395.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@6397.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@6396.4]
endmodule
module StickySelects_1( // @[:@7585.2]
  input   clock, // @[:@7586.4]
  input   reset, // @[:@7587.4]
  input   io_ins_0, // @[:@7588.4]
  input   io_ins_1, // @[:@7588.4]
  input   io_ins_2, // @[:@7588.4]
  input   io_ins_3, // @[:@7588.4]
  input   io_ins_4, // @[:@7588.4]
  input   io_ins_5, // @[:@7588.4]
  input   io_ins_6, // @[:@7588.4]
  input   io_ins_7, // @[:@7588.4]
  input   io_ins_8, // @[:@7588.4]
  output  io_outs_0, // @[:@7588.4]
  output  io_outs_1, // @[:@7588.4]
  output  io_outs_2, // @[:@7588.4]
  output  io_outs_3, // @[:@7588.4]
  output  io_outs_4, // @[:@7588.4]
  output  io_outs_5, // @[:@7588.4]
  output  io_outs_6, // @[:@7588.4]
  output  io_outs_7, // @[:@7588.4]
  output  io_outs_8 // @[:@7588.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@7590.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@7591.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@7592.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@7593.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@7594.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@7595.4]
  reg [31:0] _RAND_5;
  reg  _T_37; // @[StickySelects.scala 37:46:@7596.4]
  reg [31:0] _RAND_6;
  reg  _T_40; // @[StickySelects.scala 37:46:@7597.4]
  reg [31:0] _RAND_7;
  reg  _T_43; // @[StickySelects.scala 37:46:@7598.4]
  reg [31:0] _RAND_8;
  wire  _T_44; // @[StickySelects.scala 47:46:@7599.4]
  wire  _T_45; // @[StickySelects.scala 47:46:@7600.4]
  wire  _T_46; // @[StickySelects.scala 47:46:@7601.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@7602.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@7603.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@7604.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@7605.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@7606.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@7607.4]
  wire  _T_53; // @[StickySelects.scala 47:46:@7609.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@7610.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@7611.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@7612.4]
  wire  _T_57; // @[StickySelects.scala 47:46:@7613.4]
  wire  _T_58; // @[StickySelects.scala 47:46:@7614.4]
  wire  _T_59; // @[StickySelects.scala 47:46:@7615.4]
  wire  _T_60; // @[StickySelects.scala 49:53:@7616.4]
  wire  _T_61; // @[StickySelects.scala 49:21:@7617.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@7619.4]
  wire  _T_63; // @[StickySelects.scala 47:46:@7620.4]
  wire  _T_64; // @[StickySelects.scala 47:46:@7621.4]
  wire  _T_65; // @[StickySelects.scala 47:46:@7622.4]
  wire  _T_66; // @[StickySelects.scala 47:46:@7623.4]
  wire  _T_67; // @[StickySelects.scala 47:46:@7624.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@7625.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@7626.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@7627.4]
  wire  _T_72; // @[StickySelects.scala 47:46:@7630.4]
  wire  _T_73; // @[StickySelects.scala 47:46:@7631.4]
  wire  _T_74; // @[StickySelects.scala 47:46:@7632.4]
  wire  _T_75; // @[StickySelects.scala 47:46:@7633.4]
  wire  _T_76; // @[StickySelects.scala 47:46:@7634.4]
  wire  _T_77; // @[StickySelects.scala 47:46:@7635.4]
  wire  _T_78; // @[StickySelects.scala 49:53:@7636.4]
  wire  _T_79; // @[StickySelects.scala 49:21:@7637.4]
  wire  _T_82; // @[StickySelects.scala 47:46:@7641.4]
  wire  _T_83; // @[StickySelects.scala 47:46:@7642.4]
  wire  _T_84; // @[StickySelects.scala 47:46:@7643.4]
  wire  _T_85; // @[StickySelects.scala 47:46:@7644.4]
  wire  _T_86; // @[StickySelects.scala 47:46:@7645.4]
  wire  _T_87; // @[StickySelects.scala 49:53:@7646.4]
  wire  _T_88; // @[StickySelects.scala 49:21:@7647.4]
  wire  _T_92; // @[StickySelects.scala 47:46:@7652.4]
  wire  _T_93; // @[StickySelects.scala 47:46:@7653.4]
  wire  _T_94; // @[StickySelects.scala 47:46:@7654.4]
  wire  _T_95; // @[StickySelects.scala 47:46:@7655.4]
  wire  _T_96; // @[StickySelects.scala 49:53:@7656.4]
  wire  _T_97; // @[StickySelects.scala 49:21:@7657.4]
  wire  _T_102; // @[StickySelects.scala 47:46:@7663.4]
  wire  _T_103; // @[StickySelects.scala 47:46:@7664.4]
  wire  _T_104; // @[StickySelects.scala 47:46:@7665.4]
  wire  _T_105; // @[StickySelects.scala 49:53:@7666.4]
  wire  _T_106; // @[StickySelects.scala 49:21:@7667.4]
  wire  _T_112; // @[StickySelects.scala 47:46:@7674.4]
  wire  _T_113; // @[StickySelects.scala 47:46:@7675.4]
  wire  _T_114; // @[StickySelects.scala 49:53:@7676.4]
  wire  _T_115; // @[StickySelects.scala 49:21:@7677.4]
  wire  _T_122; // @[StickySelects.scala 47:46:@7685.4]
  wire  _T_123; // @[StickySelects.scala 49:53:@7686.4]
  wire  _T_124; // @[StickySelects.scala 49:21:@7687.4]
  assign _T_44 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@7599.4]
  assign _T_45 = _T_44 | io_ins_3; // @[StickySelects.scala 47:46:@7600.4]
  assign _T_46 = _T_45 | io_ins_4; // @[StickySelects.scala 47:46:@7601.4]
  assign _T_47 = _T_46 | io_ins_5; // @[StickySelects.scala 47:46:@7602.4]
  assign _T_48 = _T_47 | io_ins_6; // @[StickySelects.scala 47:46:@7603.4]
  assign _T_49 = _T_48 | io_ins_7; // @[StickySelects.scala 47:46:@7604.4]
  assign _T_50 = _T_49 | io_ins_8; // @[StickySelects.scala 47:46:@7605.4]
  assign _T_51 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@7606.4]
  assign _T_52 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 49:21:@7607.4]
  assign _T_53 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@7609.4]
  assign _T_54 = _T_53 | io_ins_3; // @[StickySelects.scala 47:46:@7610.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@7611.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@7612.4]
  assign _T_57 = _T_56 | io_ins_6; // @[StickySelects.scala 47:46:@7613.4]
  assign _T_58 = _T_57 | io_ins_7; // @[StickySelects.scala 47:46:@7614.4]
  assign _T_59 = _T_58 | io_ins_8; // @[StickySelects.scala 47:46:@7615.4]
  assign _T_60 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@7616.4]
  assign _T_61 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 49:21:@7617.4]
  assign _T_62 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@7619.4]
  assign _T_63 = _T_62 | io_ins_3; // @[StickySelects.scala 47:46:@7620.4]
  assign _T_64 = _T_63 | io_ins_4; // @[StickySelects.scala 47:46:@7621.4]
  assign _T_65 = _T_64 | io_ins_5; // @[StickySelects.scala 47:46:@7622.4]
  assign _T_66 = _T_65 | io_ins_6; // @[StickySelects.scala 47:46:@7623.4]
  assign _T_67 = _T_66 | io_ins_7; // @[StickySelects.scala 47:46:@7624.4]
  assign _T_68 = _T_67 | io_ins_8; // @[StickySelects.scala 47:46:@7625.4]
  assign _T_69 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@7626.4]
  assign _T_70 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 49:21:@7627.4]
  assign _T_72 = _T_62 | io_ins_2; // @[StickySelects.scala 47:46:@7630.4]
  assign _T_73 = _T_72 | io_ins_4; // @[StickySelects.scala 47:46:@7631.4]
  assign _T_74 = _T_73 | io_ins_5; // @[StickySelects.scala 47:46:@7632.4]
  assign _T_75 = _T_74 | io_ins_6; // @[StickySelects.scala 47:46:@7633.4]
  assign _T_76 = _T_75 | io_ins_7; // @[StickySelects.scala 47:46:@7634.4]
  assign _T_77 = _T_76 | io_ins_8; // @[StickySelects.scala 47:46:@7635.4]
  assign _T_78 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@7636.4]
  assign _T_79 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 49:21:@7637.4]
  assign _T_82 = _T_72 | io_ins_3; // @[StickySelects.scala 47:46:@7641.4]
  assign _T_83 = _T_82 | io_ins_5; // @[StickySelects.scala 47:46:@7642.4]
  assign _T_84 = _T_83 | io_ins_6; // @[StickySelects.scala 47:46:@7643.4]
  assign _T_85 = _T_84 | io_ins_7; // @[StickySelects.scala 47:46:@7644.4]
  assign _T_86 = _T_85 | io_ins_8; // @[StickySelects.scala 47:46:@7645.4]
  assign _T_87 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@7646.4]
  assign _T_88 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 49:21:@7647.4]
  assign _T_92 = _T_82 | io_ins_4; // @[StickySelects.scala 47:46:@7652.4]
  assign _T_93 = _T_92 | io_ins_6; // @[StickySelects.scala 47:46:@7653.4]
  assign _T_94 = _T_93 | io_ins_7; // @[StickySelects.scala 47:46:@7654.4]
  assign _T_95 = _T_94 | io_ins_8; // @[StickySelects.scala 47:46:@7655.4]
  assign _T_96 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@7656.4]
  assign _T_97 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 49:21:@7657.4]
  assign _T_102 = _T_92 | io_ins_5; // @[StickySelects.scala 47:46:@7663.4]
  assign _T_103 = _T_102 | io_ins_7; // @[StickySelects.scala 47:46:@7664.4]
  assign _T_104 = _T_103 | io_ins_8; // @[StickySelects.scala 47:46:@7665.4]
  assign _T_105 = io_ins_6 | _T_37; // @[StickySelects.scala 49:53:@7666.4]
  assign _T_106 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 49:21:@7667.4]
  assign _T_112 = _T_102 | io_ins_6; // @[StickySelects.scala 47:46:@7674.4]
  assign _T_113 = _T_112 | io_ins_8; // @[StickySelects.scala 47:46:@7675.4]
  assign _T_114 = io_ins_7 | _T_40; // @[StickySelects.scala 49:53:@7676.4]
  assign _T_115 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 49:21:@7677.4]
  assign _T_122 = _T_112 | io_ins_7; // @[StickySelects.scala 47:46:@7685.4]
  assign _T_123 = io_ins_8 | _T_43; // @[StickySelects.scala 49:53:@7686.4]
  assign _T_124 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 49:21:@7687.4]
  assign io_outs_0 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 53:57:@7689.4]
  assign io_outs_1 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 53:57:@7690.4]
  assign io_outs_2 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 53:57:@7691.4]
  assign io_outs_3 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 53:57:@7692.4]
  assign io_outs_4 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 53:57:@7693.4]
  assign io_outs_5 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 53:57:@7694.4]
  assign io_outs_6 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 53:57:@7695.4]
  assign io_outs_7 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 53:57:@7696.4]
  assign io_outs_8 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 53:57:@7697.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_37 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_40 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_43 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_51;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_59) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_60;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_69;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_77) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_78;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_86) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_87;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_95) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_96;
      end
    end
    if (reset) begin
      _T_37 <= 1'h0;
    end else begin
      if (_T_104) begin
        _T_37 <= io_ins_6;
      end else begin
        _T_37 <= _T_105;
      end
    end
    if (reset) begin
      _T_40 <= 1'h0;
    end else begin
      if (_T_113) begin
        _T_40 <= io_ins_7;
      end else begin
        _T_40 <= _T_114;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_122) begin
        _T_43 <= io_ins_8;
      end else begin
        _T_43 <= _T_123;
      end
    end
  end
endmodule
module x241_lb_0( // @[:@12409.2]
  input         clock, // @[:@12410.4]
  input         reset, // @[:@12411.4]
  input  [1:0]  io_rPort_8_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_8_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_8_ofs_0, // @[:@12412.4]
  input         io_rPort_8_en_0, // @[:@12412.4]
  input         io_rPort_8_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_8_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_7_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_7_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_7_ofs_0, // @[:@12412.4]
  input         io_rPort_7_en_0, // @[:@12412.4]
  input         io_rPort_7_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_7_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_6_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_6_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_6_ofs_0, // @[:@12412.4]
  input         io_rPort_6_en_0, // @[:@12412.4]
  input         io_rPort_6_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_6_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_5_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_5_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_5_ofs_0, // @[:@12412.4]
  input         io_rPort_5_en_0, // @[:@12412.4]
  input         io_rPort_5_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_5_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_4_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_4_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_4_ofs_0, // @[:@12412.4]
  input         io_rPort_4_en_0, // @[:@12412.4]
  input         io_rPort_4_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_4_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_3_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_3_ofs_0, // @[:@12412.4]
  input         io_rPort_3_en_0, // @[:@12412.4]
  input         io_rPort_3_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_3_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_2_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_2_ofs_0, // @[:@12412.4]
  input         io_rPort_2_en_0, // @[:@12412.4]
  input         io_rPort_2_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_2_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_1_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_1_ofs_0, // @[:@12412.4]
  input         io_rPort_1_en_0, // @[:@12412.4]
  input         io_rPort_1_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_1_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_0_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_0_ofs_0, // @[:@12412.4]
  input         io_rPort_0_en_0, // @[:@12412.4]
  input         io_rPort_0_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_0_output_0, // @[:@12412.4]
  input  [1:0]  io_wPort_0_banks_1, // @[:@12412.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@12412.4]
  input  [9:0]  io_wPort_0_ofs_0, // @[:@12412.4]
  input  [31:0] io_wPort_0_data_0, // @[:@12412.4]
  input         io_wPort_0_en_0 // @[:@12412.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@12477.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@12477.4]
  wire [9:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12477.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12477.4]
  wire [9:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12477.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@12477.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@12477.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@12477.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@12493.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@12493.4]
  wire [9:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12493.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12493.4]
  wire [9:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12493.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@12493.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@12493.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@12493.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@12509.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@12509.4]
  wire [9:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12509.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12509.4]
  wire [9:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12509.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@12509.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@12509.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@12509.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@12525.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@12525.4]
  wire [9:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12525.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12525.4]
  wire [9:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12525.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@12525.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@12525.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@12525.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@12541.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@12541.4]
  wire [9:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12541.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12541.4]
  wire [9:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12541.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@12541.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@12541.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@12541.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@12557.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@12557.4]
  wire [9:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12557.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12557.4]
  wire [9:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12557.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@12557.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@12557.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@12557.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@12573.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@12573.4]
  wire [9:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12573.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12573.4]
  wire [9:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12573.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@12573.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@12573.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@12573.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@12589.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@12589.4]
  wire [9:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12589.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12589.4]
  wire [9:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12589.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@12589.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@12589.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@12589.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@12605.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@12605.4]
  wire [9:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12605.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12605.4]
  wire [9:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12605.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@12605.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@12605.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@12605.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@12621.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@12621.4]
  wire [9:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12621.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12621.4]
  wire [9:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12621.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@12621.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@12621.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@12621.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@12637.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@12637.4]
  wire [9:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12637.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12637.4]
  wire [9:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12637.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@12637.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@12637.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@12637.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@12653.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@12653.4]
  wire [9:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12653.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12653.4]
  wire [9:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12653.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@12653.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@12653.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@12653.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_6; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_7; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_8; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_6; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_7; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_8; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_6; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_7; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_8; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_6; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_7; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_8; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_8; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_8; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_8; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_8; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_6; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_7; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_8; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_6; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_7; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_8; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_6; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_7; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_8; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_6; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_7; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_8; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_8; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_8; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_8; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_8; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_6; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_7; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_8; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_6; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_7; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_8; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_6; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_7; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_8; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_6; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_7; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_8; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_8; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_8; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_8; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_8; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@13918.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@13918.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@13918.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@13918.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@13918.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@13926.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@13926.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@13926.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@13926.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@13926.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@13934.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@13934.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@13934.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@13934.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@13934.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@13942.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@13942.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@13942.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@13942.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@13942.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@13950.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@13950.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@13950.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@13950.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@13950.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@13958.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@13958.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@13958.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@13958.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@13958.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@13966.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@13966.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@13966.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@13966.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@13966.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@13974.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@13974.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@13974.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@13974.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@13974.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@13982.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@13982.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@13982.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@13982.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@13982.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@13990.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@13990.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@13990.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@13990.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@13990.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@13998.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@13998.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@13998.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@13998.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@13998.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@14006.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@14006.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@14006.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@14006.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@14006.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@14062.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@14062.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@14062.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@14062.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@14062.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@14070.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@14070.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@14070.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@14070.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@14070.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@14078.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@14078.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@14078.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@14078.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@14078.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@14086.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@14086.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@14086.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@14086.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@14086.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@14094.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@14094.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@14094.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@14094.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@14094.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@14102.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@14102.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@14102.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@14102.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@14102.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@14110.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@14110.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@14110.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@14110.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@14110.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@14118.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@14118.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@14118.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@14118.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@14118.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@14126.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@14126.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@14126.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@14126.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@14126.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@14134.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@14134.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@14134.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@14134.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@14134.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@14142.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@14142.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@14142.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@14142.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@14142.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@14150.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@14150.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@14150.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@14150.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@14150.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@14206.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@14206.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@14206.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@14206.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@14206.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@14214.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@14214.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@14214.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@14214.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@14214.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@14222.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@14222.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@14222.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@14222.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@14222.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@14230.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@14230.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@14230.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@14230.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@14230.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@14238.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@14238.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@14238.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@14238.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@14238.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@14246.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@14246.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@14246.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@14246.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@14246.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@14254.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@14254.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@14254.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@14254.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@14254.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@14262.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@14262.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@14262.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@14262.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@14262.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@14270.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@14270.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@14270.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@14270.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@14270.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@14278.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@14278.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@14278.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@14278.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@14278.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@14286.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@14286.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@14286.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@14286.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@14286.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@14294.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@14294.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@14294.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@14294.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@14294.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@14350.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@14350.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@14350.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@14350.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@14350.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@14358.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@14358.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@14358.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@14358.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@14358.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@14366.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@14366.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@14366.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@14366.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@14366.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@14374.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@14374.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@14374.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@14374.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@14374.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@14382.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@14382.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@14382.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@14382.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@14382.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@14390.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@14390.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@14390.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@14390.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@14390.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@14398.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@14398.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@14398.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@14398.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@14398.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@14406.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@14406.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@14406.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@14406.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@14406.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@14414.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@14414.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@14414.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@14414.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@14414.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@14422.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@14422.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@14422.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@14422.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@14422.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@14430.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@14430.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@14430.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@14430.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@14430.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@14438.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@14438.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@14438.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@14438.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@14438.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@14494.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@14494.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@14494.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@14494.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@14494.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@14502.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@14502.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@14502.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@14502.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@14502.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@14510.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@14510.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@14510.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@14510.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@14510.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@14518.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@14518.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@14518.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@14518.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@14518.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@14526.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@14526.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@14526.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@14526.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@14526.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@14534.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@14534.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@14534.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@14534.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@14534.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@14542.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@14542.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@14542.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@14542.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@14542.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@14550.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@14550.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@14550.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@14550.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@14550.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@14558.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@14558.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@14558.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@14558.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@14558.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@14566.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@14566.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@14566.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@14566.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@14566.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@14574.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@14574.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@14574.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@14574.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@14574.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@14582.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@14582.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@14582.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@14582.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@14582.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@14638.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@14638.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@14638.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@14638.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@14638.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@14646.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@14646.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@14646.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@14646.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@14646.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@14654.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@14654.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@14654.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@14654.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@14654.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@14662.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@14662.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@14662.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@14662.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@14662.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@14670.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@14670.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@14670.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@14670.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@14670.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@14678.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@14678.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@14678.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@14678.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@14678.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@14686.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@14686.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@14686.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@14686.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@14686.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@14694.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@14694.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@14694.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@14694.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@14694.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@14702.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@14702.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@14702.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@14702.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@14702.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@14710.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@14710.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@14710.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@14710.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@14710.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@14718.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@14718.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@14718.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@14718.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@14718.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@14726.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@14726.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@14726.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@14726.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@14726.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@14782.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@14782.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@14782.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@14782.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@14782.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@14790.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@14790.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@14790.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@14790.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@14790.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@14798.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@14798.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@14798.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@14798.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@14798.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@14806.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@14806.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@14806.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@14806.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@14806.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@14814.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@14814.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@14814.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@14814.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@14814.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@14822.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@14822.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@14822.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@14822.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@14822.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@14830.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@14830.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@14830.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@14830.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@14830.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@14838.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@14838.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@14838.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@14838.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@14838.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@14846.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@14846.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@14846.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@14846.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@14846.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@14854.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@14854.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@14854.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@14854.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@14854.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@14870.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@14870.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@14870.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@14870.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@14870.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@14926.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@14926.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@14926.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@14926.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@14926.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@14934.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@14934.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@14934.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@14934.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@14934.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@14942.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@14942.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@14942.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@14942.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@14942.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@14950.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@14950.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@14950.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@14950.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@14950.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@14966.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@14966.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@14966.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@14966.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@14966.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@14974.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@14974.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@14974.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@14974.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@14974.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@14990.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@14990.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@14990.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@14990.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@14990.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@14998.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@14998.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@14998.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@14998.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@14998.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@15006.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@15006.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@15006.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@15006.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@15006.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@15014.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@15014.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@15014.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@15014.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@15014.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@15070.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@15070.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@15070.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@15070.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@15070.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@15078.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@15078.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@15078.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@15078.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@15078.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@15086.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@15086.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@15086.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@15086.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@15086.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@15094.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@15094.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@15094.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@15094.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@15094.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@15102.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@15102.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@15102.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@15102.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@15102.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@15110.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@15110.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@15110.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@15110.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@15110.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@15118.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@15118.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@15118.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@15118.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@15118.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@15126.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@15126.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@15126.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@15126.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@15126.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@15134.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@15134.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@15134.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@15134.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@15134.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@15142.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@15142.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@15142.4]
  wire  RetimeWrapper_105_io_in; // @[package.scala 93:22:@15142.4]
  wire  RetimeWrapper_105_io_out; // @[package.scala 93:22:@15142.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@15150.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@15150.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@15150.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@15150.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@15150.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@15158.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@15158.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@15158.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@15158.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@15158.4]
  wire  _T_316; // @[MemPrimitives.scala 82:210:@12669.4]
  wire  _T_318; // @[MemPrimitives.scala 82:210:@12670.4]
  wire  _T_319; // @[MemPrimitives.scala 82:228:@12671.4]
  wire  _T_320; // @[MemPrimitives.scala 83:102:@12672.4]
  wire [42:0] _T_322; // @[Cat.scala 30:58:@12674.4]
  wire  _T_329; // @[MemPrimitives.scala 82:210:@12682.4]
  wire  _T_330; // @[MemPrimitives.scala 82:228:@12683.4]
  wire  _T_331; // @[MemPrimitives.scala 83:102:@12684.4]
  wire [42:0] _T_333; // @[Cat.scala 30:58:@12686.4]
  wire  _T_340; // @[MemPrimitives.scala 82:210:@12694.4]
  wire  _T_341; // @[MemPrimitives.scala 82:228:@12695.4]
  wire  _T_342; // @[MemPrimitives.scala 83:102:@12696.4]
  wire [42:0] _T_344; // @[Cat.scala 30:58:@12698.4]
  wire  _T_349; // @[MemPrimitives.scala 82:210:@12705.4]
  wire  _T_352; // @[MemPrimitives.scala 82:228:@12707.4]
  wire  _T_353; // @[MemPrimitives.scala 83:102:@12708.4]
  wire [42:0] _T_355; // @[Cat.scala 30:58:@12710.4]
  wire  _T_363; // @[MemPrimitives.scala 82:228:@12719.4]
  wire  _T_364; // @[MemPrimitives.scala 83:102:@12720.4]
  wire [42:0] _T_366; // @[Cat.scala 30:58:@12722.4]
  wire  _T_374; // @[MemPrimitives.scala 82:228:@12731.4]
  wire  _T_375; // @[MemPrimitives.scala 83:102:@12732.4]
  wire [42:0] _T_377; // @[Cat.scala 30:58:@12734.4]
  wire  _T_382; // @[MemPrimitives.scala 82:210:@12741.4]
  wire  _T_385; // @[MemPrimitives.scala 82:228:@12743.4]
  wire  _T_386; // @[MemPrimitives.scala 83:102:@12744.4]
  wire [42:0] _T_388; // @[Cat.scala 30:58:@12746.4]
  wire  _T_396; // @[MemPrimitives.scala 82:228:@12755.4]
  wire  _T_397; // @[MemPrimitives.scala 83:102:@12756.4]
  wire [42:0] _T_399; // @[Cat.scala 30:58:@12758.4]
  wire  _T_407; // @[MemPrimitives.scala 82:228:@12767.4]
  wire  _T_408; // @[MemPrimitives.scala 83:102:@12768.4]
  wire [42:0] _T_410; // @[Cat.scala 30:58:@12770.4]
  wire  _T_415; // @[MemPrimitives.scala 82:210:@12777.4]
  wire  _T_418; // @[MemPrimitives.scala 82:228:@12779.4]
  wire  _T_419; // @[MemPrimitives.scala 83:102:@12780.4]
  wire [42:0] _T_421; // @[Cat.scala 30:58:@12782.4]
  wire  _T_429; // @[MemPrimitives.scala 82:228:@12791.4]
  wire  _T_430; // @[MemPrimitives.scala 83:102:@12792.4]
  wire [42:0] _T_432; // @[Cat.scala 30:58:@12794.4]
  wire  _T_440; // @[MemPrimitives.scala 82:228:@12803.4]
  wire  _T_441; // @[MemPrimitives.scala 83:102:@12804.4]
  wire [42:0] _T_443; // @[Cat.scala 30:58:@12806.4]
  wire  _T_448; // @[MemPrimitives.scala 110:210:@12813.4]
  wire  _T_450; // @[MemPrimitives.scala 110:210:@12814.4]
  wire  _T_451; // @[MemPrimitives.scala 110:228:@12815.4]
  wire  _T_454; // @[MemPrimitives.scala 110:210:@12817.4]
  wire  _T_456; // @[MemPrimitives.scala 110:210:@12818.4]
  wire  _T_457; // @[MemPrimitives.scala 110:228:@12819.4]
  wire  _T_460; // @[MemPrimitives.scala 110:210:@12821.4]
  wire  _T_462; // @[MemPrimitives.scala 110:210:@12822.4]
  wire  _T_463; // @[MemPrimitives.scala 110:228:@12823.4]
  wire  _T_466; // @[MemPrimitives.scala 110:210:@12825.4]
  wire  _T_468; // @[MemPrimitives.scala 110:210:@12826.4]
  wire  _T_469; // @[MemPrimitives.scala 110:228:@12827.4]
  wire  _T_472; // @[MemPrimitives.scala 110:210:@12829.4]
  wire  _T_474; // @[MemPrimitives.scala 110:210:@12830.4]
  wire  _T_475; // @[MemPrimitives.scala 110:228:@12831.4]
  wire  _T_478; // @[MemPrimitives.scala 110:210:@12833.4]
  wire  _T_480; // @[MemPrimitives.scala 110:210:@12834.4]
  wire  _T_481; // @[MemPrimitives.scala 110:228:@12835.4]
  wire  _T_484; // @[MemPrimitives.scala 110:210:@12837.4]
  wire  _T_486; // @[MemPrimitives.scala 110:210:@12838.4]
  wire  _T_487; // @[MemPrimitives.scala 110:228:@12839.4]
  wire  _T_490; // @[MemPrimitives.scala 110:210:@12841.4]
  wire  _T_492; // @[MemPrimitives.scala 110:210:@12842.4]
  wire  _T_493; // @[MemPrimitives.scala 110:228:@12843.4]
  wire  _T_496; // @[MemPrimitives.scala 110:210:@12845.4]
  wire  _T_498; // @[MemPrimitives.scala 110:210:@12846.4]
  wire  _T_499; // @[MemPrimitives.scala 110:228:@12847.4]
  wire  _T_501; // @[MemPrimitives.scala 126:35:@12861.4]
  wire  _T_502; // @[MemPrimitives.scala 126:35:@12862.4]
  wire  _T_503; // @[MemPrimitives.scala 126:35:@12863.4]
  wire  _T_504; // @[MemPrimitives.scala 126:35:@12864.4]
  wire  _T_505; // @[MemPrimitives.scala 126:35:@12865.4]
  wire  _T_506; // @[MemPrimitives.scala 126:35:@12866.4]
  wire  _T_507; // @[MemPrimitives.scala 126:35:@12867.4]
  wire  _T_508; // @[MemPrimitives.scala 126:35:@12868.4]
  wire  _T_509; // @[MemPrimitives.scala 126:35:@12869.4]
  wire [11:0] _T_511; // @[Cat.scala 30:58:@12871.4]
  wire [11:0] _T_513; // @[Cat.scala 30:58:@12873.4]
  wire [11:0] _T_515; // @[Cat.scala 30:58:@12875.4]
  wire [11:0] _T_517; // @[Cat.scala 30:58:@12877.4]
  wire [11:0] _T_519; // @[Cat.scala 30:58:@12879.4]
  wire [11:0] _T_521; // @[Cat.scala 30:58:@12881.4]
  wire [11:0] _T_523; // @[Cat.scala 30:58:@12883.4]
  wire [11:0] _T_525; // @[Cat.scala 30:58:@12885.4]
  wire [11:0] _T_527; // @[Cat.scala 30:58:@12887.4]
  wire [11:0] _T_528; // @[Mux.scala 31:69:@12888.4]
  wire [11:0] _T_529; // @[Mux.scala 31:69:@12889.4]
  wire [11:0] _T_530; // @[Mux.scala 31:69:@12890.4]
  wire [11:0] _T_531; // @[Mux.scala 31:69:@12891.4]
  wire [11:0] _T_532; // @[Mux.scala 31:69:@12892.4]
  wire [11:0] _T_533; // @[Mux.scala 31:69:@12893.4]
  wire [11:0] _T_534; // @[Mux.scala 31:69:@12894.4]
  wire [11:0] _T_535; // @[Mux.scala 31:69:@12895.4]
  wire  _T_542; // @[MemPrimitives.scala 110:210:@12903.4]
  wire  _T_543; // @[MemPrimitives.scala 110:228:@12904.4]
  wire  _T_548; // @[MemPrimitives.scala 110:210:@12907.4]
  wire  _T_549; // @[MemPrimitives.scala 110:228:@12908.4]
  wire  _T_554; // @[MemPrimitives.scala 110:210:@12911.4]
  wire  _T_555; // @[MemPrimitives.scala 110:228:@12912.4]
  wire  _T_560; // @[MemPrimitives.scala 110:210:@12915.4]
  wire  _T_561; // @[MemPrimitives.scala 110:228:@12916.4]
  wire  _T_566; // @[MemPrimitives.scala 110:210:@12919.4]
  wire  _T_567; // @[MemPrimitives.scala 110:228:@12920.4]
  wire  _T_572; // @[MemPrimitives.scala 110:210:@12923.4]
  wire  _T_573; // @[MemPrimitives.scala 110:228:@12924.4]
  wire  _T_578; // @[MemPrimitives.scala 110:210:@12927.4]
  wire  _T_579; // @[MemPrimitives.scala 110:228:@12928.4]
  wire  _T_584; // @[MemPrimitives.scala 110:210:@12931.4]
  wire  _T_585; // @[MemPrimitives.scala 110:228:@12932.4]
  wire  _T_590; // @[MemPrimitives.scala 110:210:@12935.4]
  wire  _T_591; // @[MemPrimitives.scala 110:228:@12936.4]
  wire  _T_593; // @[MemPrimitives.scala 126:35:@12950.4]
  wire  _T_594; // @[MemPrimitives.scala 126:35:@12951.4]
  wire  _T_595; // @[MemPrimitives.scala 126:35:@12952.4]
  wire  _T_596; // @[MemPrimitives.scala 126:35:@12953.4]
  wire  _T_597; // @[MemPrimitives.scala 126:35:@12954.4]
  wire  _T_598; // @[MemPrimitives.scala 126:35:@12955.4]
  wire  _T_599; // @[MemPrimitives.scala 126:35:@12956.4]
  wire  _T_600; // @[MemPrimitives.scala 126:35:@12957.4]
  wire  _T_601; // @[MemPrimitives.scala 126:35:@12958.4]
  wire [11:0] _T_603; // @[Cat.scala 30:58:@12960.4]
  wire [11:0] _T_605; // @[Cat.scala 30:58:@12962.4]
  wire [11:0] _T_607; // @[Cat.scala 30:58:@12964.4]
  wire [11:0] _T_609; // @[Cat.scala 30:58:@12966.4]
  wire [11:0] _T_611; // @[Cat.scala 30:58:@12968.4]
  wire [11:0] _T_613; // @[Cat.scala 30:58:@12970.4]
  wire [11:0] _T_615; // @[Cat.scala 30:58:@12972.4]
  wire [11:0] _T_617; // @[Cat.scala 30:58:@12974.4]
  wire [11:0] _T_619; // @[Cat.scala 30:58:@12976.4]
  wire [11:0] _T_620; // @[Mux.scala 31:69:@12977.4]
  wire [11:0] _T_621; // @[Mux.scala 31:69:@12978.4]
  wire [11:0] _T_622; // @[Mux.scala 31:69:@12979.4]
  wire [11:0] _T_623; // @[Mux.scala 31:69:@12980.4]
  wire [11:0] _T_624; // @[Mux.scala 31:69:@12981.4]
  wire [11:0] _T_625; // @[Mux.scala 31:69:@12982.4]
  wire [11:0] _T_626; // @[Mux.scala 31:69:@12983.4]
  wire [11:0] _T_627; // @[Mux.scala 31:69:@12984.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@12992.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@12993.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@12996.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@12997.4]
  wire  _T_646; // @[MemPrimitives.scala 110:210:@13000.4]
  wire  _T_647; // @[MemPrimitives.scala 110:228:@13001.4]
  wire  _T_652; // @[MemPrimitives.scala 110:210:@13004.4]
  wire  _T_653; // @[MemPrimitives.scala 110:228:@13005.4]
  wire  _T_658; // @[MemPrimitives.scala 110:210:@13008.4]
  wire  _T_659; // @[MemPrimitives.scala 110:228:@13009.4]
  wire  _T_664; // @[MemPrimitives.scala 110:210:@13012.4]
  wire  _T_665; // @[MemPrimitives.scala 110:228:@13013.4]
  wire  _T_670; // @[MemPrimitives.scala 110:210:@13016.4]
  wire  _T_671; // @[MemPrimitives.scala 110:228:@13017.4]
  wire  _T_676; // @[MemPrimitives.scala 110:210:@13020.4]
  wire  _T_677; // @[MemPrimitives.scala 110:228:@13021.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@13024.4]
  wire  _T_683; // @[MemPrimitives.scala 110:228:@13025.4]
  wire  _T_685; // @[MemPrimitives.scala 126:35:@13039.4]
  wire  _T_686; // @[MemPrimitives.scala 126:35:@13040.4]
  wire  _T_687; // @[MemPrimitives.scala 126:35:@13041.4]
  wire  _T_688; // @[MemPrimitives.scala 126:35:@13042.4]
  wire  _T_689; // @[MemPrimitives.scala 126:35:@13043.4]
  wire  _T_690; // @[MemPrimitives.scala 126:35:@13044.4]
  wire  _T_691; // @[MemPrimitives.scala 126:35:@13045.4]
  wire  _T_692; // @[MemPrimitives.scala 126:35:@13046.4]
  wire  _T_693; // @[MemPrimitives.scala 126:35:@13047.4]
  wire [11:0] _T_695; // @[Cat.scala 30:58:@13049.4]
  wire [11:0] _T_697; // @[Cat.scala 30:58:@13051.4]
  wire [11:0] _T_699; // @[Cat.scala 30:58:@13053.4]
  wire [11:0] _T_701; // @[Cat.scala 30:58:@13055.4]
  wire [11:0] _T_703; // @[Cat.scala 30:58:@13057.4]
  wire [11:0] _T_705; // @[Cat.scala 30:58:@13059.4]
  wire [11:0] _T_707; // @[Cat.scala 30:58:@13061.4]
  wire [11:0] _T_709; // @[Cat.scala 30:58:@13063.4]
  wire [11:0] _T_711; // @[Cat.scala 30:58:@13065.4]
  wire [11:0] _T_712; // @[Mux.scala 31:69:@13066.4]
  wire [11:0] _T_713; // @[Mux.scala 31:69:@13067.4]
  wire [11:0] _T_714; // @[Mux.scala 31:69:@13068.4]
  wire [11:0] _T_715; // @[Mux.scala 31:69:@13069.4]
  wire [11:0] _T_716; // @[Mux.scala 31:69:@13070.4]
  wire [11:0] _T_717; // @[Mux.scala 31:69:@13071.4]
  wire [11:0] _T_718; // @[Mux.scala 31:69:@13072.4]
  wire [11:0] _T_719; // @[Mux.scala 31:69:@13073.4]
  wire  _T_724; // @[MemPrimitives.scala 110:210:@13080.4]
  wire  _T_727; // @[MemPrimitives.scala 110:228:@13082.4]
  wire  _T_730; // @[MemPrimitives.scala 110:210:@13084.4]
  wire  _T_733; // @[MemPrimitives.scala 110:228:@13086.4]
  wire  _T_736; // @[MemPrimitives.scala 110:210:@13088.4]
  wire  _T_739; // @[MemPrimitives.scala 110:228:@13090.4]
  wire  _T_742; // @[MemPrimitives.scala 110:210:@13092.4]
  wire  _T_745; // @[MemPrimitives.scala 110:228:@13094.4]
  wire  _T_748; // @[MemPrimitives.scala 110:210:@13096.4]
  wire  _T_751; // @[MemPrimitives.scala 110:228:@13098.4]
  wire  _T_754; // @[MemPrimitives.scala 110:210:@13100.4]
  wire  _T_757; // @[MemPrimitives.scala 110:228:@13102.4]
  wire  _T_760; // @[MemPrimitives.scala 110:210:@13104.4]
  wire  _T_763; // @[MemPrimitives.scala 110:228:@13106.4]
  wire  _T_766; // @[MemPrimitives.scala 110:210:@13108.4]
  wire  _T_769; // @[MemPrimitives.scala 110:228:@13110.4]
  wire  _T_772; // @[MemPrimitives.scala 110:210:@13112.4]
  wire  _T_775; // @[MemPrimitives.scala 110:228:@13114.4]
  wire  _T_777; // @[MemPrimitives.scala 126:35:@13128.4]
  wire  _T_778; // @[MemPrimitives.scala 126:35:@13129.4]
  wire  _T_779; // @[MemPrimitives.scala 126:35:@13130.4]
  wire  _T_780; // @[MemPrimitives.scala 126:35:@13131.4]
  wire  _T_781; // @[MemPrimitives.scala 126:35:@13132.4]
  wire  _T_782; // @[MemPrimitives.scala 126:35:@13133.4]
  wire  _T_783; // @[MemPrimitives.scala 126:35:@13134.4]
  wire  _T_784; // @[MemPrimitives.scala 126:35:@13135.4]
  wire  _T_785; // @[MemPrimitives.scala 126:35:@13136.4]
  wire [11:0] _T_787; // @[Cat.scala 30:58:@13138.4]
  wire [11:0] _T_789; // @[Cat.scala 30:58:@13140.4]
  wire [11:0] _T_791; // @[Cat.scala 30:58:@13142.4]
  wire [11:0] _T_793; // @[Cat.scala 30:58:@13144.4]
  wire [11:0] _T_795; // @[Cat.scala 30:58:@13146.4]
  wire [11:0] _T_797; // @[Cat.scala 30:58:@13148.4]
  wire [11:0] _T_799; // @[Cat.scala 30:58:@13150.4]
  wire [11:0] _T_801; // @[Cat.scala 30:58:@13152.4]
  wire [11:0] _T_803; // @[Cat.scala 30:58:@13154.4]
  wire [11:0] _T_804; // @[Mux.scala 31:69:@13155.4]
  wire [11:0] _T_805; // @[Mux.scala 31:69:@13156.4]
  wire [11:0] _T_806; // @[Mux.scala 31:69:@13157.4]
  wire [11:0] _T_807; // @[Mux.scala 31:69:@13158.4]
  wire [11:0] _T_808; // @[Mux.scala 31:69:@13159.4]
  wire [11:0] _T_809; // @[Mux.scala 31:69:@13160.4]
  wire [11:0] _T_810; // @[Mux.scala 31:69:@13161.4]
  wire [11:0] _T_811; // @[Mux.scala 31:69:@13162.4]
  wire  _T_819; // @[MemPrimitives.scala 110:228:@13171.4]
  wire  _T_825; // @[MemPrimitives.scala 110:228:@13175.4]
  wire  _T_831; // @[MemPrimitives.scala 110:228:@13179.4]
  wire  _T_837; // @[MemPrimitives.scala 110:228:@13183.4]
  wire  _T_843; // @[MemPrimitives.scala 110:228:@13187.4]
  wire  _T_849; // @[MemPrimitives.scala 110:228:@13191.4]
  wire  _T_855; // @[MemPrimitives.scala 110:228:@13195.4]
  wire  _T_861; // @[MemPrimitives.scala 110:228:@13199.4]
  wire  _T_867; // @[MemPrimitives.scala 110:228:@13203.4]
  wire  _T_869; // @[MemPrimitives.scala 126:35:@13217.4]
  wire  _T_870; // @[MemPrimitives.scala 126:35:@13218.4]
  wire  _T_871; // @[MemPrimitives.scala 126:35:@13219.4]
  wire  _T_872; // @[MemPrimitives.scala 126:35:@13220.4]
  wire  _T_873; // @[MemPrimitives.scala 126:35:@13221.4]
  wire  _T_874; // @[MemPrimitives.scala 126:35:@13222.4]
  wire  _T_875; // @[MemPrimitives.scala 126:35:@13223.4]
  wire  _T_876; // @[MemPrimitives.scala 126:35:@13224.4]
  wire  _T_877; // @[MemPrimitives.scala 126:35:@13225.4]
  wire [11:0] _T_879; // @[Cat.scala 30:58:@13227.4]
  wire [11:0] _T_881; // @[Cat.scala 30:58:@13229.4]
  wire [11:0] _T_883; // @[Cat.scala 30:58:@13231.4]
  wire [11:0] _T_885; // @[Cat.scala 30:58:@13233.4]
  wire [11:0] _T_887; // @[Cat.scala 30:58:@13235.4]
  wire [11:0] _T_889; // @[Cat.scala 30:58:@13237.4]
  wire [11:0] _T_891; // @[Cat.scala 30:58:@13239.4]
  wire [11:0] _T_893; // @[Cat.scala 30:58:@13241.4]
  wire [11:0] _T_895; // @[Cat.scala 30:58:@13243.4]
  wire [11:0] _T_896; // @[Mux.scala 31:69:@13244.4]
  wire [11:0] _T_897; // @[Mux.scala 31:69:@13245.4]
  wire [11:0] _T_898; // @[Mux.scala 31:69:@13246.4]
  wire [11:0] _T_899; // @[Mux.scala 31:69:@13247.4]
  wire [11:0] _T_900; // @[Mux.scala 31:69:@13248.4]
  wire [11:0] _T_901; // @[Mux.scala 31:69:@13249.4]
  wire [11:0] _T_902; // @[Mux.scala 31:69:@13250.4]
  wire [11:0] _T_903; // @[Mux.scala 31:69:@13251.4]
  wire  _T_911; // @[MemPrimitives.scala 110:228:@13260.4]
  wire  _T_917; // @[MemPrimitives.scala 110:228:@13264.4]
  wire  _T_923; // @[MemPrimitives.scala 110:228:@13268.4]
  wire  _T_929; // @[MemPrimitives.scala 110:228:@13272.4]
  wire  _T_935; // @[MemPrimitives.scala 110:228:@13276.4]
  wire  _T_941; // @[MemPrimitives.scala 110:228:@13280.4]
  wire  _T_947; // @[MemPrimitives.scala 110:228:@13284.4]
  wire  _T_953; // @[MemPrimitives.scala 110:228:@13288.4]
  wire  _T_959; // @[MemPrimitives.scala 110:228:@13292.4]
  wire  _T_961; // @[MemPrimitives.scala 126:35:@13306.4]
  wire  _T_962; // @[MemPrimitives.scala 126:35:@13307.4]
  wire  _T_963; // @[MemPrimitives.scala 126:35:@13308.4]
  wire  _T_964; // @[MemPrimitives.scala 126:35:@13309.4]
  wire  _T_965; // @[MemPrimitives.scala 126:35:@13310.4]
  wire  _T_966; // @[MemPrimitives.scala 126:35:@13311.4]
  wire  _T_967; // @[MemPrimitives.scala 126:35:@13312.4]
  wire  _T_968; // @[MemPrimitives.scala 126:35:@13313.4]
  wire  _T_969; // @[MemPrimitives.scala 126:35:@13314.4]
  wire [11:0] _T_971; // @[Cat.scala 30:58:@13316.4]
  wire [11:0] _T_973; // @[Cat.scala 30:58:@13318.4]
  wire [11:0] _T_975; // @[Cat.scala 30:58:@13320.4]
  wire [11:0] _T_977; // @[Cat.scala 30:58:@13322.4]
  wire [11:0] _T_979; // @[Cat.scala 30:58:@13324.4]
  wire [11:0] _T_981; // @[Cat.scala 30:58:@13326.4]
  wire [11:0] _T_983; // @[Cat.scala 30:58:@13328.4]
  wire [11:0] _T_985; // @[Cat.scala 30:58:@13330.4]
  wire [11:0] _T_987; // @[Cat.scala 30:58:@13332.4]
  wire [11:0] _T_988; // @[Mux.scala 31:69:@13333.4]
  wire [11:0] _T_989; // @[Mux.scala 31:69:@13334.4]
  wire [11:0] _T_990; // @[Mux.scala 31:69:@13335.4]
  wire [11:0] _T_991; // @[Mux.scala 31:69:@13336.4]
  wire [11:0] _T_992; // @[Mux.scala 31:69:@13337.4]
  wire [11:0] _T_993; // @[Mux.scala 31:69:@13338.4]
  wire [11:0] _T_994; // @[Mux.scala 31:69:@13339.4]
  wire [11:0] _T_995; // @[Mux.scala 31:69:@13340.4]
  wire  _T_1000; // @[MemPrimitives.scala 110:210:@13347.4]
  wire  _T_1003; // @[MemPrimitives.scala 110:228:@13349.4]
  wire  _T_1006; // @[MemPrimitives.scala 110:210:@13351.4]
  wire  _T_1009; // @[MemPrimitives.scala 110:228:@13353.4]
  wire  _T_1012; // @[MemPrimitives.scala 110:210:@13355.4]
  wire  _T_1015; // @[MemPrimitives.scala 110:228:@13357.4]
  wire  _T_1018; // @[MemPrimitives.scala 110:210:@13359.4]
  wire  _T_1021; // @[MemPrimitives.scala 110:228:@13361.4]
  wire  _T_1024; // @[MemPrimitives.scala 110:210:@13363.4]
  wire  _T_1027; // @[MemPrimitives.scala 110:228:@13365.4]
  wire  _T_1030; // @[MemPrimitives.scala 110:210:@13367.4]
  wire  _T_1033; // @[MemPrimitives.scala 110:228:@13369.4]
  wire  _T_1036; // @[MemPrimitives.scala 110:210:@13371.4]
  wire  _T_1039; // @[MemPrimitives.scala 110:228:@13373.4]
  wire  _T_1042; // @[MemPrimitives.scala 110:210:@13375.4]
  wire  _T_1045; // @[MemPrimitives.scala 110:228:@13377.4]
  wire  _T_1048; // @[MemPrimitives.scala 110:210:@13379.4]
  wire  _T_1051; // @[MemPrimitives.scala 110:228:@13381.4]
  wire  _T_1053; // @[MemPrimitives.scala 126:35:@13395.4]
  wire  _T_1054; // @[MemPrimitives.scala 126:35:@13396.4]
  wire  _T_1055; // @[MemPrimitives.scala 126:35:@13397.4]
  wire  _T_1056; // @[MemPrimitives.scala 126:35:@13398.4]
  wire  _T_1057; // @[MemPrimitives.scala 126:35:@13399.4]
  wire  _T_1058; // @[MemPrimitives.scala 126:35:@13400.4]
  wire  _T_1059; // @[MemPrimitives.scala 126:35:@13401.4]
  wire  _T_1060; // @[MemPrimitives.scala 126:35:@13402.4]
  wire  _T_1061; // @[MemPrimitives.scala 126:35:@13403.4]
  wire [11:0] _T_1063; // @[Cat.scala 30:58:@13405.4]
  wire [11:0] _T_1065; // @[Cat.scala 30:58:@13407.4]
  wire [11:0] _T_1067; // @[Cat.scala 30:58:@13409.4]
  wire [11:0] _T_1069; // @[Cat.scala 30:58:@13411.4]
  wire [11:0] _T_1071; // @[Cat.scala 30:58:@13413.4]
  wire [11:0] _T_1073; // @[Cat.scala 30:58:@13415.4]
  wire [11:0] _T_1075; // @[Cat.scala 30:58:@13417.4]
  wire [11:0] _T_1077; // @[Cat.scala 30:58:@13419.4]
  wire [11:0] _T_1079; // @[Cat.scala 30:58:@13421.4]
  wire [11:0] _T_1080; // @[Mux.scala 31:69:@13422.4]
  wire [11:0] _T_1081; // @[Mux.scala 31:69:@13423.4]
  wire [11:0] _T_1082; // @[Mux.scala 31:69:@13424.4]
  wire [11:0] _T_1083; // @[Mux.scala 31:69:@13425.4]
  wire [11:0] _T_1084; // @[Mux.scala 31:69:@13426.4]
  wire [11:0] _T_1085; // @[Mux.scala 31:69:@13427.4]
  wire [11:0] _T_1086; // @[Mux.scala 31:69:@13428.4]
  wire [11:0] _T_1087; // @[Mux.scala 31:69:@13429.4]
  wire  _T_1095; // @[MemPrimitives.scala 110:228:@13438.4]
  wire  _T_1101; // @[MemPrimitives.scala 110:228:@13442.4]
  wire  _T_1107; // @[MemPrimitives.scala 110:228:@13446.4]
  wire  _T_1113; // @[MemPrimitives.scala 110:228:@13450.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@13454.4]
  wire  _T_1125; // @[MemPrimitives.scala 110:228:@13458.4]
  wire  _T_1131; // @[MemPrimitives.scala 110:228:@13462.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:228:@13466.4]
  wire  _T_1143; // @[MemPrimitives.scala 110:228:@13470.4]
  wire  _T_1145; // @[MemPrimitives.scala 126:35:@13484.4]
  wire  _T_1146; // @[MemPrimitives.scala 126:35:@13485.4]
  wire  _T_1147; // @[MemPrimitives.scala 126:35:@13486.4]
  wire  _T_1148; // @[MemPrimitives.scala 126:35:@13487.4]
  wire  _T_1149; // @[MemPrimitives.scala 126:35:@13488.4]
  wire  _T_1150; // @[MemPrimitives.scala 126:35:@13489.4]
  wire  _T_1151; // @[MemPrimitives.scala 126:35:@13490.4]
  wire  _T_1152; // @[MemPrimitives.scala 126:35:@13491.4]
  wire  _T_1153; // @[MemPrimitives.scala 126:35:@13492.4]
  wire [11:0] _T_1155; // @[Cat.scala 30:58:@13494.4]
  wire [11:0] _T_1157; // @[Cat.scala 30:58:@13496.4]
  wire [11:0] _T_1159; // @[Cat.scala 30:58:@13498.4]
  wire [11:0] _T_1161; // @[Cat.scala 30:58:@13500.4]
  wire [11:0] _T_1163; // @[Cat.scala 30:58:@13502.4]
  wire [11:0] _T_1165; // @[Cat.scala 30:58:@13504.4]
  wire [11:0] _T_1167; // @[Cat.scala 30:58:@13506.4]
  wire [11:0] _T_1169; // @[Cat.scala 30:58:@13508.4]
  wire [11:0] _T_1171; // @[Cat.scala 30:58:@13510.4]
  wire [11:0] _T_1172; // @[Mux.scala 31:69:@13511.4]
  wire [11:0] _T_1173; // @[Mux.scala 31:69:@13512.4]
  wire [11:0] _T_1174; // @[Mux.scala 31:69:@13513.4]
  wire [11:0] _T_1175; // @[Mux.scala 31:69:@13514.4]
  wire [11:0] _T_1176; // @[Mux.scala 31:69:@13515.4]
  wire [11:0] _T_1177; // @[Mux.scala 31:69:@13516.4]
  wire [11:0] _T_1178; // @[Mux.scala 31:69:@13517.4]
  wire [11:0] _T_1179; // @[Mux.scala 31:69:@13518.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@13527.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@13531.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@13535.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@13539.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@13543.4]
  wire  _T_1217; // @[MemPrimitives.scala 110:228:@13547.4]
  wire  _T_1223; // @[MemPrimitives.scala 110:228:@13551.4]
  wire  _T_1229; // @[MemPrimitives.scala 110:228:@13555.4]
  wire  _T_1235; // @[MemPrimitives.scala 110:228:@13559.4]
  wire  _T_1237; // @[MemPrimitives.scala 126:35:@13573.4]
  wire  _T_1238; // @[MemPrimitives.scala 126:35:@13574.4]
  wire  _T_1239; // @[MemPrimitives.scala 126:35:@13575.4]
  wire  _T_1240; // @[MemPrimitives.scala 126:35:@13576.4]
  wire  _T_1241; // @[MemPrimitives.scala 126:35:@13577.4]
  wire  _T_1242; // @[MemPrimitives.scala 126:35:@13578.4]
  wire  _T_1243; // @[MemPrimitives.scala 126:35:@13579.4]
  wire  _T_1244; // @[MemPrimitives.scala 126:35:@13580.4]
  wire  _T_1245; // @[MemPrimitives.scala 126:35:@13581.4]
  wire [11:0] _T_1247; // @[Cat.scala 30:58:@13583.4]
  wire [11:0] _T_1249; // @[Cat.scala 30:58:@13585.4]
  wire [11:0] _T_1251; // @[Cat.scala 30:58:@13587.4]
  wire [11:0] _T_1253; // @[Cat.scala 30:58:@13589.4]
  wire [11:0] _T_1255; // @[Cat.scala 30:58:@13591.4]
  wire [11:0] _T_1257; // @[Cat.scala 30:58:@13593.4]
  wire [11:0] _T_1259; // @[Cat.scala 30:58:@13595.4]
  wire [11:0] _T_1261; // @[Cat.scala 30:58:@13597.4]
  wire [11:0] _T_1263; // @[Cat.scala 30:58:@13599.4]
  wire [11:0] _T_1264; // @[Mux.scala 31:69:@13600.4]
  wire [11:0] _T_1265; // @[Mux.scala 31:69:@13601.4]
  wire [11:0] _T_1266; // @[Mux.scala 31:69:@13602.4]
  wire [11:0] _T_1267; // @[Mux.scala 31:69:@13603.4]
  wire [11:0] _T_1268; // @[Mux.scala 31:69:@13604.4]
  wire [11:0] _T_1269; // @[Mux.scala 31:69:@13605.4]
  wire [11:0] _T_1270; // @[Mux.scala 31:69:@13606.4]
  wire [11:0] _T_1271; // @[Mux.scala 31:69:@13607.4]
  wire  _T_1276; // @[MemPrimitives.scala 110:210:@13614.4]
  wire  _T_1279; // @[MemPrimitives.scala 110:228:@13616.4]
  wire  _T_1282; // @[MemPrimitives.scala 110:210:@13618.4]
  wire  _T_1285; // @[MemPrimitives.scala 110:228:@13620.4]
  wire  _T_1288; // @[MemPrimitives.scala 110:210:@13622.4]
  wire  _T_1291; // @[MemPrimitives.scala 110:228:@13624.4]
  wire  _T_1294; // @[MemPrimitives.scala 110:210:@13626.4]
  wire  _T_1297; // @[MemPrimitives.scala 110:228:@13628.4]
  wire  _T_1300; // @[MemPrimitives.scala 110:210:@13630.4]
  wire  _T_1303; // @[MemPrimitives.scala 110:228:@13632.4]
  wire  _T_1306; // @[MemPrimitives.scala 110:210:@13634.4]
  wire  _T_1309; // @[MemPrimitives.scala 110:228:@13636.4]
  wire  _T_1312; // @[MemPrimitives.scala 110:210:@13638.4]
  wire  _T_1315; // @[MemPrimitives.scala 110:228:@13640.4]
  wire  _T_1318; // @[MemPrimitives.scala 110:210:@13642.4]
  wire  _T_1321; // @[MemPrimitives.scala 110:228:@13644.4]
  wire  _T_1324; // @[MemPrimitives.scala 110:210:@13646.4]
  wire  _T_1327; // @[MemPrimitives.scala 110:228:@13648.4]
  wire  _T_1329; // @[MemPrimitives.scala 126:35:@13662.4]
  wire  _T_1330; // @[MemPrimitives.scala 126:35:@13663.4]
  wire  _T_1331; // @[MemPrimitives.scala 126:35:@13664.4]
  wire  _T_1332; // @[MemPrimitives.scala 126:35:@13665.4]
  wire  _T_1333; // @[MemPrimitives.scala 126:35:@13666.4]
  wire  _T_1334; // @[MemPrimitives.scala 126:35:@13667.4]
  wire  _T_1335; // @[MemPrimitives.scala 126:35:@13668.4]
  wire  _T_1336; // @[MemPrimitives.scala 126:35:@13669.4]
  wire  _T_1337; // @[MemPrimitives.scala 126:35:@13670.4]
  wire [11:0] _T_1339; // @[Cat.scala 30:58:@13672.4]
  wire [11:0] _T_1341; // @[Cat.scala 30:58:@13674.4]
  wire [11:0] _T_1343; // @[Cat.scala 30:58:@13676.4]
  wire [11:0] _T_1345; // @[Cat.scala 30:58:@13678.4]
  wire [11:0] _T_1347; // @[Cat.scala 30:58:@13680.4]
  wire [11:0] _T_1349; // @[Cat.scala 30:58:@13682.4]
  wire [11:0] _T_1351; // @[Cat.scala 30:58:@13684.4]
  wire [11:0] _T_1353; // @[Cat.scala 30:58:@13686.4]
  wire [11:0] _T_1355; // @[Cat.scala 30:58:@13688.4]
  wire [11:0] _T_1356; // @[Mux.scala 31:69:@13689.4]
  wire [11:0] _T_1357; // @[Mux.scala 31:69:@13690.4]
  wire [11:0] _T_1358; // @[Mux.scala 31:69:@13691.4]
  wire [11:0] _T_1359; // @[Mux.scala 31:69:@13692.4]
  wire [11:0] _T_1360; // @[Mux.scala 31:69:@13693.4]
  wire [11:0] _T_1361; // @[Mux.scala 31:69:@13694.4]
  wire [11:0] _T_1362; // @[Mux.scala 31:69:@13695.4]
  wire [11:0] _T_1363; // @[Mux.scala 31:69:@13696.4]
  wire  _T_1371; // @[MemPrimitives.scala 110:228:@13705.4]
  wire  _T_1377; // @[MemPrimitives.scala 110:228:@13709.4]
  wire  _T_1383; // @[MemPrimitives.scala 110:228:@13713.4]
  wire  _T_1389; // @[MemPrimitives.scala 110:228:@13717.4]
  wire  _T_1395; // @[MemPrimitives.scala 110:228:@13721.4]
  wire  _T_1401; // @[MemPrimitives.scala 110:228:@13725.4]
  wire  _T_1407; // @[MemPrimitives.scala 110:228:@13729.4]
  wire  _T_1413; // @[MemPrimitives.scala 110:228:@13733.4]
  wire  _T_1419; // @[MemPrimitives.scala 110:228:@13737.4]
  wire  _T_1421; // @[MemPrimitives.scala 126:35:@13751.4]
  wire  _T_1422; // @[MemPrimitives.scala 126:35:@13752.4]
  wire  _T_1423; // @[MemPrimitives.scala 126:35:@13753.4]
  wire  _T_1424; // @[MemPrimitives.scala 126:35:@13754.4]
  wire  _T_1425; // @[MemPrimitives.scala 126:35:@13755.4]
  wire  _T_1426; // @[MemPrimitives.scala 126:35:@13756.4]
  wire  _T_1427; // @[MemPrimitives.scala 126:35:@13757.4]
  wire  _T_1428; // @[MemPrimitives.scala 126:35:@13758.4]
  wire  _T_1429; // @[MemPrimitives.scala 126:35:@13759.4]
  wire [11:0] _T_1431; // @[Cat.scala 30:58:@13761.4]
  wire [11:0] _T_1433; // @[Cat.scala 30:58:@13763.4]
  wire [11:0] _T_1435; // @[Cat.scala 30:58:@13765.4]
  wire [11:0] _T_1437; // @[Cat.scala 30:58:@13767.4]
  wire [11:0] _T_1439; // @[Cat.scala 30:58:@13769.4]
  wire [11:0] _T_1441; // @[Cat.scala 30:58:@13771.4]
  wire [11:0] _T_1443; // @[Cat.scala 30:58:@13773.4]
  wire [11:0] _T_1445; // @[Cat.scala 30:58:@13775.4]
  wire [11:0] _T_1447; // @[Cat.scala 30:58:@13777.4]
  wire [11:0] _T_1448; // @[Mux.scala 31:69:@13778.4]
  wire [11:0] _T_1449; // @[Mux.scala 31:69:@13779.4]
  wire [11:0] _T_1450; // @[Mux.scala 31:69:@13780.4]
  wire [11:0] _T_1451; // @[Mux.scala 31:69:@13781.4]
  wire [11:0] _T_1452; // @[Mux.scala 31:69:@13782.4]
  wire [11:0] _T_1453; // @[Mux.scala 31:69:@13783.4]
  wire [11:0] _T_1454; // @[Mux.scala 31:69:@13784.4]
  wire [11:0] _T_1455; // @[Mux.scala 31:69:@13785.4]
  wire  _T_1463; // @[MemPrimitives.scala 110:228:@13794.4]
  wire  _T_1469; // @[MemPrimitives.scala 110:228:@13798.4]
  wire  _T_1475; // @[MemPrimitives.scala 110:228:@13802.4]
  wire  _T_1481; // @[MemPrimitives.scala 110:228:@13806.4]
  wire  _T_1487; // @[MemPrimitives.scala 110:228:@13810.4]
  wire  _T_1493; // @[MemPrimitives.scala 110:228:@13814.4]
  wire  _T_1499; // @[MemPrimitives.scala 110:228:@13818.4]
  wire  _T_1505; // @[MemPrimitives.scala 110:228:@13822.4]
  wire  _T_1511; // @[MemPrimitives.scala 110:228:@13826.4]
  wire  _T_1513; // @[MemPrimitives.scala 126:35:@13840.4]
  wire  _T_1514; // @[MemPrimitives.scala 126:35:@13841.4]
  wire  _T_1515; // @[MemPrimitives.scala 126:35:@13842.4]
  wire  _T_1516; // @[MemPrimitives.scala 126:35:@13843.4]
  wire  _T_1517; // @[MemPrimitives.scala 126:35:@13844.4]
  wire  _T_1518; // @[MemPrimitives.scala 126:35:@13845.4]
  wire  _T_1519; // @[MemPrimitives.scala 126:35:@13846.4]
  wire  _T_1520; // @[MemPrimitives.scala 126:35:@13847.4]
  wire  _T_1521; // @[MemPrimitives.scala 126:35:@13848.4]
  wire [11:0] _T_1523; // @[Cat.scala 30:58:@13850.4]
  wire [11:0] _T_1525; // @[Cat.scala 30:58:@13852.4]
  wire [11:0] _T_1527; // @[Cat.scala 30:58:@13854.4]
  wire [11:0] _T_1529; // @[Cat.scala 30:58:@13856.4]
  wire [11:0] _T_1531; // @[Cat.scala 30:58:@13858.4]
  wire [11:0] _T_1533; // @[Cat.scala 30:58:@13860.4]
  wire [11:0] _T_1535; // @[Cat.scala 30:58:@13862.4]
  wire [11:0] _T_1537; // @[Cat.scala 30:58:@13864.4]
  wire [11:0] _T_1539; // @[Cat.scala 30:58:@13866.4]
  wire [11:0] _T_1540; // @[Mux.scala 31:69:@13867.4]
  wire [11:0] _T_1541; // @[Mux.scala 31:69:@13868.4]
  wire [11:0] _T_1542; // @[Mux.scala 31:69:@13869.4]
  wire [11:0] _T_1543; // @[Mux.scala 31:69:@13870.4]
  wire [11:0] _T_1544; // @[Mux.scala 31:69:@13871.4]
  wire [11:0] _T_1545; // @[Mux.scala 31:69:@13872.4]
  wire [11:0] _T_1546; // @[Mux.scala 31:69:@13873.4]
  wire [11:0] _T_1547; // @[Mux.scala 31:69:@13874.4]
  wire  _T_1643; // @[package.scala 96:25:@14003.4 package.scala 96:25:@14004.4]
  wire [31:0] _T_1647; // @[Mux.scala 31:69:@14013.4]
  wire  _T_1640; // @[package.scala 96:25:@13995.4 package.scala 96:25:@13996.4]
  wire [31:0] _T_1648; // @[Mux.scala 31:69:@14014.4]
  wire  _T_1637; // @[package.scala 96:25:@13987.4 package.scala 96:25:@13988.4]
  wire [31:0] _T_1649; // @[Mux.scala 31:69:@14015.4]
  wire  _T_1634; // @[package.scala 96:25:@13979.4 package.scala 96:25:@13980.4]
  wire [31:0] _T_1650; // @[Mux.scala 31:69:@14016.4]
  wire  _T_1631; // @[package.scala 96:25:@13971.4 package.scala 96:25:@13972.4]
  wire [31:0] _T_1651; // @[Mux.scala 31:69:@14017.4]
  wire  _T_1628; // @[package.scala 96:25:@13963.4 package.scala 96:25:@13964.4]
  wire [31:0] _T_1652; // @[Mux.scala 31:69:@14018.4]
  wire  _T_1625; // @[package.scala 96:25:@13955.4 package.scala 96:25:@13956.4]
  wire [31:0] _T_1653; // @[Mux.scala 31:69:@14019.4]
  wire  _T_1622; // @[package.scala 96:25:@13947.4 package.scala 96:25:@13948.4]
  wire [31:0] _T_1654; // @[Mux.scala 31:69:@14020.4]
  wire  _T_1619; // @[package.scala 96:25:@13939.4 package.scala 96:25:@13940.4]
  wire [31:0] _T_1655; // @[Mux.scala 31:69:@14021.4]
  wire  _T_1616; // @[package.scala 96:25:@13931.4 package.scala 96:25:@13932.4]
  wire [31:0] _T_1656; // @[Mux.scala 31:69:@14022.4]
  wire  _T_1613; // @[package.scala 96:25:@13923.4 package.scala 96:25:@13924.4]
  wire  _T_1750; // @[package.scala 96:25:@14147.4 package.scala 96:25:@14148.4]
  wire [31:0] _T_1754; // @[Mux.scala 31:69:@14157.4]
  wire  _T_1747; // @[package.scala 96:25:@14139.4 package.scala 96:25:@14140.4]
  wire [31:0] _T_1755; // @[Mux.scala 31:69:@14158.4]
  wire  _T_1744; // @[package.scala 96:25:@14131.4 package.scala 96:25:@14132.4]
  wire [31:0] _T_1756; // @[Mux.scala 31:69:@14159.4]
  wire  _T_1741; // @[package.scala 96:25:@14123.4 package.scala 96:25:@14124.4]
  wire [31:0] _T_1757; // @[Mux.scala 31:69:@14160.4]
  wire  _T_1738; // @[package.scala 96:25:@14115.4 package.scala 96:25:@14116.4]
  wire [31:0] _T_1758; // @[Mux.scala 31:69:@14161.4]
  wire  _T_1735; // @[package.scala 96:25:@14107.4 package.scala 96:25:@14108.4]
  wire [31:0] _T_1759; // @[Mux.scala 31:69:@14162.4]
  wire  _T_1732; // @[package.scala 96:25:@14099.4 package.scala 96:25:@14100.4]
  wire [31:0] _T_1760; // @[Mux.scala 31:69:@14163.4]
  wire  _T_1729; // @[package.scala 96:25:@14091.4 package.scala 96:25:@14092.4]
  wire [31:0] _T_1761; // @[Mux.scala 31:69:@14164.4]
  wire  _T_1726; // @[package.scala 96:25:@14083.4 package.scala 96:25:@14084.4]
  wire [31:0] _T_1762; // @[Mux.scala 31:69:@14165.4]
  wire  _T_1723; // @[package.scala 96:25:@14075.4 package.scala 96:25:@14076.4]
  wire [31:0] _T_1763; // @[Mux.scala 31:69:@14166.4]
  wire  _T_1720; // @[package.scala 96:25:@14067.4 package.scala 96:25:@14068.4]
  wire  _T_1857; // @[package.scala 96:25:@14291.4 package.scala 96:25:@14292.4]
  wire [31:0] _T_1861; // @[Mux.scala 31:69:@14301.4]
  wire  _T_1854; // @[package.scala 96:25:@14283.4 package.scala 96:25:@14284.4]
  wire [31:0] _T_1862; // @[Mux.scala 31:69:@14302.4]
  wire  _T_1851; // @[package.scala 96:25:@14275.4 package.scala 96:25:@14276.4]
  wire [31:0] _T_1863; // @[Mux.scala 31:69:@14303.4]
  wire  _T_1848; // @[package.scala 96:25:@14267.4 package.scala 96:25:@14268.4]
  wire [31:0] _T_1864; // @[Mux.scala 31:69:@14304.4]
  wire  _T_1845; // @[package.scala 96:25:@14259.4 package.scala 96:25:@14260.4]
  wire [31:0] _T_1865; // @[Mux.scala 31:69:@14305.4]
  wire  _T_1842; // @[package.scala 96:25:@14251.4 package.scala 96:25:@14252.4]
  wire [31:0] _T_1866; // @[Mux.scala 31:69:@14306.4]
  wire  _T_1839; // @[package.scala 96:25:@14243.4 package.scala 96:25:@14244.4]
  wire [31:0] _T_1867; // @[Mux.scala 31:69:@14307.4]
  wire  _T_1836; // @[package.scala 96:25:@14235.4 package.scala 96:25:@14236.4]
  wire [31:0] _T_1868; // @[Mux.scala 31:69:@14308.4]
  wire  _T_1833; // @[package.scala 96:25:@14227.4 package.scala 96:25:@14228.4]
  wire [31:0] _T_1869; // @[Mux.scala 31:69:@14309.4]
  wire  _T_1830; // @[package.scala 96:25:@14219.4 package.scala 96:25:@14220.4]
  wire [31:0] _T_1870; // @[Mux.scala 31:69:@14310.4]
  wire  _T_1827; // @[package.scala 96:25:@14211.4 package.scala 96:25:@14212.4]
  wire  _T_1964; // @[package.scala 96:25:@14435.4 package.scala 96:25:@14436.4]
  wire [31:0] _T_1968; // @[Mux.scala 31:69:@14445.4]
  wire  _T_1961; // @[package.scala 96:25:@14427.4 package.scala 96:25:@14428.4]
  wire [31:0] _T_1969; // @[Mux.scala 31:69:@14446.4]
  wire  _T_1958; // @[package.scala 96:25:@14419.4 package.scala 96:25:@14420.4]
  wire [31:0] _T_1970; // @[Mux.scala 31:69:@14447.4]
  wire  _T_1955; // @[package.scala 96:25:@14411.4 package.scala 96:25:@14412.4]
  wire [31:0] _T_1971; // @[Mux.scala 31:69:@14448.4]
  wire  _T_1952; // @[package.scala 96:25:@14403.4 package.scala 96:25:@14404.4]
  wire [31:0] _T_1972; // @[Mux.scala 31:69:@14449.4]
  wire  _T_1949; // @[package.scala 96:25:@14395.4 package.scala 96:25:@14396.4]
  wire [31:0] _T_1973; // @[Mux.scala 31:69:@14450.4]
  wire  _T_1946; // @[package.scala 96:25:@14387.4 package.scala 96:25:@14388.4]
  wire [31:0] _T_1974; // @[Mux.scala 31:69:@14451.4]
  wire  _T_1943; // @[package.scala 96:25:@14379.4 package.scala 96:25:@14380.4]
  wire [31:0] _T_1975; // @[Mux.scala 31:69:@14452.4]
  wire  _T_1940; // @[package.scala 96:25:@14371.4 package.scala 96:25:@14372.4]
  wire [31:0] _T_1976; // @[Mux.scala 31:69:@14453.4]
  wire  _T_1937; // @[package.scala 96:25:@14363.4 package.scala 96:25:@14364.4]
  wire [31:0] _T_1977; // @[Mux.scala 31:69:@14454.4]
  wire  _T_1934; // @[package.scala 96:25:@14355.4 package.scala 96:25:@14356.4]
  wire  _T_2071; // @[package.scala 96:25:@14579.4 package.scala 96:25:@14580.4]
  wire [31:0] _T_2075; // @[Mux.scala 31:69:@14589.4]
  wire  _T_2068; // @[package.scala 96:25:@14571.4 package.scala 96:25:@14572.4]
  wire [31:0] _T_2076; // @[Mux.scala 31:69:@14590.4]
  wire  _T_2065; // @[package.scala 96:25:@14563.4 package.scala 96:25:@14564.4]
  wire [31:0] _T_2077; // @[Mux.scala 31:69:@14591.4]
  wire  _T_2062; // @[package.scala 96:25:@14555.4 package.scala 96:25:@14556.4]
  wire [31:0] _T_2078; // @[Mux.scala 31:69:@14592.4]
  wire  _T_2059; // @[package.scala 96:25:@14547.4 package.scala 96:25:@14548.4]
  wire [31:0] _T_2079; // @[Mux.scala 31:69:@14593.4]
  wire  _T_2056; // @[package.scala 96:25:@14539.4 package.scala 96:25:@14540.4]
  wire [31:0] _T_2080; // @[Mux.scala 31:69:@14594.4]
  wire  _T_2053; // @[package.scala 96:25:@14531.4 package.scala 96:25:@14532.4]
  wire [31:0] _T_2081; // @[Mux.scala 31:69:@14595.4]
  wire  _T_2050; // @[package.scala 96:25:@14523.4 package.scala 96:25:@14524.4]
  wire [31:0] _T_2082; // @[Mux.scala 31:69:@14596.4]
  wire  _T_2047; // @[package.scala 96:25:@14515.4 package.scala 96:25:@14516.4]
  wire [31:0] _T_2083; // @[Mux.scala 31:69:@14597.4]
  wire  _T_2044; // @[package.scala 96:25:@14507.4 package.scala 96:25:@14508.4]
  wire [31:0] _T_2084; // @[Mux.scala 31:69:@14598.4]
  wire  _T_2041; // @[package.scala 96:25:@14499.4 package.scala 96:25:@14500.4]
  wire  _T_2178; // @[package.scala 96:25:@14723.4 package.scala 96:25:@14724.4]
  wire [31:0] _T_2182; // @[Mux.scala 31:69:@14733.4]
  wire  _T_2175; // @[package.scala 96:25:@14715.4 package.scala 96:25:@14716.4]
  wire [31:0] _T_2183; // @[Mux.scala 31:69:@14734.4]
  wire  _T_2172; // @[package.scala 96:25:@14707.4 package.scala 96:25:@14708.4]
  wire [31:0] _T_2184; // @[Mux.scala 31:69:@14735.4]
  wire  _T_2169; // @[package.scala 96:25:@14699.4 package.scala 96:25:@14700.4]
  wire [31:0] _T_2185; // @[Mux.scala 31:69:@14736.4]
  wire  _T_2166; // @[package.scala 96:25:@14691.4 package.scala 96:25:@14692.4]
  wire [31:0] _T_2186; // @[Mux.scala 31:69:@14737.4]
  wire  _T_2163; // @[package.scala 96:25:@14683.4 package.scala 96:25:@14684.4]
  wire [31:0] _T_2187; // @[Mux.scala 31:69:@14738.4]
  wire  _T_2160; // @[package.scala 96:25:@14675.4 package.scala 96:25:@14676.4]
  wire [31:0] _T_2188; // @[Mux.scala 31:69:@14739.4]
  wire  _T_2157; // @[package.scala 96:25:@14667.4 package.scala 96:25:@14668.4]
  wire [31:0] _T_2189; // @[Mux.scala 31:69:@14740.4]
  wire  _T_2154; // @[package.scala 96:25:@14659.4 package.scala 96:25:@14660.4]
  wire [31:0] _T_2190; // @[Mux.scala 31:69:@14741.4]
  wire  _T_2151; // @[package.scala 96:25:@14651.4 package.scala 96:25:@14652.4]
  wire [31:0] _T_2191; // @[Mux.scala 31:69:@14742.4]
  wire  _T_2148; // @[package.scala 96:25:@14643.4 package.scala 96:25:@14644.4]
  wire  _T_2285; // @[package.scala 96:25:@14867.4 package.scala 96:25:@14868.4]
  wire [31:0] _T_2289; // @[Mux.scala 31:69:@14877.4]
  wire  _T_2282; // @[package.scala 96:25:@14859.4 package.scala 96:25:@14860.4]
  wire [31:0] _T_2290; // @[Mux.scala 31:69:@14878.4]
  wire  _T_2279; // @[package.scala 96:25:@14851.4 package.scala 96:25:@14852.4]
  wire [31:0] _T_2291; // @[Mux.scala 31:69:@14879.4]
  wire  _T_2276; // @[package.scala 96:25:@14843.4 package.scala 96:25:@14844.4]
  wire [31:0] _T_2292; // @[Mux.scala 31:69:@14880.4]
  wire  _T_2273; // @[package.scala 96:25:@14835.4 package.scala 96:25:@14836.4]
  wire [31:0] _T_2293; // @[Mux.scala 31:69:@14881.4]
  wire  _T_2270; // @[package.scala 96:25:@14827.4 package.scala 96:25:@14828.4]
  wire [31:0] _T_2294; // @[Mux.scala 31:69:@14882.4]
  wire  _T_2267; // @[package.scala 96:25:@14819.4 package.scala 96:25:@14820.4]
  wire [31:0] _T_2295; // @[Mux.scala 31:69:@14883.4]
  wire  _T_2264; // @[package.scala 96:25:@14811.4 package.scala 96:25:@14812.4]
  wire [31:0] _T_2296; // @[Mux.scala 31:69:@14884.4]
  wire  _T_2261; // @[package.scala 96:25:@14803.4 package.scala 96:25:@14804.4]
  wire [31:0] _T_2297; // @[Mux.scala 31:69:@14885.4]
  wire  _T_2258; // @[package.scala 96:25:@14795.4 package.scala 96:25:@14796.4]
  wire [31:0] _T_2298; // @[Mux.scala 31:69:@14886.4]
  wire  _T_2255; // @[package.scala 96:25:@14787.4 package.scala 96:25:@14788.4]
  wire  _T_2392; // @[package.scala 96:25:@15011.4 package.scala 96:25:@15012.4]
  wire [31:0] _T_2396; // @[Mux.scala 31:69:@15021.4]
  wire  _T_2389; // @[package.scala 96:25:@15003.4 package.scala 96:25:@15004.4]
  wire [31:0] _T_2397; // @[Mux.scala 31:69:@15022.4]
  wire  _T_2386; // @[package.scala 96:25:@14995.4 package.scala 96:25:@14996.4]
  wire [31:0] _T_2398; // @[Mux.scala 31:69:@15023.4]
  wire  _T_2383; // @[package.scala 96:25:@14987.4 package.scala 96:25:@14988.4]
  wire [31:0] _T_2399; // @[Mux.scala 31:69:@15024.4]
  wire  _T_2380; // @[package.scala 96:25:@14979.4 package.scala 96:25:@14980.4]
  wire [31:0] _T_2400; // @[Mux.scala 31:69:@15025.4]
  wire  _T_2377; // @[package.scala 96:25:@14971.4 package.scala 96:25:@14972.4]
  wire [31:0] _T_2401; // @[Mux.scala 31:69:@15026.4]
  wire  _T_2374; // @[package.scala 96:25:@14963.4 package.scala 96:25:@14964.4]
  wire [31:0] _T_2402; // @[Mux.scala 31:69:@15027.4]
  wire  _T_2371; // @[package.scala 96:25:@14955.4 package.scala 96:25:@14956.4]
  wire [31:0] _T_2403; // @[Mux.scala 31:69:@15028.4]
  wire  _T_2368; // @[package.scala 96:25:@14947.4 package.scala 96:25:@14948.4]
  wire [31:0] _T_2404; // @[Mux.scala 31:69:@15029.4]
  wire  _T_2365; // @[package.scala 96:25:@14939.4 package.scala 96:25:@14940.4]
  wire [31:0] _T_2405; // @[Mux.scala 31:69:@15030.4]
  wire  _T_2362; // @[package.scala 96:25:@14931.4 package.scala 96:25:@14932.4]
  wire  _T_2499; // @[package.scala 96:25:@15155.4 package.scala 96:25:@15156.4]
  wire [31:0] _T_2503; // @[Mux.scala 31:69:@15165.4]
  wire  _T_2496; // @[package.scala 96:25:@15147.4 package.scala 96:25:@15148.4]
  wire [31:0] _T_2504; // @[Mux.scala 31:69:@15166.4]
  wire  _T_2493; // @[package.scala 96:25:@15139.4 package.scala 96:25:@15140.4]
  wire [31:0] _T_2505; // @[Mux.scala 31:69:@15167.4]
  wire  _T_2490; // @[package.scala 96:25:@15131.4 package.scala 96:25:@15132.4]
  wire [31:0] _T_2506; // @[Mux.scala 31:69:@15168.4]
  wire  _T_2487; // @[package.scala 96:25:@15123.4 package.scala 96:25:@15124.4]
  wire [31:0] _T_2507; // @[Mux.scala 31:69:@15169.4]
  wire  _T_2484; // @[package.scala 96:25:@15115.4 package.scala 96:25:@15116.4]
  wire [31:0] _T_2508; // @[Mux.scala 31:69:@15170.4]
  wire  _T_2481; // @[package.scala 96:25:@15107.4 package.scala 96:25:@15108.4]
  wire [31:0] _T_2509; // @[Mux.scala 31:69:@15171.4]
  wire  _T_2478; // @[package.scala 96:25:@15099.4 package.scala 96:25:@15100.4]
  wire [31:0] _T_2510; // @[Mux.scala 31:69:@15172.4]
  wire  _T_2475; // @[package.scala 96:25:@15091.4 package.scala 96:25:@15092.4]
  wire [31:0] _T_2511; // @[Mux.scala 31:69:@15173.4]
  wire  _T_2472; // @[package.scala 96:25:@15083.4 package.scala 96:25:@15084.4]
  wire [31:0] _T_2512; // @[Mux.scala 31:69:@15174.4]
  wire  _T_2469; // @[package.scala 96:25:@15075.4 package.scala 96:25:@15076.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@12477.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@12493.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@12509.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@12525.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@12541.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@12557.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@12573.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@12589.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@12605.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@12621.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@12637.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@12653.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 124:33:@12849.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_ins_6(StickySelects_io_ins_6),
    .io_ins_7(StickySelects_io_ins_7),
    .io_ins_8(StickySelects_io_ins_8),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5),
    .io_outs_6(StickySelects_io_outs_6),
    .io_outs_7(StickySelects_io_outs_7),
    .io_outs_8(StickySelects_io_outs_8)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@12938.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_ins_6(StickySelects_1_io_ins_6),
    .io_ins_7(StickySelects_1_io_ins_7),
    .io_ins_8(StickySelects_1_io_ins_8),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5),
    .io_outs_6(StickySelects_1_io_outs_6),
    .io_outs_7(StickySelects_1_io_outs_7),
    .io_outs_8(StickySelects_1_io_outs_8)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@13027.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_ins_8(StickySelects_2_io_ins_8),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7),
    .io_outs_8(StickySelects_2_io_outs_8)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@13116.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_ins_8(StickySelects_3_io_ins_8),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7),
    .io_outs_8(StickySelects_3_io_outs_8)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@13205.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_ins_6(StickySelects_4_io_ins_6),
    .io_ins_7(StickySelects_4_io_ins_7),
    .io_ins_8(StickySelects_4_io_ins_8),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5),
    .io_outs_6(StickySelects_4_io_outs_6),
    .io_outs_7(StickySelects_4_io_outs_7),
    .io_outs_8(StickySelects_4_io_outs_8)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@13294.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_ins_6(StickySelects_5_io_ins_6),
    .io_ins_7(StickySelects_5_io_ins_7),
    .io_ins_8(StickySelects_5_io_ins_8),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5),
    .io_outs_6(StickySelects_5_io_outs_6),
    .io_outs_7(StickySelects_5_io_outs_7),
    .io_outs_8(StickySelects_5_io_outs_8)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@13383.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_ins_8(StickySelects_6_io_ins_8),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7),
    .io_outs_8(StickySelects_6_io_outs_8)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@13472.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_ins_8(StickySelects_7_io_ins_8),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7),
    .io_outs_8(StickySelects_7_io_outs_8)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@13561.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_ins_6(StickySelects_8_io_ins_6),
    .io_ins_7(StickySelects_8_io_ins_7),
    .io_ins_8(StickySelects_8_io_ins_8),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5),
    .io_outs_6(StickySelects_8_io_outs_6),
    .io_outs_7(StickySelects_8_io_outs_7),
    .io_outs_8(StickySelects_8_io_outs_8)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@13650.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_ins_6(StickySelects_9_io_ins_6),
    .io_ins_7(StickySelects_9_io_ins_7),
    .io_ins_8(StickySelects_9_io_ins_8),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5),
    .io_outs_6(StickySelects_9_io_outs_6),
    .io_outs_7(StickySelects_9_io_outs_7),
    .io_outs_8(StickySelects_9_io_outs_8)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@13739.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_ins_8(StickySelects_10_io_ins_8),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7),
    .io_outs_8(StickySelects_10_io_outs_8)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@13828.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_ins_8(StickySelects_11_io_ins_8),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7),
    .io_outs_8(StickySelects_11_io_outs_8)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@13918.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@13926.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@13934.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@13942.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@13950.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@13958.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@13966.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@13974.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@13982.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@13990.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@13998.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@14006.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@14062.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@14070.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@14078.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@14086.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@14094.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@14102.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@14110.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@14118.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@14126.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@14134.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@14142.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@14150.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@14206.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@14214.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@14222.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@14230.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@14238.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@14246.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@14254.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@14262.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@14270.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@14278.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@14286.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@14294.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@14350.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@14358.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@14366.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@14374.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@14382.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@14390.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@14398.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@14406.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@14414.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@14422.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@14430.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@14438.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@14494.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@14502.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@14510.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@14518.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@14526.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@14534.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@14542.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@14550.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@14558.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@14566.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@14574.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@14582.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@14638.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@14646.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@14654.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@14662.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@14670.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@14678.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@14686.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@14694.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@14702.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@14710.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@14718.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@14726.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@14782.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@14790.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@14798.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@14806.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@14814.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@14822.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@14830.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@14838.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@14846.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@14854.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@14862.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@14870.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@14926.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@14934.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@14942.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@14950.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@14958.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@14966.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@14974.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@14982.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@14990.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@14998.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@15006.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@15014.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_96 ( // @[package.scala 93:22:@15070.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_97 ( // @[package.scala 93:22:@15078.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_98 ( // @[package.scala 93:22:@15086.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_99 ( // @[package.scala 93:22:@15094.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_100 ( // @[package.scala 93:22:@15102.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_101 ( // @[package.scala 93:22:@15110.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_102 ( // @[package.scala 93:22:@15118.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_103 ( // @[package.scala 93:22:@15126.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_104 ( // @[package.scala 93:22:@15134.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_105 ( // @[package.scala 93:22:@15142.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_106 ( // @[package.scala 93:22:@15150.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_107 ( // @[package.scala 93:22:@15158.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  assign _T_316 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@12669.4]
  assign _T_318 = io_wPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 82:210:@12670.4]
  assign _T_319 = _T_316 & _T_318; // @[MemPrimitives.scala 82:228:@12671.4]
  assign _T_320 = io_wPort_0_en_0 & _T_319; // @[MemPrimitives.scala 83:102:@12672.4]
  assign _T_322 = {_T_320,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12674.4]
  assign _T_329 = io_wPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 82:210:@12682.4]
  assign _T_330 = _T_316 & _T_329; // @[MemPrimitives.scala 82:228:@12683.4]
  assign _T_331 = io_wPort_0_en_0 & _T_330; // @[MemPrimitives.scala 83:102:@12684.4]
  assign _T_333 = {_T_331,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12686.4]
  assign _T_340 = io_wPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 82:210:@12694.4]
  assign _T_341 = _T_316 & _T_340; // @[MemPrimitives.scala 82:228:@12695.4]
  assign _T_342 = io_wPort_0_en_0 & _T_341; // @[MemPrimitives.scala 83:102:@12696.4]
  assign _T_344 = {_T_342,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12698.4]
  assign _T_349 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@12705.4]
  assign _T_352 = _T_349 & _T_318; // @[MemPrimitives.scala 82:228:@12707.4]
  assign _T_353 = io_wPort_0_en_0 & _T_352; // @[MemPrimitives.scala 83:102:@12708.4]
  assign _T_355 = {_T_353,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12710.4]
  assign _T_363 = _T_349 & _T_329; // @[MemPrimitives.scala 82:228:@12719.4]
  assign _T_364 = io_wPort_0_en_0 & _T_363; // @[MemPrimitives.scala 83:102:@12720.4]
  assign _T_366 = {_T_364,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12722.4]
  assign _T_374 = _T_349 & _T_340; // @[MemPrimitives.scala 82:228:@12731.4]
  assign _T_375 = io_wPort_0_en_0 & _T_374; // @[MemPrimitives.scala 83:102:@12732.4]
  assign _T_377 = {_T_375,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12734.4]
  assign _T_382 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@12741.4]
  assign _T_385 = _T_382 & _T_318; // @[MemPrimitives.scala 82:228:@12743.4]
  assign _T_386 = io_wPort_0_en_0 & _T_385; // @[MemPrimitives.scala 83:102:@12744.4]
  assign _T_388 = {_T_386,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12746.4]
  assign _T_396 = _T_382 & _T_329; // @[MemPrimitives.scala 82:228:@12755.4]
  assign _T_397 = io_wPort_0_en_0 & _T_396; // @[MemPrimitives.scala 83:102:@12756.4]
  assign _T_399 = {_T_397,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12758.4]
  assign _T_407 = _T_382 & _T_340; // @[MemPrimitives.scala 82:228:@12767.4]
  assign _T_408 = io_wPort_0_en_0 & _T_407; // @[MemPrimitives.scala 83:102:@12768.4]
  assign _T_410 = {_T_408,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12770.4]
  assign _T_415 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@12777.4]
  assign _T_418 = _T_415 & _T_318; // @[MemPrimitives.scala 82:228:@12779.4]
  assign _T_419 = io_wPort_0_en_0 & _T_418; // @[MemPrimitives.scala 83:102:@12780.4]
  assign _T_421 = {_T_419,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12782.4]
  assign _T_429 = _T_415 & _T_329; // @[MemPrimitives.scala 82:228:@12791.4]
  assign _T_430 = io_wPort_0_en_0 & _T_429; // @[MemPrimitives.scala 83:102:@12792.4]
  assign _T_432 = {_T_430,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12794.4]
  assign _T_440 = _T_415 & _T_340; // @[MemPrimitives.scala 82:228:@12803.4]
  assign _T_441 = io_wPort_0_en_0 & _T_440; // @[MemPrimitives.scala 83:102:@12804.4]
  assign _T_443 = {_T_441,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12806.4]
  assign _T_448 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12813.4]
  assign _T_450 = io_rPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12814.4]
  assign _T_451 = _T_448 & _T_450; // @[MemPrimitives.scala 110:228:@12815.4]
  assign _T_454 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12817.4]
  assign _T_456 = io_rPort_1_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12818.4]
  assign _T_457 = _T_454 & _T_456; // @[MemPrimitives.scala 110:228:@12819.4]
  assign _T_460 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12821.4]
  assign _T_462 = io_rPort_2_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12822.4]
  assign _T_463 = _T_460 & _T_462; // @[MemPrimitives.scala 110:228:@12823.4]
  assign _T_466 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12825.4]
  assign _T_468 = io_rPort_3_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12826.4]
  assign _T_469 = _T_466 & _T_468; // @[MemPrimitives.scala 110:228:@12827.4]
  assign _T_472 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12829.4]
  assign _T_474 = io_rPort_4_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12830.4]
  assign _T_475 = _T_472 & _T_474; // @[MemPrimitives.scala 110:228:@12831.4]
  assign _T_478 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12833.4]
  assign _T_480 = io_rPort_5_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12834.4]
  assign _T_481 = _T_478 & _T_480; // @[MemPrimitives.scala 110:228:@12835.4]
  assign _T_484 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12837.4]
  assign _T_486 = io_rPort_6_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12838.4]
  assign _T_487 = _T_484 & _T_486; // @[MemPrimitives.scala 110:228:@12839.4]
  assign _T_490 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12841.4]
  assign _T_492 = io_rPort_7_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12842.4]
  assign _T_493 = _T_490 & _T_492; // @[MemPrimitives.scala 110:228:@12843.4]
  assign _T_496 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12845.4]
  assign _T_498 = io_rPort_8_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12846.4]
  assign _T_499 = _T_496 & _T_498; // @[MemPrimitives.scala 110:228:@12847.4]
  assign _T_501 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@12861.4]
  assign _T_502 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@12862.4]
  assign _T_503 = StickySelects_io_outs_2; // @[MemPrimitives.scala 126:35:@12863.4]
  assign _T_504 = StickySelects_io_outs_3; // @[MemPrimitives.scala 126:35:@12864.4]
  assign _T_505 = StickySelects_io_outs_4; // @[MemPrimitives.scala 126:35:@12865.4]
  assign _T_506 = StickySelects_io_outs_5; // @[MemPrimitives.scala 126:35:@12866.4]
  assign _T_507 = StickySelects_io_outs_6; // @[MemPrimitives.scala 126:35:@12867.4]
  assign _T_508 = StickySelects_io_outs_7; // @[MemPrimitives.scala 126:35:@12868.4]
  assign _T_509 = StickySelects_io_outs_8; // @[MemPrimitives.scala 126:35:@12869.4]
  assign _T_511 = {_T_501,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12871.4]
  assign _T_513 = {_T_502,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12873.4]
  assign _T_515 = {_T_503,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12875.4]
  assign _T_517 = {_T_504,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12877.4]
  assign _T_519 = {_T_505,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12879.4]
  assign _T_521 = {_T_506,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12881.4]
  assign _T_523 = {_T_507,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12883.4]
  assign _T_525 = {_T_508,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12885.4]
  assign _T_527 = {_T_509,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12887.4]
  assign _T_528 = _T_508 ? _T_525 : _T_527; // @[Mux.scala 31:69:@12888.4]
  assign _T_529 = _T_507 ? _T_523 : _T_528; // @[Mux.scala 31:69:@12889.4]
  assign _T_530 = _T_506 ? _T_521 : _T_529; // @[Mux.scala 31:69:@12890.4]
  assign _T_531 = _T_505 ? _T_519 : _T_530; // @[Mux.scala 31:69:@12891.4]
  assign _T_532 = _T_504 ? _T_517 : _T_531; // @[Mux.scala 31:69:@12892.4]
  assign _T_533 = _T_503 ? _T_515 : _T_532; // @[Mux.scala 31:69:@12893.4]
  assign _T_534 = _T_502 ? _T_513 : _T_533; // @[Mux.scala 31:69:@12894.4]
  assign _T_535 = _T_501 ? _T_511 : _T_534; // @[Mux.scala 31:69:@12895.4]
  assign _T_542 = io_rPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12903.4]
  assign _T_543 = _T_448 & _T_542; // @[MemPrimitives.scala 110:228:@12904.4]
  assign _T_548 = io_rPort_1_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12907.4]
  assign _T_549 = _T_454 & _T_548; // @[MemPrimitives.scala 110:228:@12908.4]
  assign _T_554 = io_rPort_2_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12911.4]
  assign _T_555 = _T_460 & _T_554; // @[MemPrimitives.scala 110:228:@12912.4]
  assign _T_560 = io_rPort_3_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12915.4]
  assign _T_561 = _T_466 & _T_560; // @[MemPrimitives.scala 110:228:@12916.4]
  assign _T_566 = io_rPort_4_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12919.4]
  assign _T_567 = _T_472 & _T_566; // @[MemPrimitives.scala 110:228:@12920.4]
  assign _T_572 = io_rPort_5_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12923.4]
  assign _T_573 = _T_478 & _T_572; // @[MemPrimitives.scala 110:228:@12924.4]
  assign _T_578 = io_rPort_6_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12927.4]
  assign _T_579 = _T_484 & _T_578; // @[MemPrimitives.scala 110:228:@12928.4]
  assign _T_584 = io_rPort_7_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12931.4]
  assign _T_585 = _T_490 & _T_584; // @[MemPrimitives.scala 110:228:@12932.4]
  assign _T_590 = io_rPort_8_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12935.4]
  assign _T_591 = _T_496 & _T_590; // @[MemPrimitives.scala 110:228:@12936.4]
  assign _T_593 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@12950.4]
  assign _T_594 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@12951.4]
  assign _T_595 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@12952.4]
  assign _T_596 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@12953.4]
  assign _T_597 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 126:35:@12954.4]
  assign _T_598 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 126:35:@12955.4]
  assign _T_599 = StickySelects_1_io_outs_6; // @[MemPrimitives.scala 126:35:@12956.4]
  assign _T_600 = StickySelects_1_io_outs_7; // @[MemPrimitives.scala 126:35:@12957.4]
  assign _T_601 = StickySelects_1_io_outs_8; // @[MemPrimitives.scala 126:35:@12958.4]
  assign _T_603 = {_T_593,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12960.4]
  assign _T_605 = {_T_594,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12962.4]
  assign _T_607 = {_T_595,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12964.4]
  assign _T_609 = {_T_596,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12966.4]
  assign _T_611 = {_T_597,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12968.4]
  assign _T_613 = {_T_598,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12970.4]
  assign _T_615 = {_T_599,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12972.4]
  assign _T_617 = {_T_600,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12974.4]
  assign _T_619 = {_T_601,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12976.4]
  assign _T_620 = _T_600 ? _T_617 : _T_619; // @[Mux.scala 31:69:@12977.4]
  assign _T_621 = _T_599 ? _T_615 : _T_620; // @[Mux.scala 31:69:@12978.4]
  assign _T_622 = _T_598 ? _T_613 : _T_621; // @[Mux.scala 31:69:@12979.4]
  assign _T_623 = _T_597 ? _T_611 : _T_622; // @[Mux.scala 31:69:@12980.4]
  assign _T_624 = _T_596 ? _T_609 : _T_623; // @[Mux.scala 31:69:@12981.4]
  assign _T_625 = _T_595 ? _T_607 : _T_624; // @[Mux.scala 31:69:@12982.4]
  assign _T_626 = _T_594 ? _T_605 : _T_625; // @[Mux.scala 31:69:@12983.4]
  assign _T_627 = _T_593 ? _T_603 : _T_626; // @[Mux.scala 31:69:@12984.4]
  assign _T_634 = io_rPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@12992.4]
  assign _T_635 = _T_448 & _T_634; // @[MemPrimitives.scala 110:228:@12993.4]
  assign _T_640 = io_rPort_1_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@12996.4]
  assign _T_641 = _T_454 & _T_640; // @[MemPrimitives.scala 110:228:@12997.4]
  assign _T_646 = io_rPort_2_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13000.4]
  assign _T_647 = _T_460 & _T_646; // @[MemPrimitives.scala 110:228:@13001.4]
  assign _T_652 = io_rPort_3_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13004.4]
  assign _T_653 = _T_466 & _T_652; // @[MemPrimitives.scala 110:228:@13005.4]
  assign _T_658 = io_rPort_4_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13008.4]
  assign _T_659 = _T_472 & _T_658; // @[MemPrimitives.scala 110:228:@13009.4]
  assign _T_664 = io_rPort_5_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13012.4]
  assign _T_665 = _T_478 & _T_664; // @[MemPrimitives.scala 110:228:@13013.4]
  assign _T_670 = io_rPort_6_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13016.4]
  assign _T_671 = _T_484 & _T_670; // @[MemPrimitives.scala 110:228:@13017.4]
  assign _T_676 = io_rPort_7_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13020.4]
  assign _T_677 = _T_490 & _T_676; // @[MemPrimitives.scala 110:228:@13021.4]
  assign _T_682 = io_rPort_8_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13024.4]
  assign _T_683 = _T_496 & _T_682; // @[MemPrimitives.scala 110:228:@13025.4]
  assign _T_685 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@13039.4]
  assign _T_686 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@13040.4]
  assign _T_687 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 126:35:@13041.4]
  assign _T_688 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 126:35:@13042.4]
  assign _T_689 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 126:35:@13043.4]
  assign _T_690 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 126:35:@13044.4]
  assign _T_691 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 126:35:@13045.4]
  assign _T_692 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 126:35:@13046.4]
  assign _T_693 = StickySelects_2_io_outs_8; // @[MemPrimitives.scala 126:35:@13047.4]
  assign _T_695 = {_T_685,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13049.4]
  assign _T_697 = {_T_686,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13051.4]
  assign _T_699 = {_T_687,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13053.4]
  assign _T_701 = {_T_688,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13055.4]
  assign _T_703 = {_T_689,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13057.4]
  assign _T_705 = {_T_690,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13059.4]
  assign _T_707 = {_T_691,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13061.4]
  assign _T_709 = {_T_692,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13063.4]
  assign _T_711 = {_T_693,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13065.4]
  assign _T_712 = _T_692 ? _T_709 : _T_711; // @[Mux.scala 31:69:@13066.4]
  assign _T_713 = _T_691 ? _T_707 : _T_712; // @[Mux.scala 31:69:@13067.4]
  assign _T_714 = _T_690 ? _T_705 : _T_713; // @[Mux.scala 31:69:@13068.4]
  assign _T_715 = _T_689 ? _T_703 : _T_714; // @[Mux.scala 31:69:@13069.4]
  assign _T_716 = _T_688 ? _T_701 : _T_715; // @[Mux.scala 31:69:@13070.4]
  assign _T_717 = _T_687 ? _T_699 : _T_716; // @[Mux.scala 31:69:@13071.4]
  assign _T_718 = _T_686 ? _T_697 : _T_717; // @[Mux.scala 31:69:@13072.4]
  assign _T_719 = _T_685 ? _T_695 : _T_718; // @[Mux.scala 31:69:@13073.4]
  assign _T_724 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13080.4]
  assign _T_727 = _T_724 & _T_450; // @[MemPrimitives.scala 110:228:@13082.4]
  assign _T_730 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13084.4]
  assign _T_733 = _T_730 & _T_456; // @[MemPrimitives.scala 110:228:@13086.4]
  assign _T_736 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13088.4]
  assign _T_739 = _T_736 & _T_462; // @[MemPrimitives.scala 110:228:@13090.4]
  assign _T_742 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13092.4]
  assign _T_745 = _T_742 & _T_468; // @[MemPrimitives.scala 110:228:@13094.4]
  assign _T_748 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13096.4]
  assign _T_751 = _T_748 & _T_474; // @[MemPrimitives.scala 110:228:@13098.4]
  assign _T_754 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13100.4]
  assign _T_757 = _T_754 & _T_480; // @[MemPrimitives.scala 110:228:@13102.4]
  assign _T_760 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13104.4]
  assign _T_763 = _T_760 & _T_486; // @[MemPrimitives.scala 110:228:@13106.4]
  assign _T_766 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13108.4]
  assign _T_769 = _T_766 & _T_492; // @[MemPrimitives.scala 110:228:@13110.4]
  assign _T_772 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13112.4]
  assign _T_775 = _T_772 & _T_498; // @[MemPrimitives.scala 110:228:@13114.4]
  assign _T_777 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@13128.4]
  assign _T_778 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@13129.4]
  assign _T_779 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@13130.4]
  assign _T_780 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@13131.4]
  assign _T_781 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 126:35:@13132.4]
  assign _T_782 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 126:35:@13133.4]
  assign _T_783 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 126:35:@13134.4]
  assign _T_784 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 126:35:@13135.4]
  assign _T_785 = StickySelects_3_io_outs_8; // @[MemPrimitives.scala 126:35:@13136.4]
  assign _T_787 = {_T_777,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13138.4]
  assign _T_789 = {_T_778,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13140.4]
  assign _T_791 = {_T_779,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13142.4]
  assign _T_793 = {_T_780,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13144.4]
  assign _T_795 = {_T_781,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13146.4]
  assign _T_797 = {_T_782,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13148.4]
  assign _T_799 = {_T_783,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13150.4]
  assign _T_801 = {_T_784,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13152.4]
  assign _T_803 = {_T_785,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13154.4]
  assign _T_804 = _T_784 ? _T_801 : _T_803; // @[Mux.scala 31:69:@13155.4]
  assign _T_805 = _T_783 ? _T_799 : _T_804; // @[Mux.scala 31:69:@13156.4]
  assign _T_806 = _T_782 ? _T_797 : _T_805; // @[Mux.scala 31:69:@13157.4]
  assign _T_807 = _T_781 ? _T_795 : _T_806; // @[Mux.scala 31:69:@13158.4]
  assign _T_808 = _T_780 ? _T_793 : _T_807; // @[Mux.scala 31:69:@13159.4]
  assign _T_809 = _T_779 ? _T_791 : _T_808; // @[Mux.scala 31:69:@13160.4]
  assign _T_810 = _T_778 ? _T_789 : _T_809; // @[Mux.scala 31:69:@13161.4]
  assign _T_811 = _T_777 ? _T_787 : _T_810; // @[Mux.scala 31:69:@13162.4]
  assign _T_819 = _T_724 & _T_542; // @[MemPrimitives.scala 110:228:@13171.4]
  assign _T_825 = _T_730 & _T_548; // @[MemPrimitives.scala 110:228:@13175.4]
  assign _T_831 = _T_736 & _T_554; // @[MemPrimitives.scala 110:228:@13179.4]
  assign _T_837 = _T_742 & _T_560; // @[MemPrimitives.scala 110:228:@13183.4]
  assign _T_843 = _T_748 & _T_566; // @[MemPrimitives.scala 110:228:@13187.4]
  assign _T_849 = _T_754 & _T_572; // @[MemPrimitives.scala 110:228:@13191.4]
  assign _T_855 = _T_760 & _T_578; // @[MemPrimitives.scala 110:228:@13195.4]
  assign _T_861 = _T_766 & _T_584; // @[MemPrimitives.scala 110:228:@13199.4]
  assign _T_867 = _T_772 & _T_590; // @[MemPrimitives.scala 110:228:@13203.4]
  assign _T_869 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@13217.4]
  assign _T_870 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@13218.4]
  assign _T_871 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 126:35:@13219.4]
  assign _T_872 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 126:35:@13220.4]
  assign _T_873 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 126:35:@13221.4]
  assign _T_874 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 126:35:@13222.4]
  assign _T_875 = StickySelects_4_io_outs_6; // @[MemPrimitives.scala 126:35:@13223.4]
  assign _T_876 = StickySelects_4_io_outs_7; // @[MemPrimitives.scala 126:35:@13224.4]
  assign _T_877 = StickySelects_4_io_outs_8; // @[MemPrimitives.scala 126:35:@13225.4]
  assign _T_879 = {_T_869,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13227.4]
  assign _T_881 = {_T_870,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13229.4]
  assign _T_883 = {_T_871,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13231.4]
  assign _T_885 = {_T_872,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13233.4]
  assign _T_887 = {_T_873,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13235.4]
  assign _T_889 = {_T_874,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13237.4]
  assign _T_891 = {_T_875,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13239.4]
  assign _T_893 = {_T_876,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13241.4]
  assign _T_895 = {_T_877,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13243.4]
  assign _T_896 = _T_876 ? _T_893 : _T_895; // @[Mux.scala 31:69:@13244.4]
  assign _T_897 = _T_875 ? _T_891 : _T_896; // @[Mux.scala 31:69:@13245.4]
  assign _T_898 = _T_874 ? _T_889 : _T_897; // @[Mux.scala 31:69:@13246.4]
  assign _T_899 = _T_873 ? _T_887 : _T_898; // @[Mux.scala 31:69:@13247.4]
  assign _T_900 = _T_872 ? _T_885 : _T_899; // @[Mux.scala 31:69:@13248.4]
  assign _T_901 = _T_871 ? _T_883 : _T_900; // @[Mux.scala 31:69:@13249.4]
  assign _T_902 = _T_870 ? _T_881 : _T_901; // @[Mux.scala 31:69:@13250.4]
  assign _T_903 = _T_869 ? _T_879 : _T_902; // @[Mux.scala 31:69:@13251.4]
  assign _T_911 = _T_724 & _T_634; // @[MemPrimitives.scala 110:228:@13260.4]
  assign _T_917 = _T_730 & _T_640; // @[MemPrimitives.scala 110:228:@13264.4]
  assign _T_923 = _T_736 & _T_646; // @[MemPrimitives.scala 110:228:@13268.4]
  assign _T_929 = _T_742 & _T_652; // @[MemPrimitives.scala 110:228:@13272.4]
  assign _T_935 = _T_748 & _T_658; // @[MemPrimitives.scala 110:228:@13276.4]
  assign _T_941 = _T_754 & _T_664; // @[MemPrimitives.scala 110:228:@13280.4]
  assign _T_947 = _T_760 & _T_670; // @[MemPrimitives.scala 110:228:@13284.4]
  assign _T_953 = _T_766 & _T_676; // @[MemPrimitives.scala 110:228:@13288.4]
  assign _T_959 = _T_772 & _T_682; // @[MemPrimitives.scala 110:228:@13292.4]
  assign _T_961 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@13306.4]
  assign _T_962 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@13307.4]
  assign _T_963 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@13308.4]
  assign _T_964 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@13309.4]
  assign _T_965 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 126:35:@13310.4]
  assign _T_966 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 126:35:@13311.4]
  assign _T_967 = StickySelects_5_io_outs_6; // @[MemPrimitives.scala 126:35:@13312.4]
  assign _T_968 = StickySelects_5_io_outs_7; // @[MemPrimitives.scala 126:35:@13313.4]
  assign _T_969 = StickySelects_5_io_outs_8; // @[MemPrimitives.scala 126:35:@13314.4]
  assign _T_971 = {_T_961,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13316.4]
  assign _T_973 = {_T_962,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13318.4]
  assign _T_975 = {_T_963,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13320.4]
  assign _T_977 = {_T_964,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13322.4]
  assign _T_979 = {_T_965,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13324.4]
  assign _T_981 = {_T_966,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13326.4]
  assign _T_983 = {_T_967,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13328.4]
  assign _T_985 = {_T_968,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13330.4]
  assign _T_987 = {_T_969,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13332.4]
  assign _T_988 = _T_968 ? _T_985 : _T_987; // @[Mux.scala 31:69:@13333.4]
  assign _T_989 = _T_967 ? _T_983 : _T_988; // @[Mux.scala 31:69:@13334.4]
  assign _T_990 = _T_966 ? _T_981 : _T_989; // @[Mux.scala 31:69:@13335.4]
  assign _T_991 = _T_965 ? _T_979 : _T_990; // @[Mux.scala 31:69:@13336.4]
  assign _T_992 = _T_964 ? _T_977 : _T_991; // @[Mux.scala 31:69:@13337.4]
  assign _T_993 = _T_963 ? _T_975 : _T_992; // @[Mux.scala 31:69:@13338.4]
  assign _T_994 = _T_962 ? _T_973 : _T_993; // @[Mux.scala 31:69:@13339.4]
  assign _T_995 = _T_961 ? _T_971 : _T_994; // @[Mux.scala 31:69:@13340.4]
  assign _T_1000 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13347.4]
  assign _T_1003 = _T_1000 & _T_450; // @[MemPrimitives.scala 110:228:@13349.4]
  assign _T_1006 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13351.4]
  assign _T_1009 = _T_1006 & _T_456; // @[MemPrimitives.scala 110:228:@13353.4]
  assign _T_1012 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13355.4]
  assign _T_1015 = _T_1012 & _T_462; // @[MemPrimitives.scala 110:228:@13357.4]
  assign _T_1018 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13359.4]
  assign _T_1021 = _T_1018 & _T_468; // @[MemPrimitives.scala 110:228:@13361.4]
  assign _T_1024 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13363.4]
  assign _T_1027 = _T_1024 & _T_474; // @[MemPrimitives.scala 110:228:@13365.4]
  assign _T_1030 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13367.4]
  assign _T_1033 = _T_1030 & _T_480; // @[MemPrimitives.scala 110:228:@13369.4]
  assign _T_1036 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13371.4]
  assign _T_1039 = _T_1036 & _T_486; // @[MemPrimitives.scala 110:228:@13373.4]
  assign _T_1042 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13375.4]
  assign _T_1045 = _T_1042 & _T_492; // @[MemPrimitives.scala 110:228:@13377.4]
  assign _T_1048 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13379.4]
  assign _T_1051 = _T_1048 & _T_498; // @[MemPrimitives.scala 110:228:@13381.4]
  assign _T_1053 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@13395.4]
  assign _T_1054 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@13396.4]
  assign _T_1055 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 126:35:@13397.4]
  assign _T_1056 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 126:35:@13398.4]
  assign _T_1057 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 126:35:@13399.4]
  assign _T_1058 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 126:35:@13400.4]
  assign _T_1059 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 126:35:@13401.4]
  assign _T_1060 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 126:35:@13402.4]
  assign _T_1061 = StickySelects_6_io_outs_8; // @[MemPrimitives.scala 126:35:@13403.4]
  assign _T_1063 = {_T_1053,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13405.4]
  assign _T_1065 = {_T_1054,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13407.4]
  assign _T_1067 = {_T_1055,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13409.4]
  assign _T_1069 = {_T_1056,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13411.4]
  assign _T_1071 = {_T_1057,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13413.4]
  assign _T_1073 = {_T_1058,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13415.4]
  assign _T_1075 = {_T_1059,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13417.4]
  assign _T_1077 = {_T_1060,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13419.4]
  assign _T_1079 = {_T_1061,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13421.4]
  assign _T_1080 = _T_1060 ? _T_1077 : _T_1079; // @[Mux.scala 31:69:@13422.4]
  assign _T_1081 = _T_1059 ? _T_1075 : _T_1080; // @[Mux.scala 31:69:@13423.4]
  assign _T_1082 = _T_1058 ? _T_1073 : _T_1081; // @[Mux.scala 31:69:@13424.4]
  assign _T_1083 = _T_1057 ? _T_1071 : _T_1082; // @[Mux.scala 31:69:@13425.4]
  assign _T_1084 = _T_1056 ? _T_1069 : _T_1083; // @[Mux.scala 31:69:@13426.4]
  assign _T_1085 = _T_1055 ? _T_1067 : _T_1084; // @[Mux.scala 31:69:@13427.4]
  assign _T_1086 = _T_1054 ? _T_1065 : _T_1085; // @[Mux.scala 31:69:@13428.4]
  assign _T_1087 = _T_1053 ? _T_1063 : _T_1086; // @[Mux.scala 31:69:@13429.4]
  assign _T_1095 = _T_1000 & _T_542; // @[MemPrimitives.scala 110:228:@13438.4]
  assign _T_1101 = _T_1006 & _T_548; // @[MemPrimitives.scala 110:228:@13442.4]
  assign _T_1107 = _T_1012 & _T_554; // @[MemPrimitives.scala 110:228:@13446.4]
  assign _T_1113 = _T_1018 & _T_560; // @[MemPrimitives.scala 110:228:@13450.4]
  assign _T_1119 = _T_1024 & _T_566; // @[MemPrimitives.scala 110:228:@13454.4]
  assign _T_1125 = _T_1030 & _T_572; // @[MemPrimitives.scala 110:228:@13458.4]
  assign _T_1131 = _T_1036 & _T_578; // @[MemPrimitives.scala 110:228:@13462.4]
  assign _T_1137 = _T_1042 & _T_584; // @[MemPrimitives.scala 110:228:@13466.4]
  assign _T_1143 = _T_1048 & _T_590; // @[MemPrimitives.scala 110:228:@13470.4]
  assign _T_1145 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@13484.4]
  assign _T_1146 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@13485.4]
  assign _T_1147 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@13486.4]
  assign _T_1148 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@13487.4]
  assign _T_1149 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 126:35:@13488.4]
  assign _T_1150 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 126:35:@13489.4]
  assign _T_1151 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 126:35:@13490.4]
  assign _T_1152 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 126:35:@13491.4]
  assign _T_1153 = StickySelects_7_io_outs_8; // @[MemPrimitives.scala 126:35:@13492.4]
  assign _T_1155 = {_T_1145,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13494.4]
  assign _T_1157 = {_T_1146,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13496.4]
  assign _T_1159 = {_T_1147,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13498.4]
  assign _T_1161 = {_T_1148,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13500.4]
  assign _T_1163 = {_T_1149,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13502.4]
  assign _T_1165 = {_T_1150,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13504.4]
  assign _T_1167 = {_T_1151,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13506.4]
  assign _T_1169 = {_T_1152,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13508.4]
  assign _T_1171 = {_T_1153,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13510.4]
  assign _T_1172 = _T_1152 ? _T_1169 : _T_1171; // @[Mux.scala 31:69:@13511.4]
  assign _T_1173 = _T_1151 ? _T_1167 : _T_1172; // @[Mux.scala 31:69:@13512.4]
  assign _T_1174 = _T_1150 ? _T_1165 : _T_1173; // @[Mux.scala 31:69:@13513.4]
  assign _T_1175 = _T_1149 ? _T_1163 : _T_1174; // @[Mux.scala 31:69:@13514.4]
  assign _T_1176 = _T_1148 ? _T_1161 : _T_1175; // @[Mux.scala 31:69:@13515.4]
  assign _T_1177 = _T_1147 ? _T_1159 : _T_1176; // @[Mux.scala 31:69:@13516.4]
  assign _T_1178 = _T_1146 ? _T_1157 : _T_1177; // @[Mux.scala 31:69:@13517.4]
  assign _T_1179 = _T_1145 ? _T_1155 : _T_1178; // @[Mux.scala 31:69:@13518.4]
  assign _T_1187 = _T_1000 & _T_634; // @[MemPrimitives.scala 110:228:@13527.4]
  assign _T_1193 = _T_1006 & _T_640; // @[MemPrimitives.scala 110:228:@13531.4]
  assign _T_1199 = _T_1012 & _T_646; // @[MemPrimitives.scala 110:228:@13535.4]
  assign _T_1205 = _T_1018 & _T_652; // @[MemPrimitives.scala 110:228:@13539.4]
  assign _T_1211 = _T_1024 & _T_658; // @[MemPrimitives.scala 110:228:@13543.4]
  assign _T_1217 = _T_1030 & _T_664; // @[MemPrimitives.scala 110:228:@13547.4]
  assign _T_1223 = _T_1036 & _T_670; // @[MemPrimitives.scala 110:228:@13551.4]
  assign _T_1229 = _T_1042 & _T_676; // @[MemPrimitives.scala 110:228:@13555.4]
  assign _T_1235 = _T_1048 & _T_682; // @[MemPrimitives.scala 110:228:@13559.4]
  assign _T_1237 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@13573.4]
  assign _T_1238 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@13574.4]
  assign _T_1239 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 126:35:@13575.4]
  assign _T_1240 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 126:35:@13576.4]
  assign _T_1241 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 126:35:@13577.4]
  assign _T_1242 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 126:35:@13578.4]
  assign _T_1243 = StickySelects_8_io_outs_6; // @[MemPrimitives.scala 126:35:@13579.4]
  assign _T_1244 = StickySelects_8_io_outs_7; // @[MemPrimitives.scala 126:35:@13580.4]
  assign _T_1245 = StickySelects_8_io_outs_8; // @[MemPrimitives.scala 126:35:@13581.4]
  assign _T_1247 = {_T_1237,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13583.4]
  assign _T_1249 = {_T_1238,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13585.4]
  assign _T_1251 = {_T_1239,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13587.4]
  assign _T_1253 = {_T_1240,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13589.4]
  assign _T_1255 = {_T_1241,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13591.4]
  assign _T_1257 = {_T_1242,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13593.4]
  assign _T_1259 = {_T_1243,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13595.4]
  assign _T_1261 = {_T_1244,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13597.4]
  assign _T_1263 = {_T_1245,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13599.4]
  assign _T_1264 = _T_1244 ? _T_1261 : _T_1263; // @[Mux.scala 31:69:@13600.4]
  assign _T_1265 = _T_1243 ? _T_1259 : _T_1264; // @[Mux.scala 31:69:@13601.4]
  assign _T_1266 = _T_1242 ? _T_1257 : _T_1265; // @[Mux.scala 31:69:@13602.4]
  assign _T_1267 = _T_1241 ? _T_1255 : _T_1266; // @[Mux.scala 31:69:@13603.4]
  assign _T_1268 = _T_1240 ? _T_1253 : _T_1267; // @[Mux.scala 31:69:@13604.4]
  assign _T_1269 = _T_1239 ? _T_1251 : _T_1268; // @[Mux.scala 31:69:@13605.4]
  assign _T_1270 = _T_1238 ? _T_1249 : _T_1269; // @[Mux.scala 31:69:@13606.4]
  assign _T_1271 = _T_1237 ? _T_1247 : _T_1270; // @[Mux.scala 31:69:@13607.4]
  assign _T_1276 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13614.4]
  assign _T_1279 = _T_1276 & _T_450; // @[MemPrimitives.scala 110:228:@13616.4]
  assign _T_1282 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13618.4]
  assign _T_1285 = _T_1282 & _T_456; // @[MemPrimitives.scala 110:228:@13620.4]
  assign _T_1288 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13622.4]
  assign _T_1291 = _T_1288 & _T_462; // @[MemPrimitives.scala 110:228:@13624.4]
  assign _T_1294 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13626.4]
  assign _T_1297 = _T_1294 & _T_468; // @[MemPrimitives.scala 110:228:@13628.4]
  assign _T_1300 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13630.4]
  assign _T_1303 = _T_1300 & _T_474; // @[MemPrimitives.scala 110:228:@13632.4]
  assign _T_1306 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13634.4]
  assign _T_1309 = _T_1306 & _T_480; // @[MemPrimitives.scala 110:228:@13636.4]
  assign _T_1312 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13638.4]
  assign _T_1315 = _T_1312 & _T_486; // @[MemPrimitives.scala 110:228:@13640.4]
  assign _T_1318 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13642.4]
  assign _T_1321 = _T_1318 & _T_492; // @[MemPrimitives.scala 110:228:@13644.4]
  assign _T_1324 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13646.4]
  assign _T_1327 = _T_1324 & _T_498; // @[MemPrimitives.scala 110:228:@13648.4]
  assign _T_1329 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@13662.4]
  assign _T_1330 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@13663.4]
  assign _T_1331 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@13664.4]
  assign _T_1332 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@13665.4]
  assign _T_1333 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 126:35:@13666.4]
  assign _T_1334 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 126:35:@13667.4]
  assign _T_1335 = StickySelects_9_io_outs_6; // @[MemPrimitives.scala 126:35:@13668.4]
  assign _T_1336 = StickySelects_9_io_outs_7; // @[MemPrimitives.scala 126:35:@13669.4]
  assign _T_1337 = StickySelects_9_io_outs_8; // @[MemPrimitives.scala 126:35:@13670.4]
  assign _T_1339 = {_T_1329,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13672.4]
  assign _T_1341 = {_T_1330,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13674.4]
  assign _T_1343 = {_T_1331,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13676.4]
  assign _T_1345 = {_T_1332,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13678.4]
  assign _T_1347 = {_T_1333,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13680.4]
  assign _T_1349 = {_T_1334,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13682.4]
  assign _T_1351 = {_T_1335,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13684.4]
  assign _T_1353 = {_T_1336,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13686.4]
  assign _T_1355 = {_T_1337,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13688.4]
  assign _T_1356 = _T_1336 ? _T_1353 : _T_1355; // @[Mux.scala 31:69:@13689.4]
  assign _T_1357 = _T_1335 ? _T_1351 : _T_1356; // @[Mux.scala 31:69:@13690.4]
  assign _T_1358 = _T_1334 ? _T_1349 : _T_1357; // @[Mux.scala 31:69:@13691.4]
  assign _T_1359 = _T_1333 ? _T_1347 : _T_1358; // @[Mux.scala 31:69:@13692.4]
  assign _T_1360 = _T_1332 ? _T_1345 : _T_1359; // @[Mux.scala 31:69:@13693.4]
  assign _T_1361 = _T_1331 ? _T_1343 : _T_1360; // @[Mux.scala 31:69:@13694.4]
  assign _T_1362 = _T_1330 ? _T_1341 : _T_1361; // @[Mux.scala 31:69:@13695.4]
  assign _T_1363 = _T_1329 ? _T_1339 : _T_1362; // @[Mux.scala 31:69:@13696.4]
  assign _T_1371 = _T_1276 & _T_542; // @[MemPrimitives.scala 110:228:@13705.4]
  assign _T_1377 = _T_1282 & _T_548; // @[MemPrimitives.scala 110:228:@13709.4]
  assign _T_1383 = _T_1288 & _T_554; // @[MemPrimitives.scala 110:228:@13713.4]
  assign _T_1389 = _T_1294 & _T_560; // @[MemPrimitives.scala 110:228:@13717.4]
  assign _T_1395 = _T_1300 & _T_566; // @[MemPrimitives.scala 110:228:@13721.4]
  assign _T_1401 = _T_1306 & _T_572; // @[MemPrimitives.scala 110:228:@13725.4]
  assign _T_1407 = _T_1312 & _T_578; // @[MemPrimitives.scala 110:228:@13729.4]
  assign _T_1413 = _T_1318 & _T_584; // @[MemPrimitives.scala 110:228:@13733.4]
  assign _T_1419 = _T_1324 & _T_590; // @[MemPrimitives.scala 110:228:@13737.4]
  assign _T_1421 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@13751.4]
  assign _T_1422 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@13752.4]
  assign _T_1423 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 126:35:@13753.4]
  assign _T_1424 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 126:35:@13754.4]
  assign _T_1425 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 126:35:@13755.4]
  assign _T_1426 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 126:35:@13756.4]
  assign _T_1427 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 126:35:@13757.4]
  assign _T_1428 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 126:35:@13758.4]
  assign _T_1429 = StickySelects_10_io_outs_8; // @[MemPrimitives.scala 126:35:@13759.4]
  assign _T_1431 = {_T_1421,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13761.4]
  assign _T_1433 = {_T_1422,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13763.4]
  assign _T_1435 = {_T_1423,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13765.4]
  assign _T_1437 = {_T_1424,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13767.4]
  assign _T_1439 = {_T_1425,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13769.4]
  assign _T_1441 = {_T_1426,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13771.4]
  assign _T_1443 = {_T_1427,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13773.4]
  assign _T_1445 = {_T_1428,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13775.4]
  assign _T_1447 = {_T_1429,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13777.4]
  assign _T_1448 = _T_1428 ? _T_1445 : _T_1447; // @[Mux.scala 31:69:@13778.4]
  assign _T_1449 = _T_1427 ? _T_1443 : _T_1448; // @[Mux.scala 31:69:@13779.4]
  assign _T_1450 = _T_1426 ? _T_1441 : _T_1449; // @[Mux.scala 31:69:@13780.4]
  assign _T_1451 = _T_1425 ? _T_1439 : _T_1450; // @[Mux.scala 31:69:@13781.4]
  assign _T_1452 = _T_1424 ? _T_1437 : _T_1451; // @[Mux.scala 31:69:@13782.4]
  assign _T_1453 = _T_1423 ? _T_1435 : _T_1452; // @[Mux.scala 31:69:@13783.4]
  assign _T_1454 = _T_1422 ? _T_1433 : _T_1453; // @[Mux.scala 31:69:@13784.4]
  assign _T_1455 = _T_1421 ? _T_1431 : _T_1454; // @[Mux.scala 31:69:@13785.4]
  assign _T_1463 = _T_1276 & _T_634; // @[MemPrimitives.scala 110:228:@13794.4]
  assign _T_1469 = _T_1282 & _T_640; // @[MemPrimitives.scala 110:228:@13798.4]
  assign _T_1475 = _T_1288 & _T_646; // @[MemPrimitives.scala 110:228:@13802.4]
  assign _T_1481 = _T_1294 & _T_652; // @[MemPrimitives.scala 110:228:@13806.4]
  assign _T_1487 = _T_1300 & _T_658; // @[MemPrimitives.scala 110:228:@13810.4]
  assign _T_1493 = _T_1306 & _T_664; // @[MemPrimitives.scala 110:228:@13814.4]
  assign _T_1499 = _T_1312 & _T_670; // @[MemPrimitives.scala 110:228:@13818.4]
  assign _T_1505 = _T_1318 & _T_676; // @[MemPrimitives.scala 110:228:@13822.4]
  assign _T_1511 = _T_1324 & _T_682; // @[MemPrimitives.scala 110:228:@13826.4]
  assign _T_1513 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@13840.4]
  assign _T_1514 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@13841.4]
  assign _T_1515 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@13842.4]
  assign _T_1516 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@13843.4]
  assign _T_1517 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 126:35:@13844.4]
  assign _T_1518 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 126:35:@13845.4]
  assign _T_1519 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 126:35:@13846.4]
  assign _T_1520 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 126:35:@13847.4]
  assign _T_1521 = StickySelects_11_io_outs_8; // @[MemPrimitives.scala 126:35:@13848.4]
  assign _T_1523 = {_T_1513,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13850.4]
  assign _T_1525 = {_T_1514,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13852.4]
  assign _T_1527 = {_T_1515,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13854.4]
  assign _T_1529 = {_T_1516,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13856.4]
  assign _T_1531 = {_T_1517,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13858.4]
  assign _T_1533 = {_T_1518,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13860.4]
  assign _T_1535 = {_T_1519,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13862.4]
  assign _T_1537 = {_T_1520,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13864.4]
  assign _T_1539 = {_T_1521,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13866.4]
  assign _T_1540 = _T_1520 ? _T_1537 : _T_1539; // @[Mux.scala 31:69:@13867.4]
  assign _T_1541 = _T_1519 ? _T_1535 : _T_1540; // @[Mux.scala 31:69:@13868.4]
  assign _T_1542 = _T_1518 ? _T_1533 : _T_1541; // @[Mux.scala 31:69:@13869.4]
  assign _T_1543 = _T_1517 ? _T_1531 : _T_1542; // @[Mux.scala 31:69:@13870.4]
  assign _T_1544 = _T_1516 ? _T_1529 : _T_1543; // @[Mux.scala 31:69:@13871.4]
  assign _T_1545 = _T_1515 ? _T_1527 : _T_1544; // @[Mux.scala 31:69:@13872.4]
  assign _T_1546 = _T_1514 ? _T_1525 : _T_1545; // @[Mux.scala 31:69:@13873.4]
  assign _T_1547 = _T_1513 ? _T_1523 : _T_1546; // @[Mux.scala 31:69:@13874.4]
  assign _T_1643 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@14003.4 package.scala 96:25:@14004.4]
  assign _T_1647 = _T_1643 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14013.4]
  assign _T_1640 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@13995.4 package.scala 96:25:@13996.4]
  assign _T_1648 = _T_1640 ? Mem1D_9_io_output : _T_1647; // @[Mux.scala 31:69:@14014.4]
  assign _T_1637 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@13987.4 package.scala 96:25:@13988.4]
  assign _T_1649 = _T_1637 ? Mem1D_8_io_output : _T_1648; // @[Mux.scala 31:69:@14015.4]
  assign _T_1634 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@13979.4 package.scala 96:25:@13980.4]
  assign _T_1650 = _T_1634 ? Mem1D_7_io_output : _T_1649; // @[Mux.scala 31:69:@14016.4]
  assign _T_1631 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@13971.4 package.scala 96:25:@13972.4]
  assign _T_1651 = _T_1631 ? Mem1D_6_io_output : _T_1650; // @[Mux.scala 31:69:@14017.4]
  assign _T_1628 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@13963.4 package.scala 96:25:@13964.4]
  assign _T_1652 = _T_1628 ? Mem1D_5_io_output : _T_1651; // @[Mux.scala 31:69:@14018.4]
  assign _T_1625 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@13955.4 package.scala 96:25:@13956.4]
  assign _T_1653 = _T_1625 ? Mem1D_4_io_output : _T_1652; // @[Mux.scala 31:69:@14019.4]
  assign _T_1622 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@13947.4 package.scala 96:25:@13948.4]
  assign _T_1654 = _T_1622 ? Mem1D_3_io_output : _T_1653; // @[Mux.scala 31:69:@14020.4]
  assign _T_1619 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@13939.4 package.scala 96:25:@13940.4]
  assign _T_1655 = _T_1619 ? Mem1D_2_io_output : _T_1654; // @[Mux.scala 31:69:@14021.4]
  assign _T_1616 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@13931.4 package.scala 96:25:@13932.4]
  assign _T_1656 = _T_1616 ? Mem1D_1_io_output : _T_1655; // @[Mux.scala 31:69:@14022.4]
  assign _T_1613 = RetimeWrapper_io_out; // @[package.scala 96:25:@13923.4 package.scala 96:25:@13924.4]
  assign _T_1750 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@14147.4 package.scala 96:25:@14148.4]
  assign _T_1754 = _T_1750 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14157.4]
  assign _T_1747 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@14139.4 package.scala 96:25:@14140.4]
  assign _T_1755 = _T_1747 ? Mem1D_9_io_output : _T_1754; // @[Mux.scala 31:69:@14158.4]
  assign _T_1744 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@14131.4 package.scala 96:25:@14132.4]
  assign _T_1756 = _T_1744 ? Mem1D_8_io_output : _T_1755; // @[Mux.scala 31:69:@14159.4]
  assign _T_1741 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@14123.4 package.scala 96:25:@14124.4]
  assign _T_1757 = _T_1741 ? Mem1D_7_io_output : _T_1756; // @[Mux.scala 31:69:@14160.4]
  assign _T_1738 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@14115.4 package.scala 96:25:@14116.4]
  assign _T_1758 = _T_1738 ? Mem1D_6_io_output : _T_1757; // @[Mux.scala 31:69:@14161.4]
  assign _T_1735 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@14107.4 package.scala 96:25:@14108.4]
  assign _T_1759 = _T_1735 ? Mem1D_5_io_output : _T_1758; // @[Mux.scala 31:69:@14162.4]
  assign _T_1732 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@14099.4 package.scala 96:25:@14100.4]
  assign _T_1760 = _T_1732 ? Mem1D_4_io_output : _T_1759; // @[Mux.scala 31:69:@14163.4]
  assign _T_1729 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@14091.4 package.scala 96:25:@14092.4]
  assign _T_1761 = _T_1729 ? Mem1D_3_io_output : _T_1760; // @[Mux.scala 31:69:@14164.4]
  assign _T_1726 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@14083.4 package.scala 96:25:@14084.4]
  assign _T_1762 = _T_1726 ? Mem1D_2_io_output : _T_1761; // @[Mux.scala 31:69:@14165.4]
  assign _T_1723 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@14075.4 package.scala 96:25:@14076.4]
  assign _T_1763 = _T_1723 ? Mem1D_1_io_output : _T_1762; // @[Mux.scala 31:69:@14166.4]
  assign _T_1720 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@14067.4 package.scala 96:25:@14068.4]
  assign _T_1857 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@14291.4 package.scala 96:25:@14292.4]
  assign _T_1861 = _T_1857 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14301.4]
  assign _T_1854 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@14283.4 package.scala 96:25:@14284.4]
  assign _T_1862 = _T_1854 ? Mem1D_9_io_output : _T_1861; // @[Mux.scala 31:69:@14302.4]
  assign _T_1851 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@14275.4 package.scala 96:25:@14276.4]
  assign _T_1863 = _T_1851 ? Mem1D_8_io_output : _T_1862; // @[Mux.scala 31:69:@14303.4]
  assign _T_1848 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@14267.4 package.scala 96:25:@14268.4]
  assign _T_1864 = _T_1848 ? Mem1D_7_io_output : _T_1863; // @[Mux.scala 31:69:@14304.4]
  assign _T_1845 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@14259.4 package.scala 96:25:@14260.4]
  assign _T_1865 = _T_1845 ? Mem1D_6_io_output : _T_1864; // @[Mux.scala 31:69:@14305.4]
  assign _T_1842 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@14251.4 package.scala 96:25:@14252.4]
  assign _T_1866 = _T_1842 ? Mem1D_5_io_output : _T_1865; // @[Mux.scala 31:69:@14306.4]
  assign _T_1839 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@14243.4 package.scala 96:25:@14244.4]
  assign _T_1867 = _T_1839 ? Mem1D_4_io_output : _T_1866; // @[Mux.scala 31:69:@14307.4]
  assign _T_1836 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@14235.4 package.scala 96:25:@14236.4]
  assign _T_1868 = _T_1836 ? Mem1D_3_io_output : _T_1867; // @[Mux.scala 31:69:@14308.4]
  assign _T_1833 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@14227.4 package.scala 96:25:@14228.4]
  assign _T_1869 = _T_1833 ? Mem1D_2_io_output : _T_1868; // @[Mux.scala 31:69:@14309.4]
  assign _T_1830 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@14219.4 package.scala 96:25:@14220.4]
  assign _T_1870 = _T_1830 ? Mem1D_1_io_output : _T_1869; // @[Mux.scala 31:69:@14310.4]
  assign _T_1827 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@14211.4 package.scala 96:25:@14212.4]
  assign _T_1964 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@14435.4 package.scala 96:25:@14436.4]
  assign _T_1968 = _T_1964 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14445.4]
  assign _T_1961 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@14427.4 package.scala 96:25:@14428.4]
  assign _T_1969 = _T_1961 ? Mem1D_9_io_output : _T_1968; // @[Mux.scala 31:69:@14446.4]
  assign _T_1958 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@14419.4 package.scala 96:25:@14420.4]
  assign _T_1970 = _T_1958 ? Mem1D_8_io_output : _T_1969; // @[Mux.scala 31:69:@14447.4]
  assign _T_1955 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@14411.4 package.scala 96:25:@14412.4]
  assign _T_1971 = _T_1955 ? Mem1D_7_io_output : _T_1970; // @[Mux.scala 31:69:@14448.4]
  assign _T_1952 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@14403.4 package.scala 96:25:@14404.4]
  assign _T_1972 = _T_1952 ? Mem1D_6_io_output : _T_1971; // @[Mux.scala 31:69:@14449.4]
  assign _T_1949 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@14395.4 package.scala 96:25:@14396.4]
  assign _T_1973 = _T_1949 ? Mem1D_5_io_output : _T_1972; // @[Mux.scala 31:69:@14450.4]
  assign _T_1946 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@14387.4 package.scala 96:25:@14388.4]
  assign _T_1974 = _T_1946 ? Mem1D_4_io_output : _T_1973; // @[Mux.scala 31:69:@14451.4]
  assign _T_1943 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@14379.4 package.scala 96:25:@14380.4]
  assign _T_1975 = _T_1943 ? Mem1D_3_io_output : _T_1974; // @[Mux.scala 31:69:@14452.4]
  assign _T_1940 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@14371.4 package.scala 96:25:@14372.4]
  assign _T_1976 = _T_1940 ? Mem1D_2_io_output : _T_1975; // @[Mux.scala 31:69:@14453.4]
  assign _T_1937 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@14363.4 package.scala 96:25:@14364.4]
  assign _T_1977 = _T_1937 ? Mem1D_1_io_output : _T_1976; // @[Mux.scala 31:69:@14454.4]
  assign _T_1934 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@14355.4 package.scala 96:25:@14356.4]
  assign _T_2071 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@14579.4 package.scala 96:25:@14580.4]
  assign _T_2075 = _T_2071 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14589.4]
  assign _T_2068 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@14571.4 package.scala 96:25:@14572.4]
  assign _T_2076 = _T_2068 ? Mem1D_9_io_output : _T_2075; // @[Mux.scala 31:69:@14590.4]
  assign _T_2065 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@14563.4 package.scala 96:25:@14564.4]
  assign _T_2077 = _T_2065 ? Mem1D_8_io_output : _T_2076; // @[Mux.scala 31:69:@14591.4]
  assign _T_2062 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@14555.4 package.scala 96:25:@14556.4]
  assign _T_2078 = _T_2062 ? Mem1D_7_io_output : _T_2077; // @[Mux.scala 31:69:@14592.4]
  assign _T_2059 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@14547.4 package.scala 96:25:@14548.4]
  assign _T_2079 = _T_2059 ? Mem1D_6_io_output : _T_2078; // @[Mux.scala 31:69:@14593.4]
  assign _T_2056 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@14539.4 package.scala 96:25:@14540.4]
  assign _T_2080 = _T_2056 ? Mem1D_5_io_output : _T_2079; // @[Mux.scala 31:69:@14594.4]
  assign _T_2053 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@14531.4 package.scala 96:25:@14532.4]
  assign _T_2081 = _T_2053 ? Mem1D_4_io_output : _T_2080; // @[Mux.scala 31:69:@14595.4]
  assign _T_2050 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@14523.4 package.scala 96:25:@14524.4]
  assign _T_2082 = _T_2050 ? Mem1D_3_io_output : _T_2081; // @[Mux.scala 31:69:@14596.4]
  assign _T_2047 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@14515.4 package.scala 96:25:@14516.4]
  assign _T_2083 = _T_2047 ? Mem1D_2_io_output : _T_2082; // @[Mux.scala 31:69:@14597.4]
  assign _T_2044 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@14507.4 package.scala 96:25:@14508.4]
  assign _T_2084 = _T_2044 ? Mem1D_1_io_output : _T_2083; // @[Mux.scala 31:69:@14598.4]
  assign _T_2041 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@14499.4 package.scala 96:25:@14500.4]
  assign _T_2178 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@14723.4 package.scala 96:25:@14724.4]
  assign _T_2182 = _T_2178 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14733.4]
  assign _T_2175 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@14715.4 package.scala 96:25:@14716.4]
  assign _T_2183 = _T_2175 ? Mem1D_9_io_output : _T_2182; // @[Mux.scala 31:69:@14734.4]
  assign _T_2172 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@14707.4 package.scala 96:25:@14708.4]
  assign _T_2184 = _T_2172 ? Mem1D_8_io_output : _T_2183; // @[Mux.scala 31:69:@14735.4]
  assign _T_2169 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@14699.4 package.scala 96:25:@14700.4]
  assign _T_2185 = _T_2169 ? Mem1D_7_io_output : _T_2184; // @[Mux.scala 31:69:@14736.4]
  assign _T_2166 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@14691.4 package.scala 96:25:@14692.4]
  assign _T_2186 = _T_2166 ? Mem1D_6_io_output : _T_2185; // @[Mux.scala 31:69:@14737.4]
  assign _T_2163 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@14683.4 package.scala 96:25:@14684.4]
  assign _T_2187 = _T_2163 ? Mem1D_5_io_output : _T_2186; // @[Mux.scala 31:69:@14738.4]
  assign _T_2160 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@14675.4 package.scala 96:25:@14676.4]
  assign _T_2188 = _T_2160 ? Mem1D_4_io_output : _T_2187; // @[Mux.scala 31:69:@14739.4]
  assign _T_2157 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@14667.4 package.scala 96:25:@14668.4]
  assign _T_2189 = _T_2157 ? Mem1D_3_io_output : _T_2188; // @[Mux.scala 31:69:@14740.4]
  assign _T_2154 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@14659.4 package.scala 96:25:@14660.4]
  assign _T_2190 = _T_2154 ? Mem1D_2_io_output : _T_2189; // @[Mux.scala 31:69:@14741.4]
  assign _T_2151 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@14651.4 package.scala 96:25:@14652.4]
  assign _T_2191 = _T_2151 ? Mem1D_1_io_output : _T_2190; // @[Mux.scala 31:69:@14742.4]
  assign _T_2148 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@14643.4 package.scala 96:25:@14644.4]
  assign _T_2285 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@14867.4 package.scala 96:25:@14868.4]
  assign _T_2289 = _T_2285 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14877.4]
  assign _T_2282 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@14859.4 package.scala 96:25:@14860.4]
  assign _T_2290 = _T_2282 ? Mem1D_9_io_output : _T_2289; // @[Mux.scala 31:69:@14878.4]
  assign _T_2279 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@14851.4 package.scala 96:25:@14852.4]
  assign _T_2291 = _T_2279 ? Mem1D_8_io_output : _T_2290; // @[Mux.scala 31:69:@14879.4]
  assign _T_2276 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@14843.4 package.scala 96:25:@14844.4]
  assign _T_2292 = _T_2276 ? Mem1D_7_io_output : _T_2291; // @[Mux.scala 31:69:@14880.4]
  assign _T_2273 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@14835.4 package.scala 96:25:@14836.4]
  assign _T_2293 = _T_2273 ? Mem1D_6_io_output : _T_2292; // @[Mux.scala 31:69:@14881.4]
  assign _T_2270 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@14827.4 package.scala 96:25:@14828.4]
  assign _T_2294 = _T_2270 ? Mem1D_5_io_output : _T_2293; // @[Mux.scala 31:69:@14882.4]
  assign _T_2267 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@14819.4 package.scala 96:25:@14820.4]
  assign _T_2295 = _T_2267 ? Mem1D_4_io_output : _T_2294; // @[Mux.scala 31:69:@14883.4]
  assign _T_2264 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@14811.4 package.scala 96:25:@14812.4]
  assign _T_2296 = _T_2264 ? Mem1D_3_io_output : _T_2295; // @[Mux.scala 31:69:@14884.4]
  assign _T_2261 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@14803.4 package.scala 96:25:@14804.4]
  assign _T_2297 = _T_2261 ? Mem1D_2_io_output : _T_2296; // @[Mux.scala 31:69:@14885.4]
  assign _T_2258 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@14795.4 package.scala 96:25:@14796.4]
  assign _T_2298 = _T_2258 ? Mem1D_1_io_output : _T_2297; // @[Mux.scala 31:69:@14886.4]
  assign _T_2255 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@14787.4 package.scala 96:25:@14788.4]
  assign _T_2392 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@15011.4 package.scala 96:25:@15012.4]
  assign _T_2396 = _T_2392 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@15021.4]
  assign _T_2389 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@15003.4 package.scala 96:25:@15004.4]
  assign _T_2397 = _T_2389 ? Mem1D_9_io_output : _T_2396; // @[Mux.scala 31:69:@15022.4]
  assign _T_2386 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@14995.4 package.scala 96:25:@14996.4]
  assign _T_2398 = _T_2386 ? Mem1D_8_io_output : _T_2397; // @[Mux.scala 31:69:@15023.4]
  assign _T_2383 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@14987.4 package.scala 96:25:@14988.4]
  assign _T_2399 = _T_2383 ? Mem1D_7_io_output : _T_2398; // @[Mux.scala 31:69:@15024.4]
  assign _T_2380 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@14979.4 package.scala 96:25:@14980.4]
  assign _T_2400 = _T_2380 ? Mem1D_6_io_output : _T_2399; // @[Mux.scala 31:69:@15025.4]
  assign _T_2377 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@14971.4 package.scala 96:25:@14972.4]
  assign _T_2401 = _T_2377 ? Mem1D_5_io_output : _T_2400; // @[Mux.scala 31:69:@15026.4]
  assign _T_2374 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@14963.4 package.scala 96:25:@14964.4]
  assign _T_2402 = _T_2374 ? Mem1D_4_io_output : _T_2401; // @[Mux.scala 31:69:@15027.4]
  assign _T_2371 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@14955.4 package.scala 96:25:@14956.4]
  assign _T_2403 = _T_2371 ? Mem1D_3_io_output : _T_2402; // @[Mux.scala 31:69:@15028.4]
  assign _T_2368 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@14947.4 package.scala 96:25:@14948.4]
  assign _T_2404 = _T_2368 ? Mem1D_2_io_output : _T_2403; // @[Mux.scala 31:69:@15029.4]
  assign _T_2365 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@14939.4 package.scala 96:25:@14940.4]
  assign _T_2405 = _T_2365 ? Mem1D_1_io_output : _T_2404; // @[Mux.scala 31:69:@15030.4]
  assign _T_2362 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@14931.4 package.scala 96:25:@14932.4]
  assign _T_2499 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@15155.4 package.scala 96:25:@15156.4]
  assign _T_2503 = _T_2499 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@15165.4]
  assign _T_2496 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@15147.4 package.scala 96:25:@15148.4]
  assign _T_2504 = _T_2496 ? Mem1D_9_io_output : _T_2503; // @[Mux.scala 31:69:@15166.4]
  assign _T_2493 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@15139.4 package.scala 96:25:@15140.4]
  assign _T_2505 = _T_2493 ? Mem1D_8_io_output : _T_2504; // @[Mux.scala 31:69:@15167.4]
  assign _T_2490 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@15131.4 package.scala 96:25:@15132.4]
  assign _T_2506 = _T_2490 ? Mem1D_7_io_output : _T_2505; // @[Mux.scala 31:69:@15168.4]
  assign _T_2487 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@15123.4 package.scala 96:25:@15124.4]
  assign _T_2507 = _T_2487 ? Mem1D_6_io_output : _T_2506; // @[Mux.scala 31:69:@15169.4]
  assign _T_2484 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@15115.4 package.scala 96:25:@15116.4]
  assign _T_2508 = _T_2484 ? Mem1D_5_io_output : _T_2507; // @[Mux.scala 31:69:@15170.4]
  assign _T_2481 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@15107.4 package.scala 96:25:@15108.4]
  assign _T_2509 = _T_2481 ? Mem1D_4_io_output : _T_2508; // @[Mux.scala 31:69:@15171.4]
  assign _T_2478 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@15099.4 package.scala 96:25:@15100.4]
  assign _T_2510 = _T_2478 ? Mem1D_3_io_output : _T_2509; // @[Mux.scala 31:69:@15172.4]
  assign _T_2475 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@15091.4 package.scala 96:25:@15092.4]
  assign _T_2511 = _T_2475 ? Mem1D_2_io_output : _T_2510; // @[Mux.scala 31:69:@15173.4]
  assign _T_2472 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@15083.4 package.scala 96:25:@15084.4]
  assign _T_2512 = _T_2472 ? Mem1D_1_io_output : _T_2511; // @[Mux.scala 31:69:@15174.4]
  assign _T_2469 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@15075.4 package.scala 96:25:@15076.4]
  assign io_rPort_8_output_0 = _T_2469 ? Mem1D_io_output : _T_2512; // @[MemPrimitives.scala 152:13:@15176.4]
  assign io_rPort_7_output_0 = _T_2362 ? Mem1D_io_output : _T_2405; // @[MemPrimitives.scala 152:13:@15032.4]
  assign io_rPort_6_output_0 = _T_2255 ? Mem1D_io_output : _T_2298; // @[MemPrimitives.scala 152:13:@14888.4]
  assign io_rPort_5_output_0 = _T_2148 ? Mem1D_io_output : _T_2191; // @[MemPrimitives.scala 152:13:@14744.4]
  assign io_rPort_4_output_0 = _T_2041 ? Mem1D_io_output : _T_2084; // @[MemPrimitives.scala 152:13:@14600.4]
  assign io_rPort_3_output_0 = _T_1934 ? Mem1D_io_output : _T_1977; // @[MemPrimitives.scala 152:13:@14456.4]
  assign io_rPort_2_output_0 = _T_1827 ? Mem1D_io_output : _T_1870; // @[MemPrimitives.scala 152:13:@14312.4]
  assign io_rPort_1_output_0 = _T_1720 ? Mem1D_io_output : _T_1763; // @[MemPrimitives.scala 152:13:@14168.4]
  assign io_rPort_0_output_0 = _T_1613 ? Mem1D_io_output : _T_1656; // @[MemPrimitives.scala 152:13:@14024.4]
  assign Mem1D_clock = clock; // @[:@12478.4]
  assign Mem1D_reset = reset; // @[:@12479.4]
  assign Mem1D_io_r_ofs_0 = _T_535[9:0]; // @[MemPrimitives.scala 131:28:@12899.4]
  assign Mem1D_io_r_backpressure = _T_535[10]; // @[MemPrimitives.scala 132:32:@12900.4]
  assign Mem1D_io_w_ofs_0 = _T_322[9:0]; // @[MemPrimitives.scala 94:28:@12678.4]
  assign Mem1D_io_w_data_0 = _T_322[41:10]; // @[MemPrimitives.scala 95:29:@12679.4]
  assign Mem1D_io_w_en_0 = _T_322[42]; // @[MemPrimitives.scala 96:27:@12680.4]
  assign Mem1D_1_clock = clock; // @[:@12494.4]
  assign Mem1D_1_reset = reset; // @[:@12495.4]
  assign Mem1D_1_io_r_ofs_0 = _T_627[9:0]; // @[MemPrimitives.scala 131:28:@12988.4]
  assign Mem1D_1_io_r_backpressure = _T_627[10]; // @[MemPrimitives.scala 132:32:@12989.4]
  assign Mem1D_1_io_w_ofs_0 = _T_333[9:0]; // @[MemPrimitives.scala 94:28:@12690.4]
  assign Mem1D_1_io_w_data_0 = _T_333[41:10]; // @[MemPrimitives.scala 95:29:@12691.4]
  assign Mem1D_1_io_w_en_0 = _T_333[42]; // @[MemPrimitives.scala 96:27:@12692.4]
  assign Mem1D_2_clock = clock; // @[:@12510.4]
  assign Mem1D_2_reset = reset; // @[:@12511.4]
  assign Mem1D_2_io_r_ofs_0 = _T_719[9:0]; // @[MemPrimitives.scala 131:28:@13077.4]
  assign Mem1D_2_io_r_backpressure = _T_719[10]; // @[MemPrimitives.scala 132:32:@13078.4]
  assign Mem1D_2_io_w_ofs_0 = _T_344[9:0]; // @[MemPrimitives.scala 94:28:@12702.4]
  assign Mem1D_2_io_w_data_0 = _T_344[41:10]; // @[MemPrimitives.scala 95:29:@12703.4]
  assign Mem1D_2_io_w_en_0 = _T_344[42]; // @[MemPrimitives.scala 96:27:@12704.4]
  assign Mem1D_3_clock = clock; // @[:@12526.4]
  assign Mem1D_3_reset = reset; // @[:@12527.4]
  assign Mem1D_3_io_r_ofs_0 = _T_811[9:0]; // @[MemPrimitives.scala 131:28:@13166.4]
  assign Mem1D_3_io_r_backpressure = _T_811[10]; // @[MemPrimitives.scala 132:32:@13167.4]
  assign Mem1D_3_io_w_ofs_0 = _T_355[9:0]; // @[MemPrimitives.scala 94:28:@12714.4]
  assign Mem1D_3_io_w_data_0 = _T_355[41:10]; // @[MemPrimitives.scala 95:29:@12715.4]
  assign Mem1D_3_io_w_en_0 = _T_355[42]; // @[MemPrimitives.scala 96:27:@12716.4]
  assign Mem1D_4_clock = clock; // @[:@12542.4]
  assign Mem1D_4_reset = reset; // @[:@12543.4]
  assign Mem1D_4_io_r_ofs_0 = _T_903[9:0]; // @[MemPrimitives.scala 131:28:@13255.4]
  assign Mem1D_4_io_r_backpressure = _T_903[10]; // @[MemPrimitives.scala 132:32:@13256.4]
  assign Mem1D_4_io_w_ofs_0 = _T_366[9:0]; // @[MemPrimitives.scala 94:28:@12726.4]
  assign Mem1D_4_io_w_data_0 = _T_366[41:10]; // @[MemPrimitives.scala 95:29:@12727.4]
  assign Mem1D_4_io_w_en_0 = _T_366[42]; // @[MemPrimitives.scala 96:27:@12728.4]
  assign Mem1D_5_clock = clock; // @[:@12558.4]
  assign Mem1D_5_reset = reset; // @[:@12559.4]
  assign Mem1D_5_io_r_ofs_0 = _T_995[9:0]; // @[MemPrimitives.scala 131:28:@13344.4]
  assign Mem1D_5_io_r_backpressure = _T_995[10]; // @[MemPrimitives.scala 132:32:@13345.4]
  assign Mem1D_5_io_w_ofs_0 = _T_377[9:0]; // @[MemPrimitives.scala 94:28:@12738.4]
  assign Mem1D_5_io_w_data_0 = _T_377[41:10]; // @[MemPrimitives.scala 95:29:@12739.4]
  assign Mem1D_5_io_w_en_0 = _T_377[42]; // @[MemPrimitives.scala 96:27:@12740.4]
  assign Mem1D_6_clock = clock; // @[:@12574.4]
  assign Mem1D_6_reset = reset; // @[:@12575.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1087[9:0]; // @[MemPrimitives.scala 131:28:@13433.4]
  assign Mem1D_6_io_r_backpressure = _T_1087[10]; // @[MemPrimitives.scala 132:32:@13434.4]
  assign Mem1D_6_io_w_ofs_0 = _T_388[9:0]; // @[MemPrimitives.scala 94:28:@12750.4]
  assign Mem1D_6_io_w_data_0 = _T_388[41:10]; // @[MemPrimitives.scala 95:29:@12751.4]
  assign Mem1D_6_io_w_en_0 = _T_388[42]; // @[MemPrimitives.scala 96:27:@12752.4]
  assign Mem1D_7_clock = clock; // @[:@12590.4]
  assign Mem1D_7_reset = reset; // @[:@12591.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1179[9:0]; // @[MemPrimitives.scala 131:28:@13522.4]
  assign Mem1D_7_io_r_backpressure = _T_1179[10]; // @[MemPrimitives.scala 132:32:@13523.4]
  assign Mem1D_7_io_w_ofs_0 = _T_399[9:0]; // @[MemPrimitives.scala 94:28:@12762.4]
  assign Mem1D_7_io_w_data_0 = _T_399[41:10]; // @[MemPrimitives.scala 95:29:@12763.4]
  assign Mem1D_7_io_w_en_0 = _T_399[42]; // @[MemPrimitives.scala 96:27:@12764.4]
  assign Mem1D_8_clock = clock; // @[:@12606.4]
  assign Mem1D_8_reset = reset; // @[:@12607.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1271[9:0]; // @[MemPrimitives.scala 131:28:@13611.4]
  assign Mem1D_8_io_r_backpressure = _T_1271[10]; // @[MemPrimitives.scala 132:32:@13612.4]
  assign Mem1D_8_io_w_ofs_0 = _T_410[9:0]; // @[MemPrimitives.scala 94:28:@12774.4]
  assign Mem1D_8_io_w_data_0 = _T_410[41:10]; // @[MemPrimitives.scala 95:29:@12775.4]
  assign Mem1D_8_io_w_en_0 = _T_410[42]; // @[MemPrimitives.scala 96:27:@12776.4]
  assign Mem1D_9_clock = clock; // @[:@12622.4]
  assign Mem1D_9_reset = reset; // @[:@12623.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1363[9:0]; // @[MemPrimitives.scala 131:28:@13700.4]
  assign Mem1D_9_io_r_backpressure = _T_1363[10]; // @[MemPrimitives.scala 132:32:@13701.4]
  assign Mem1D_9_io_w_ofs_0 = _T_421[9:0]; // @[MemPrimitives.scala 94:28:@12786.4]
  assign Mem1D_9_io_w_data_0 = _T_421[41:10]; // @[MemPrimitives.scala 95:29:@12787.4]
  assign Mem1D_9_io_w_en_0 = _T_421[42]; // @[MemPrimitives.scala 96:27:@12788.4]
  assign Mem1D_10_clock = clock; // @[:@12638.4]
  assign Mem1D_10_reset = reset; // @[:@12639.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1455[9:0]; // @[MemPrimitives.scala 131:28:@13789.4]
  assign Mem1D_10_io_r_backpressure = _T_1455[10]; // @[MemPrimitives.scala 132:32:@13790.4]
  assign Mem1D_10_io_w_ofs_0 = _T_432[9:0]; // @[MemPrimitives.scala 94:28:@12798.4]
  assign Mem1D_10_io_w_data_0 = _T_432[41:10]; // @[MemPrimitives.scala 95:29:@12799.4]
  assign Mem1D_10_io_w_en_0 = _T_432[42]; // @[MemPrimitives.scala 96:27:@12800.4]
  assign Mem1D_11_clock = clock; // @[:@12654.4]
  assign Mem1D_11_reset = reset; // @[:@12655.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1547[9:0]; // @[MemPrimitives.scala 131:28:@13878.4]
  assign Mem1D_11_io_r_backpressure = _T_1547[10]; // @[MemPrimitives.scala 132:32:@13879.4]
  assign Mem1D_11_io_w_ofs_0 = _T_443[9:0]; // @[MemPrimitives.scala 94:28:@12810.4]
  assign Mem1D_11_io_w_data_0 = _T_443[41:10]; // @[MemPrimitives.scala 95:29:@12811.4]
  assign Mem1D_11_io_w_en_0 = _T_443[42]; // @[MemPrimitives.scala 96:27:@12812.4]
  assign StickySelects_clock = clock; // @[:@12850.4]
  assign StickySelects_reset = reset; // @[:@12851.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_451; // @[MemPrimitives.scala 125:64:@12852.4]
  assign StickySelects_io_ins_1 = io_rPort_1_en_0 & _T_457; // @[MemPrimitives.scala 125:64:@12853.4]
  assign StickySelects_io_ins_2 = io_rPort_2_en_0 & _T_463; // @[MemPrimitives.scala 125:64:@12854.4]
  assign StickySelects_io_ins_3 = io_rPort_3_en_0 & _T_469; // @[MemPrimitives.scala 125:64:@12855.4]
  assign StickySelects_io_ins_4 = io_rPort_4_en_0 & _T_475; // @[MemPrimitives.scala 125:64:@12856.4]
  assign StickySelects_io_ins_5 = io_rPort_5_en_0 & _T_481; // @[MemPrimitives.scala 125:64:@12857.4]
  assign StickySelects_io_ins_6 = io_rPort_6_en_0 & _T_487; // @[MemPrimitives.scala 125:64:@12858.4]
  assign StickySelects_io_ins_7 = io_rPort_7_en_0 & _T_493; // @[MemPrimitives.scala 125:64:@12859.4]
  assign StickySelects_io_ins_8 = io_rPort_8_en_0 & _T_499; // @[MemPrimitives.scala 125:64:@12860.4]
  assign StickySelects_1_clock = clock; // @[:@12939.4]
  assign StickySelects_1_reset = reset; // @[:@12940.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_543; // @[MemPrimitives.scala 125:64:@12941.4]
  assign StickySelects_1_io_ins_1 = io_rPort_1_en_0 & _T_549; // @[MemPrimitives.scala 125:64:@12942.4]
  assign StickySelects_1_io_ins_2 = io_rPort_2_en_0 & _T_555; // @[MemPrimitives.scala 125:64:@12943.4]
  assign StickySelects_1_io_ins_3 = io_rPort_3_en_0 & _T_561; // @[MemPrimitives.scala 125:64:@12944.4]
  assign StickySelects_1_io_ins_4 = io_rPort_4_en_0 & _T_567; // @[MemPrimitives.scala 125:64:@12945.4]
  assign StickySelects_1_io_ins_5 = io_rPort_5_en_0 & _T_573; // @[MemPrimitives.scala 125:64:@12946.4]
  assign StickySelects_1_io_ins_6 = io_rPort_6_en_0 & _T_579; // @[MemPrimitives.scala 125:64:@12947.4]
  assign StickySelects_1_io_ins_7 = io_rPort_7_en_0 & _T_585; // @[MemPrimitives.scala 125:64:@12948.4]
  assign StickySelects_1_io_ins_8 = io_rPort_8_en_0 & _T_591; // @[MemPrimitives.scala 125:64:@12949.4]
  assign StickySelects_2_clock = clock; // @[:@13028.4]
  assign StickySelects_2_reset = reset; // @[:@13029.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_635; // @[MemPrimitives.scala 125:64:@13030.4]
  assign StickySelects_2_io_ins_1 = io_rPort_1_en_0 & _T_641; // @[MemPrimitives.scala 125:64:@13031.4]
  assign StickySelects_2_io_ins_2 = io_rPort_2_en_0 & _T_647; // @[MemPrimitives.scala 125:64:@13032.4]
  assign StickySelects_2_io_ins_3 = io_rPort_3_en_0 & _T_653; // @[MemPrimitives.scala 125:64:@13033.4]
  assign StickySelects_2_io_ins_4 = io_rPort_4_en_0 & _T_659; // @[MemPrimitives.scala 125:64:@13034.4]
  assign StickySelects_2_io_ins_5 = io_rPort_5_en_0 & _T_665; // @[MemPrimitives.scala 125:64:@13035.4]
  assign StickySelects_2_io_ins_6 = io_rPort_6_en_0 & _T_671; // @[MemPrimitives.scala 125:64:@13036.4]
  assign StickySelects_2_io_ins_7 = io_rPort_7_en_0 & _T_677; // @[MemPrimitives.scala 125:64:@13037.4]
  assign StickySelects_2_io_ins_8 = io_rPort_8_en_0 & _T_683; // @[MemPrimitives.scala 125:64:@13038.4]
  assign StickySelects_3_clock = clock; // @[:@13117.4]
  assign StickySelects_3_reset = reset; // @[:@13118.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_727; // @[MemPrimitives.scala 125:64:@13119.4]
  assign StickySelects_3_io_ins_1 = io_rPort_1_en_0 & _T_733; // @[MemPrimitives.scala 125:64:@13120.4]
  assign StickySelects_3_io_ins_2 = io_rPort_2_en_0 & _T_739; // @[MemPrimitives.scala 125:64:@13121.4]
  assign StickySelects_3_io_ins_3 = io_rPort_3_en_0 & _T_745; // @[MemPrimitives.scala 125:64:@13122.4]
  assign StickySelects_3_io_ins_4 = io_rPort_4_en_0 & _T_751; // @[MemPrimitives.scala 125:64:@13123.4]
  assign StickySelects_3_io_ins_5 = io_rPort_5_en_0 & _T_757; // @[MemPrimitives.scala 125:64:@13124.4]
  assign StickySelects_3_io_ins_6 = io_rPort_6_en_0 & _T_763; // @[MemPrimitives.scala 125:64:@13125.4]
  assign StickySelects_3_io_ins_7 = io_rPort_7_en_0 & _T_769; // @[MemPrimitives.scala 125:64:@13126.4]
  assign StickySelects_3_io_ins_8 = io_rPort_8_en_0 & _T_775; // @[MemPrimitives.scala 125:64:@13127.4]
  assign StickySelects_4_clock = clock; // @[:@13206.4]
  assign StickySelects_4_reset = reset; // @[:@13207.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_819; // @[MemPrimitives.scala 125:64:@13208.4]
  assign StickySelects_4_io_ins_1 = io_rPort_1_en_0 & _T_825; // @[MemPrimitives.scala 125:64:@13209.4]
  assign StickySelects_4_io_ins_2 = io_rPort_2_en_0 & _T_831; // @[MemPrimitives.scala 125:64:@13210.4]
  assign StickySelects_4_io_ins_3 = io_rPort_3_en_0 & _T_837; // @[MemPrimitives.scala 125:64:@13211.4]
  assign StickySelects_4_io_ins_4 = io_rPort_4_en_0 & _T_843; // @[MemPrimitives.scala 125:64:@13212.4]
  assign StickySelects_4_io_ins_5 = io_rPort_5_en_0 & _T_849; // @[MemPrimitives.scala 125:64:@13213.4]
  assign StickySelects_4_io_ins_6 = io_rPort_6_en_0 & _T_855; // @[MemPrimitives.scala 125:64:@13214.4]
  assign StickySelects_4_io_ins_7 = io_rPort_7_en_0 & _T_861; // @[MemPrimitives.scala 125:64:@13215.4]
  assign StickySelects_4_io_ins_8 = io_rPort_8_en_0 & _T_867; // @[MemPrimitives.scala 125:64:@13216.4]
  assign StickySelects_5_clock = clock; // @[:@13295.4]
  assign StickySelects_5_reset = reset; // @[:@13296.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_911; // @[MemPrimitives.scala 125:64:@13297.4]
  assign StickySelects_5_io_ins_1 = io_rPort_1_en_0 & _T_917; // @[MemPrimitives.scala 125:64:@13298.4]
  assign StickySelects_5_io_ins_2 = io_rPort_2_en_0 & _T_923; // @[MemPrimitives.scala 125:64:@13299.4]
  assign StickySelects_5_io_ins_3 = io_rPort_3_en_0 & _T_929; // @[MemPrimitives.scala 125:64:@13300.4]
  assign StickySelects_5_io_ins_4 = io_rPort_4_en_0 & _T_935; // @[MemPrimitives.scala 125:64:@13301.4]
  assign StickySelects_5_io_ins_5 = io_rPort_5_en_0 & _T_941; // @[MemPrimitives.scala 125:64:@13302.4]
  assign StickySelects_5_io_ins_6 = io_rPort_6_en_0 & _T_947; // @[MemPrimitives.scala 125:64:@13303.4]
  assign StickySelects_5_io_ins_7 = io_rPort_7_en_0 & _T_953; // @[MemPrimitives.scala 125:64:@13304.4]
  assign StickySelects_5_io_ins_8 = io_rPort_8_en_0 & _T_959; // @[MemPrimitives.scala 125:64:@13305.4]
  assign StickySelects_6_clock = clock; // @[:@13384.4]
  assign StickySelects_6_reset = reset; // @[:@13385.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_1003; // @[MemPrimitives.scala 125:64:@13386.4]
  assign StickySelects_6_io_ins_1 = io_rPort_1_en_0 & _T_1009; // @[MemPrimitives.scala 125:64:@13387.4]
  assign StickySelects_6_io_ins_2 = io_rPort_2_en_0 & _T_1015; // @[MemPrimitives.scala 125:64:@13388.4]
  assign StickySelects_6_io_ins_3 = io_rPort_3_en_0 & _T_1021; // @[MemPrimitives.scala 125:64:@13389.4]
  assign StickySelects_6_io_ins_4 = io_rPort_4_en_0 & _T_1027; // @[MemPrimitives.scala 125:64:@13390.4]
  assign StickySelects_6_io_ins_5 = io_rPort_5_en_0 & _T_1033; // @[MemPrimitives.scala 125:64:@13391.4]
  assign StickySelects_6_io_ins_6 = io_rPort_6_en_0 & _T_1039; // @[MemPrimitives.scala 125:64:@13392.4]
  assign StickySelects_6_io_ins_7 = io_rPort_7_en_0 & _T_1045; // @[MemPrimitives.scala 125:64:@13393.4]
  assign StickySelects_6_io_ins_8 = io_rPort_8_en_0 & _T_1051; // @[MemPrimitives.scala 125:64:@13394.4]
  assign StickySelects_7_clock = clock; // @[:@13473.4]
  assign StickySelects_7_reset = reset; // @[:@13474.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1095; // @[MemPrimitives.scala 125:64:@13475.4]
  assign StickySelects_7_io_ins_1 = io_rPort_1_en_0 & _T_1101; // @[MemPrimitives.scala 125:64:@13476.4]
  assign StickySelects_7_io_ins_2 = io_rPort_2_en_0 & _T_1107; // @[MemPrimitives.scala 125:64:@13477.4]
  assign StickySelects_7_io_ins_3 = io_rPort_3_en_0 & _T_1113; // @[MemPrimitives.scala 125:64:@13478.4]
  assign StickySelects_7_io_ins_4 = io_rPort_4_en_0 & _T_1119; // @[MemPrimitives.scala 125:64:@13479.4]
  assign StickySelects_7_io_ins_5 = io_rPort_5_en_0 & _T_1125; // @[MemPrimitives.scala 125:64:@13480.4]
  assign StickySelects_7_io_ins_6 = io_rPort_6_en_0 & _T_1131; // @[MemPrimitives.scala 125:64:@13481.4]
  assign StickySelects_7_io_ins_7 = io_rPort_7_en_0 & _T_1137; // @[MemPrimitives.scala 125:64:@13482.4]
  assign StickySelects_7_io_ins_8 = io_rPort_8_en_0 & _T_1143; // @[MemPrimitives.scala 125:64:@13483.4]
  assign StickySelects_8_clock = clock; // @[:@13562.4]
  assign StickySelects_8_reset = reset; // @[:@13563.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1187; // @[MemPrimitives.scala 125:64:@13564.4]
  assign StickySelects_8_io_ins_1 = io_rPort_1_en_0 & _T_1193; // @[MemPrimitives.scala 125:64:@13565.4]
  assign StickySelects_8_io_ins_2 = io_rPort_2_en_0 & _T_1199; // @[MemPrimitives.scala 125:64:@13566.4]
  assign StickySelects_8_io_ins_3 = io_rPort_3_en_0 & _T_1205; // @[MemPrimitives.scala 125:64:@13567.4]
  assign StickySelects_8_io_ins_4 = io_rPort_4_en_0 & _T_1211; // @[MemPrimitives.scala 125:64:@13568.4]
  assign StickySelects_8_io_ins_5 = io_rPort_5_en_0 & _T_1217; // @[MemPrimitives.scala 125:64:@13569.4]
  assign StickySelects_8_io_ins_6 = io_rPort_6_en_0 & _T_1223; // @[MemPrimitives.scala 125:64:@13570.4]
  assign StickySelects_8_io_ins_7 = io_rPort_7_en_0 & _T_1229; // @[MemPrimitives.scala 125:64:@13571.4]
  assign StickySelects_8_io_ins_8 = io_rPort_8_en_0 & _T_1235; // @[MemPrimitives.scala 125:64:@13572.4]
  assign StickySelects_9_clock = clock; // @[:@13651.4]
  assign StickySelects_9_reset = reset; // @[:@13652.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_1279; // @[MemPrimitives.scala 125:64:@13653.4]
  assign StickySelects_9_io_ins_1 = io_rPort_1_en_0 & _T_1285; // @[MemPrimitives.scala 125:64:@13654.4]
  assign StickySelects_9_io_ins_2 = io_rPort_2_en_0 & _T_1291; // @[MemPrimitives.scala 125:64:@13655.4]
  assign StickySelects_9_io_ins_3 = io_rPort_3_en_0 & _T_1297; // @[MemPrimitives.scala 125:64:@13656.4]
  assign StickySelects_9_io_ins_4 = io_rPort_4_en_0 & _T_1303; // @[MemPrimitives.scala 125:64:@13657.4]
  assign StickySelects_9_io_ins_5 = io_rPort_5_en_0 & _T_1309; // @[MemPrimitives.scala 125:64:@13658.4]
  assign StickySelects_9_io_ins_6 = io_rPort_6_en_0 & _T_1315; // @[MemPrimitives.scala 125:64:@13659.4]
  assign StickySelects_9_io_ins_7 = io_rPort_7_en_0 & _T_1321; // @[MemPrimitives.scala 125:64:@13660.4]
  assign StickySelects_9_io_ins_8 = io_rPort_8_en_0 & _T_1327; // @[MemPrimitives.scala 125:64:@13661.4]
  assign StickySelects_10_clock = clock; // @[:@13740.4]
  assign StickySelects_10_reset = reset; // @[:@13741.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_1371; // @[MemPrimitives.scala 125:64:@13742.4]
  assign StickySelects_10_io_ins_1 = io_rPort_1_en_0 & _T_1377; // @[MemPrimitives.scala 125:64:@13743.4]
  assign StickySelects_10_io_ins_2 = io_rPort_2_en_0 & _T_1383; // @[MemPrimitives.scala 125:64:@13744.4]
  assign StickySelects_10_io_ins_3 = io_rPort_3_en_0 & _T_1389; // @[MemPrimitives.scala 125:64:@13745.4]
  assign StickySelects_10_io_ins_4 = io_rPort_4_en_0 & _T_1395; // @[MemPrimitives.scala 125:64:@13746.4]
  assign StickySelects_10_io_ins_5 = io_rPort_5_en_0 & _T_1401; // @[MemPrimitives.scala 125:64:@13747.4]
  assign StickySelects_10_io_ins_6 = io_rPort_6_en_0 & _T_1407; // @[MemPrimitives.scala 125:64:@13748.4]
  assign StickySelects_10_io_ins_7 = io_rPort_7_en_0 & _T_1413; // @[MemPrimitives.scala 125:64:@13749.4]
  assign StickySelects_10_io_ins_8 = io_rPort_8_en_0 & _T_1419; // @[MemPrimitives.scala 125:64:@13750.4]
  assign StickySelects_11_clock = clock; // @[:@13829.4]
  assign StickySelects_11_reset = reset; // @[:@13830.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_1463; // @[MemPrimitives.scala 125:64:@13831.4]
  assign StickySelects_11_io_ins_1 = io_rPort_1_en_0 & _T_1469; // @[MemPrimitives.scala 125:64:@13832.4]
  assign StickySelects_11_io_ins_2 = io_rPort_2_en_0 & _T_1475; // @[MemPrimitives.scala 125:64:@13833.4]
  assign StickySelects_11_io_ins_3 = io_rPort_3_en_0 & _T_1481; // @[MemPrimitives.scala 125:64:@13834.4]
  assign StickySelects_11_io_ins_4 = io_rPort_4_en_0 & _T_1487; // @[MemPrimitives.scala 125:64:@13835.4]
  assign StickySelects_11_io_ins_5 = io_rPort_5_en_0 & _T_1493; // @[MemPrimitives.scala 125:64:@13836.4]
  assign StickySelects_11_io_ins_6 = io_rPort_6_en_0 & _T_1499; // @[MemPrimitives.scala 125:64:@13837.4]
  assign StickySelects_11_io_ins_7 = io_rPort_7_en_0 & _T_1505; // @[MemPrimitives.scala 125:64:@13838.4]
  assign StickySelects_11_io_ins_8 = io_rPort_8_en_0 & _T_1511; // @[MemPrimitives.scala 125:64:@13839.4]
  assign RetimeWrapper_clock = clock; // @[:@13919.4]
  assign RetimeWrapper_reset = reset; // @[:@13920.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13922.4]
  assign RetimeWrapper_io_in = _T_451 & io_rPort_0_en_0; // @[package.scala 94:16:@13921.4]
  assign RetimeWrapper_1_clock = clock; // @[:@13927.4]
  assign RetimeWrapper_1_reset = reset; // @[:@13928.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13930.4]
  assign RetimeWrapper_1_io_in = _T_543 & io_rPort_0_en_0; // @[package.scala 94:16:@13929.4]
  assign RetimeWrapper_2_clock = clock; // @[:@13935.4]
  assign RetimeWrapper_2_reset = reset; // @[:@13936.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13938.4]
  assign RetimeWrapper_2_io_in = _T_635 & io_rPort_0_en_0; // @[package.scala 94:16:@13937.4]
  assign RetimeWrapper_3_clock = clock; // @[:@13943.4]
  assign RetimeWrapper_3_reset = reset; // @[:@13944.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13946.4]
  assign RetimeWrapper_3_io_in = _T_727 & io_rPort_0_en_0; // @[package.scala 94:16:@13945.4]
  assign RetimeWrapper_4_clock = clock; // @[:@13951.4]
  assign RetimeWrapper_4_reset = reset; // @[:@13952.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13954.4]
  assign RetimeWrapper_4_io_in = _T_819 & io_rPort_0_en_0; // @[package.scala 94:16:@13953.4]
  assign RetimeWrapper_5_clock = clock; // @[:@13959.4]
  assign RetimeWrapper_5_reset = reset; // @[:@13960.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13962.4]
  assign RetimeWrapper_5_io_in = _T_911 & io_rPort_0_en_0; // @[package.scala 94:16:@13961.4]
  assign RetimeWrapper_6_clock = clock; // @[:@13967.4]
  assign RetimeWrapper_6_reset = reset; // @[:@13968.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13970.4]
  assign RetimeWrapper_6_io_in = _T_1003 & io_rPort_0_en_0; // @[package.scala 94:16:@13969.4]
  assign RetimeWrapper_7_clock = clock; // @[:@13975.4]
  assign RetimeWrapper_7_reset = reset; // @[:@13976.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13978.4]
  assign RetimeWrapper_7_io_in = _T_1095 & io_rPort_0_en_0; // @[package.scala 94:16:@13977.4]
  assign RetimeWrapper_8_clock = clock; // @[:@13983.4]
  assign RetimeWrapper_8_reset = reset; // @[:@13984.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13986.4]
  assign RetimeWrapper_8_io_in = _T_1187 & io_rPort_0_en_0; // @[package.scala 94:16:@13985.4]
  assign RetimeWrapper_9_clock = clock; // @[:@13991.4]
  assign RetimeWrapper_9_reset = reset; // @[:@13992.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13994.4]
  assign RetimeWrapper_9_io_in = _T_1279 & io_rPort_0_en_0; // @[package.scala 94:16:@13993.4]
  assign RetimeWrapper_10_clock = clock; // @[:@13999.4]
  assign RetimeWrapper_10_reset = reset; // @[:@14000.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14002.4]
  assign RetimeWrapper_10_io_in = _T_1371 & io_rPort_0_en_0; // @[package.scala 94:16:@14001.4]
  assign RetimeWrapper_11_clock = clock; // @[:@14007.4]
  assign RetimeWrapper_11_reset = reset; // @[:@14008.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14010.4]
  assign RetimeWrapper_11_io_in = _T_1463 & io_rPort_0_en_0; // @[package.scala 94:16:@14009.4]
  assign RetimeWrapper_12_clock = clock; // @[:@14063.4]
  assign RetimeWrapper_12_reset = reset; // @[:@14064.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14066.4]
  assign RetimeWrapper_12_io_in = _T_457 & io_rPort_1_en_0; // @[package.scala 94:16:@14065.4]
  assign RetimeWrapper_13_clock = clock; // @[:@14071.4]
  assign RetimeWrapper_13_reset = reset; // @[:@14072.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14074.4]
  assign RetimeWrapper_13_io_in = _T_549 & io_rPort_1_en_0; // @[package.scala 94:16:@14073.4]
  assign RetimeWrapper_14_clock = clock; // @[:@14079.4]
  assign RetimeWrapper_14_reset = reset; // @[:@14080.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14082.4]
  assign RetimeWrapper_14_io_in = _T_641 & io_rPort_1_en_0; // @[package.scala 94:16:@14081.4]
  assign RetimeWrapper_15_clock = clock; // @[:@14087.4]
  assign RetimeWrapper_15_reset = reset; // @[:@14088.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14090.4]
  assign RetimeWrapper_15_io_in = _T_733 & io_rPort_1_en_0; // @[package.scala 94:16:@14089.4]
  assign RetimeWrapper_16_clock = clock; // @[:@14095.4]
  assign RetimeWrapper_16_reset = reset; // @[:@14096.4]
  assign RetimeWrapper_16_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14098.4]
  assign RetimeWrapper_16_io_in = _T_825 & io_rPort_1_en_0; // @[package.scala 94:16:@14097.4]
  assign RetimeWrapper_17_clock = clock; // @[:@14103.4]
  assign RetimeWrapper_17_reset = reset; // @[:@14104.4]
  assign RetimeWrapper_17_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14106.4]
  assign RetimeWrapper_17_io_in = _T_917 & io_rPort_1_en_0; // @[package.scala 94:16:@14105.4]
  assign RetimeWrapper_18_clock = clock; // @[:@14111.4]
  assign RetimeWrapper_18_reset = reset; // @[:@14112.4]
  assign RetimeWrapper_18_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14114.4]
  assign RetimeWrapper_18_io_in = _T_1009 & io_rPort_1_en_0; // @[package.scala 94:16:@14113.4]
  assign RetimeWrapper_19_clock = clock; // @[:@14119.4]
  assign RetimeWrapper_19_reset = reset; // @[:@14120.4]
  assign RetimeWrapper_19_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14122.4]
  assign RetimeWrapper_19_io_in = _T_1101 & io_rPort_1_en_0; // @[package.scala 94:16:@14121.4]
  assign RetimeWrapper_20_clock = clock; // @[:@14127.4]
  assign RetimeWrapper_20_reset = reset; // @[:@14128.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14130.4]
  assign RetimeWrapper_20_io_in = _T_1193 & io_rPort_1_en_0; // @[package.scala 94:16:@14129.4]
  assign RetimeWrapper_21_clock = clock; // @[:@14135.4]
  assign RetimeWrapper_21_reset = reset; // @[:@14136.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14138.4]
  assign RetimeWrapper_21_io_in = _T_1285 & io_rPort_1_en_0; // @[package.scala 94:16:@14137.4]
  assign RetimeWrapper_22_clock = clock; // @[:@14143.4]
  assign RetimeWrapper_22_reset = reset; // @[:@14144.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14146.4]
  assign RetimeWrapper_22_io_in = _T_1377 & io_rPort_1_en_0; // @[package.scala 94:16:@14145.4]
  assign RetimeWrapper_23_clock = clock; // @[:@14151.4]
  assign RetimeWrapper_23_reset = reset; // @[:@14152.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14154.4]
  assign RetimeWrapper_23_io_in = _T_1469 & io_rPort_1_en_0; // @[package.scala 94:16:@14153.4]
  assign RetimeWrapper_24_clock = clock; // @[:@14207.4]
  assign RetimeWrapper_24_reset = reset; // @[:@14208.4]
  assign RetimeWrapper_24_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14210.4]
  assign RetimeWrapper_24_io_in = _T_463 & io_rPort_2_en_0; // @[package.scala 94:16:@14209.4]
  assign RetimeWrapper_25_clock = clock; // @[:@14215.4]
  assign RetimeWrapper_25_reset = reset; // @[:@14216.4]
  assign RetimeWrapper_25_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14218.4]
  assign RetimeWrapper_25_io_in = _T_555 & io_rPort_2_en_0; // @[package.scala 94:16:@14217.4]
  assign RetimeWrapper_26_clock = clock; // @[:@14223.4]
  assign RetimeWrapper_26_reset = reset; // @[:@14224.4]
  assign RetimeWrapper_26_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14226.4]
  assign RetimeWrapper_26_io_in = _T_647 & io_rPort_2_en_0; // @[package.scala 94:16:@14225.4]
  assign RetimeWrapper_27_clock = clock; // @[:@14231.4]
  assign RetimeWrapper_27_reset = reset; // @[:@14232.4]
  assign RetimeWrapper_27_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14234.4]
  assign RetimeWrapper_27_io_in = _T_739 & io_rPort_2_en_0; // @[package.scala 94:16:@14233.4]
  assign RetimeWrapper_28_clock = clock; // @[:@14239.4]
  assign RetimeWrapper_28_reset = reset; // @[:@14240.4]
  assign RetimeWrapper_28_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14242.4]
  assign RetimeWrapper_28_io_in = _T_831 & io_rPort_2_en_0; // @[package.scala 94:16:@14241.4]
  assign RetimeWrapper_29_clock = clock; // @[:@14247.4]
  assign RetimeWrapper_29_reset = reset; // @[:@14248.4]
  assign RetimeWrapper_29_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14250.4]
  assign RetimeWrapper_29_io_in = _T_923 & io_rPort_2_en_0; // @[package.scala 94:16:@14249.4]
  assign RetimeWrapper_30_clock = clock; // @[:@14255.4]
  assign RetimeWrapper_30_reset = reset; // @[:@14256.4]
  assign RetimeWrapper_30_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14258.4]
  assign RetimeWrapper_30_io_in = _T_1015 & io_rPort_2_en_0; // @[package.scala 94:16:@14257.4]
  assign RetimeWrapper_31_clock = clock; // @[:@14263.4]
  assign RetimeWrapper_31_reset = reset; // @[:@14264.4]
  assign RetimeWrapper_31_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14266.4]
  assign RetimeWrapper_31_io_in = _T_1107 & io_rPort_2_en_0; // @[package.scala 94:16:@14265.4]
  assign RetimeWrapper_32_clock = clock; // @[:@14271.4]
  assign RetimeWrapper_32_reset = reset; // @[:@14272.4]
  assign RetimeWrapper_32_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14274.4]
  assign RetimeWrapper_32_io_in = _T_1199 & io_rPort_2_en_0; // @[package.scala 94:16:@14273.4]
  assign RetimeWrapper_33_clock = clock; // @[:@14279.4]
  assign RetimeWrapper_33_reset = reset; // @[:@14280.4]
  assign RetimeWrapper_33_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14282.4]
  assign RetimeWrapper_33_io_in = _T_1291 & io_rPort_2_en_0; // @[package.scala 94:16:@14281.4]
  assign RetimeWrapper_34_clock = clock; // @[:@14287.4]
  assign RetimeWrapper_34_reset = reset; // @[:@14288.4]
  assign RetimeWrapper_34_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14290.4]
  assign RetimeWrapper_34_io_in = _T_1383 & io_rPort_2_en_0; // @[package.scala 94:16:@14289.4]
  assign RetimeWrapper_35_clock = clock; // @[:@14295.4]
  assign RetimeWrapper_35_reset = reset; // @[:@14296.4]
  assign RetimeWrapper_35_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14298.4]
  assign RetimeWrapper_35_io_in = _T_1475 & io_rPort_2_en_0; // @[package.scala 94:16:@14297.4]
  assign RetimeWrapper_36_clock = clock; // @[:@14351.4]
  assign RetimeWrapper_36_reset = reset; // @[:@14352.4]
  assign RetimeWrapper_36_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14354.4]
  assign RetimeWrapper_36_io_in = _T_469 & io_rPort_3_en_0; // @[package.scala 94:16:@14353.4]
  assign RetimeWrapper_37_clock = clock; // @[:@14359.4]
  assign RetimeWrapper_37_reset = reset; // @[:@14360.4]
  assign RetimeWrapper_37_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14362.4]
  assign RetimeWrapper_37_io_in = _T_561 & io_rPort_3_en_0; // @[package.scala 94:16:@14361.4]
  assign RetimeWrapper_38_clock = clock; // @[:@14367.4]
  assign RetimeWrapper_38_reset = reset; // @[:@14368.4]
  assign RetimeWrapper_38_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14370.4]
  assign RetimeWrapper_38_io_in = _T_653 & io_rPort_3_en_0; // @[package.scala 94:16:@14369.4]
  assign RetimeWrapper_39_clock = clock; // @[:@14375.4]
  assign RetimeWrapper_39_reset = reset; // @[:@14376.4]
  assign RetimeWrapper_39_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14378.4]
  assign RetimeWrapper_39_io_in = _T_745 & io_rPort_3_en_0; // @[package.scala 94:16:@14377.4]
  assign RetimeWrapper_40_clock = clock; // @[:@14383.4]
  assign RetimeWrapper_40_reset = reset; // @[:@14384.4]
  assign RetimeWrapper_40_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14386.4]
  assign RetimeWrapper_40_io_in = _T_837 & io_rPort_3_en_0; // @[package.scala 94:16:@14385.4]
  assign RetimeWrapper_41_clock = clock; // @[:@14391.4]
  assign RetimeWrapper_41_reset = reset; // @[:@14392.4]
  assign RetimeWrapper_41_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14394.4]
  assign RetimeWrapper_41_io_in = _T_929 & io_rPort_3_en_0; // @[package.scala 94:16:@14393.4]
  assign RetimeWrapper_42_clock = clock; // @[:@14399.4]
  assign RetimeWrapper_42_reset = reset; // @[:@14400.4]
  assign RetimeWrapper_42_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14402.4]
  assign RetimeWrapper_42_io_in = _T_1021 & io_rPort_3_en_0; // @[package.scala 94:16:@14401.4]
  assign RetimeWrapper_43_clock = clock; // @[:@14407.4]
  assign RetimeWrapper_43_reset = reset; // @[:@14408.4]
  assign RetimeWrapper_43_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14410.4]
  assign RetimeWrapper_43_io_in = _T_1113 & io_rPort_3_en_0; // @[package.scala 94:16:@14409.4]
  assign RetimeWrapper_44_clock = clock; // @[:@14415.4]
  assign RetimeWrapper_44_reset = reset; // @[:@14416.4]
  assign RetimeWrapper_44_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14418.4]
  assign RetimeWrapper_44_io_in = _T_1205 & io_rPort_3_en_0; // @[package.scala 94:16:@14417.4]
  assign RetimeWrapper_45_clock = clock; // @[:@14423.4]
  assign RetimeWrapper_45_reset = reset; // @[:@14424.4]
  assign RetimeWrapper_45_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14426.4]
  assign RetimeWrapper_45_io_in = _T_1297 & io_rPort_3_en_0; // @[package.scala 94:16:@14425.4]
  assign RetimeWrapper_46_clock = clock; // @[:@14431.4]
  assign RetimeWrapper_46_reset = reset; // @[:@14432.4]
  assign RetimeWrapper_46_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14434.4]
  assign RetimeWrapper_46_io_in = _T_1389 & io_rPort_3_en_0; // @[package.scala 94:16:@14433.4]
  assign RetimeWrapper_47_clock = clock; // @[:@14439.4]
  assign RetimeWrapper_47_reset = reset; // @[:@14440.4]
  assign RetimeWrapper_47_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14442.4]
  assign RetimeWrapper_47_io_in = _T_1481 & io_rPort_3_en_0; // @[package.scala 94:16:@14441.4]
  assign RetimeWrapper_48_clock = clock; // @[:@14495.4]
  assign RetimeWrapper_48_reset = reset; // @[:@14496.4]
  assign RetimeWrapper_48_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14498.4]
  assign RetimeWrapper_48_io_in = _T_475 & io_rPort_4_en_0; // @[package.scala 94:16:@14497.4]
  assign RetimeWrapper_49_clock = clock; // @[:@14503.4]
  assign RetimeWrapper_49_reset = reset; // @[:@14504.4]
  assign RetimeWrapper_49_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14506.4]
  assign RetimeWrapper_49_io_in = _T_567 & io_rPort_4_en_0; // @[package.scala 94:16:@14505.4]
  assign RetimeWrapper_50_clock = clock; // @[:@14511.4]
  assign RetimeWrapper_50_reset = reset; // @[:@14512.4]
  assign RetimeWrapper_50_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14514.4]
  assign RetimeWrapper_50_io_in = _T_659 & io_rPort_4_en_0; // @[package.scala 94:16:@14513.4]
  assign RetimeWrapper_51_clock = clock; // @[:@14519.4]
  assign RetimeWrapper_51_reset = reset; // @[:@14520.4]
  assign RetimeWrapper_51_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14522.4]
  assign RetimeWrapper_51_io_in = _T_751 & io_rPort_4_en_0; // @[package.scala 94:16:@14521.4]
  assign RetimeWrapper_52_clock = clock; // @[:@14527.4]
  assign RetimeWrapper_52_reset = reset; // @[:@14528.4]
  assign RetimeWrapper_52_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14530.4]
  assign RetimeWrapper_52_io_in = _T_843 & io_rPort_4_en_0; // @[package.scala 94:16:@14529.4]
  assign RetimeWrapper_53_clock = clock; // @[:@14535.4]
  assign RetimeWrapper_53_reset = reset; // @[:@14536.4]
  assign RetimeWrapper_53_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14538.4]
  assign RetimeWrapper_53_io_in = _T_935 & io_rPort_4_en_0; // @[package.scala 94:16:@14537.4]
  assign RetimeWrapper_54_clock = clock; // @[:@14543.4]
  assign RetimeWrapper_54_reset = reset; // @[:@14544.4]
  assign RetimeWrapper_54_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14546.4]
  assign RetimeWrapper_54_io_in = _T_1027 & io_rPort_4_en_0; // @[package.scala 94:16:@14545.4]
  assign RetimeWrapper_55_clock = clock; // @[:@14551.4]
  assign RetimeWrapper_55_reset = reset; // @[:@14552.4]
  assign RetimeWrapper_55_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14554.4]
  assign RetimeWrapper_55_io_in = _T_1119 & io_rPort_4_en_0; // @[package.scala 94:16:@14553.4]
  assign RetimeWrapper_56_clock = clock; // @[:@14559.4]
  assign RetimeWrapper_56_reset = reset; // @[:@14560.4]
  assign RetimeWrapper_56_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14562.4]
  assign RetimeWrapper_56_io_in = _T_1211 & io_rPort_4_en_0; // @[package.scala 94:16:@14561.4]
  assign RetimeWrapper_57_clock = clock; // @[:@14567.4]
  assign RetimeWrapper_57_reset = reset; // @[:@14568.4]
  assign RetimeWrapper_57_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14570.4]
  assign RetimeWrapper_57_io_in = _T_1303 & io_rPort_4_en_0; // @[package.scala 94:16:@14569.4]
  assign RetimeWrapper_58_clock = clock; // @[:@14575.4]
  assign RetimeWrapper_58_reset = reset; // @[:@14576.4]
  assign RetimeWrapper_58_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14578.4]
  assign RetimeWrapper_58_io_in = _T_1395 & io_rPort_4_en_0; // @[package.scala 94:16:@14577.4]
  assign RetimeWrapper_59_clock = clock; // @[:@14583.4]
  assign RetimeWrapper_59_reset = reset; // @[:@14584.4]
  assign RetimeWrapper_59_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14586.4]
  assign RetimeWrapper_59_io_in = _T_1487 & io_rPort_4_en_0; // @[package.scala 94:16:@14585.4]
  assign RetimeWrapper_60_clock = clock; // @[:@14639.4]
  assign RetimeWrapper_60_reset = reset; // @[:@14640.4]
  assign RetimeWrapper_60_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14642.4]
  assign RetimeWrapper_60_io_in = _T_481 & io_rPort_5_en_0; // @[package.scala 94:16:@14641.4]
  assign RetimeWrapper_61_clock = clock; // @[:@14647.4]
  assign RetimeWrapper_61_reset = reset; // @[:@14648.4]
  assign RetimeWrapper_61_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14650.4]
  assign RetimeWrapper_61_io_in = _T_573 & io_rPort_5_en_0; // @[package.scala 94:16:@14649.4]
  assign RetimeWrapper_62_clock = clock; // @[:@14655.4]
  assign RetimeWrapper_62_reset = reset; // @[:@14656.4]
  assign RetimeWrapper_62_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14658.4]
  assign RetimeWrapper_62_io_in = _T_665 & io_rPort_5_en_0; // @[package.scala 94:16:@14657.4]
  assign RetimeWrapper_63_clock = clock; // @[:@14663.4]
  assign RetimeWrapper_63_reset = reset; // @[:@14664.4]
  assign RetimeWrapper_63_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14666.4]
  assign RetimeWrapper_63_io_in = _T_757 & io_rPort_5_en_0; // @[package.scala 94:16:@14665.4]
  assign RetimeWrapper_64_clock = clock; // @[:@14671.4]
  assign RetimeWrapper_64_reset = reset; // @[:@14672.4]
  assign RetimeWrapper_64_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14674.4]
  assign RetimeWrapper_64_io_in = _T_849 & io_rPort_5_en_0; // @[package.scala 94:16:@14673.4]
  assign RetimeWrapper_65_clock = clock; // @[:@14679.4]
  assign RetimeWrapper_65_reset = reset; // @[:@14680.4]
  assign RetimeWrapper_65_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14682.4]
  assign RetimeWrapper_65_io_in = _T_941 & io_rPort_5_en_0; // @[package.scala 94:16:@14681.4]
  assign RetimeWrapper_66_clock = clock; // @[:@14687.4]
  assign RetimeWrapper_66_reset = reset; // @[:@14688.4]
  assign RetimeWrapper_66_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14690.4]
  assign RetimeWrapper_66_io_in = _T_1033 & io_rPort_5_en_0; // @[package.scala 94:16:@14689.4]
  assign RetimeWrapper_67_clock = clock; // @[:@14695.4]
  assign RetimeWrapper_67_reset = reset; // @[:@14696.4]
  assign RetimeWrapper_67_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14698.4]
  assign RetimeWrapper_67_io_in = _T_1125 & io_rPort_5_en_0; // @[package.scala 94:16:@14697.4]
  assign RetimeWrapper_68_clock = clock; // @[:@14703.4]
  assign RetimeWrapper_68_reset = reset; // @[:@14704.4]
  assign RetimeWrapper_68_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14706.4]
  assign RetimeWrapper_68_io_in = _T_1217 & io_rPort_5_en_0; // @[package.scala 94:16:@14705.4]
  assign RetimeWrapper_69_clock = clock; // @[:@14711.4]
  assign RetimeWrapper_69_reset = reset; // @[:@14712.4]
  assign RetimeWrapper_69_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14714.4]
  assign RetimeWrapper_69_io_in = _T_1309 & io_rPort_5_en_0; // @[package.scala 94:16:@14713.4]
  assign RetimeWrapper_70_clock = clock; // @[:@14719.4]
  assign RetimeWrapper_70_reset = reset; // @[:@14720.4]
  assign RetimeWrapper_70_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14722.4]
  assign RetimeWrapper_70_io_in = _T_1401 & io_rPort_5_en_0; // @[package.scala 94:16:@14721.4]
  assign RetimeWrapper_71_clock = clock; // @[:@14727.4]
  assign RetimeWrapper_71_reset = reset; // @[:@14728.4]
  assign RetimeWrapper_71_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14730.4]
  assign RetimeWrapper_71_io_in = _T_1493 & io_rPort_5_en_0; // @[package.scala 94:16:@14729.4]
  assign RetimeWrapper_72_clock = clock; // @[:@14783.4]
  assign RetimeWrapper_72_reset = reset; // @[:@14784.4]
  assign RetimeWrapper_72_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14786.4]
  assign RetimeWrapper_72_io_in = _T_487 & io_rPort_6_en_0; // @[package.scala 94:16:@14785.4]
  assign RetimeWrapper_73_clock = clock; // @[:@14791.4]
  assign RetimeWrapper_73_reset = reset; // @[:@14792.4]
  assign RetimeWrapper_73_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14794.4]
  assign RetimeWrapper_73_io_in = _T_579 & io_rPort_6_en_0; // @[package.scala 94:16:@14793.4]
  assign RetimeWrapper_74_clock = clock; // @[:@14799.4]
  assign RetimeWrapper_74_reset = reset; // @[:@14800.4]
  assign RetimeWrapper_74_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14802.4]
  assign RetimeWrapper_74_io_in = _T_671 & io_rPort_6_en_0; // @[package.scala 94:16:@14801.4]
  assign RetimeWrapper_75_clock = clock; // @[:@14807.4]
  assign RetimeWrapper_75_reset = reset; // @[:@14808.4]
  assign RetimeWrapper_75_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14810.4]
  assign RetimeWrapper_75_io_in = _T_763 & io_rPort_6_en_0; // @[package.scala 94:16:@14809.4]
  assign RetimeWrapper_76_clock = clock; // @[:@14815.4]
  assign RetimeWrapper_76_reset = reset; // @[:@14816.4]
  assign RetimeWrapper_76_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14818.4]
  assign RetimeWrapper_76_io_in = _T_855 & io_rPort_6_en_0; // @[package.scala 94:16:@14817.4]
  assign RetimeWrapper_77_clock = clock; // @[:@14823.4]
  assign RetimeWrapper_77_reset = reset; // @[:@14824.4]
  assign RetimeWrapper_77_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14826.4]
  assign RetimeWrapper_77_io_in = _T_947 & io_rPort_6_en_0; // @[package.scala 94:16:@14825.4]
  assign RetimeWrapper_78_clock = clock; // @[:@14831.4]
  assign RetimeWrapper_78_reset = reset; // @[:@14832.4]
  assign RetimeWrapper_78_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14834.4]
  assign RetimeWrapper_78_io_in = _T_1039 & io_rPort_6_en_0; // @[package.scala 94:16:@14833.4]
  assign RetimeWrapper_79_clock = clock; // @[:@14839.4]
  assign RetimeWrapper_79_reset = reset; // @[:@14840.4]
  assign RetimeWrapper_79_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14842.4]
  assign RetimeWrapper_79_io_in = _T_1131 & io_rPort_6_en_0; // @[package.scala 94:16:@14841.4]
  assign RetimeWrapper_80_clock = clock; // @[:@14847.4]
  assign RetimeWrapper_80_reset = reset; // @[:@14848.4]
  assign RetimeWrapper_80_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14850.4]
  assign RetimeWrapper_80_io_in = _T_1223 & io_rPort_6_en_0; // @[package.scala 94:16:@14849.4]
  assign RetimeWrapper_81_clock = clock; // @[:@14855.4]
  assign RetimeWrapper_81_reset = reset; // @[:@14856.4]
  assign RetimeWrapper_81_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14858.4]
  assign RetimeWrapper_81_io_in = _T_1315 & io_rPort_6_en_0; // @[package.scala 94:16:@14857.4]
  assign RetimeWrapper_82_clock = clock; // @[:@14863.4]
  assign RetimeWrapper_82_reset = reset; // @[:@14864.4]
  assign RetimeWrapper_82_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14866.4]
  assign RetimeWrapper_82_io_in = _T_1407 & io_rPort_6_en_0; // @[package.scala 94:16:@14865.4]
  assign RetimeWrapper_83_clock = clock; // @[:@14871.4]
  assign RetimeWrapper_83_reset = reset; // @[:@14872.4]
  assign RetimeWrapper_83_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14874.4]
  assign RetimeWrapper_83_io_in = _T_1499 & io_rPort_6_en_0; // @[package.scala 94:16:@14873.4]
  assign RetimeWrapper_84_clock = clock; // @[:@14927.4]
  assign RetimeWrapper_84_reset = reset; // @[:@14928.4]
  assign RetimeWrapper_84_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14930.4]
  assign RetimeWrapper_84_io_in = _T_493 & io_rPort_7_en_0; // @[package.scala 94:16:@14929.4]
  assign RetimeWrapper_85_clock = clock; // @[:@14935.4]
  assign RetimeWrapper_85_reset = reset; // @[:@14936.4]
  assign RetimeWrapper_85_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14938.4]
  assign RetimeWrapper_85_io_in = _T_585 & io_rPort_7_en_0; // @[package.scala 94:16:@14937.4]
  assign RetimeWrapper_86_clock = clock; // @[:@14943.4]
  assign RetimeWrapper_86_reset = reset; // @[:@14944.4]
  assign RetimeWrapper_86_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14946.4]
  assign RetimeWrapper_86_io_in = _T_677 & io_rPort_7_en_0; // @[package.scala 94:16:@14945.4]
  assign RetimeWrapper_87_clock = clock; // @[:@14951.4]
  assign RetimeWrapper_87_reset = reset; // @[:@14952.4]
  assign RetimeWrapper_87_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14954.4]
  assign RetimeWrapper_87_io_in = _T_769 & io_rPort_7_en_0; // @[package.scala 94:16:@14953.4]
  assign RetimeWrapper_88_clock = clock; // @[:@14959.4]
  assign RetimeWrapper_88_reset = reset; // @[:@14960.4]
  assign RetimeWrapper_88_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14962.4]
  assign RetimeWrapper_88_io_in = _T_861 & io_rPort_7_en_0; // @[package.scala 94:16:@14961.4]
  assign RetimeWrapper_89_clock = clock; // @[:@14967.4]
  assign RetimeWrapper_89_reset = reset; // @[:@14968.4]
  assign RetimeWrapper_89_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14970.4]
  assign RetimeWrapper_89_io_in = _T_953 & io_rPort_7_en_0; // @[package.scala 94:16:@14969.4]
  assign RetimeWrapper_90_clock = clock; // @[:@14975.4]
  assign RetimeWrapper_90_reset = reset; // @[:@14976.4]
  assign RetimeWrapper_90_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14978.4]
  assign RetimeWrapper_90_io_in = _T_1045 & io_rPort_7_en_0; // @[package.scala 94:16:@14977.4]
  assign RetimeWrapper_91_clock = clock; // @[:@14983.4]
  assign RetimeWrapper_91_reset = reset; // @[:@14984.4]
  assign RetimeWrapper_91_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14986.4]
  assign RetimeWrapper_91_io_in = _T_1137 & io_rPort_7_en_0; // @[package.scala 94:16:@14985.4]
  assign RetimeWrapper_92_clock = clock; // @[:@14991.4]
  assign RetimeWrapper_92_reset = reset; // @[:@14992.4]
  assign RetimeWrapper_92_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14994.4]
  assign RetimeWrapper_92_io_in = _T_1229 & io_rPort_7_en_0; // @[package.scala 94:16:@14993.4]
  assign RetimeWrapper_93_clock = clock; // @[:@14999.4]
  assign RetimeWrapper_93_reset = reset; // @[:@15000.4]
  assign RetimeWrapper_93_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15002.4]
  assign RetimeWrapper_93_io_in = _T_1321 & io_rPort_7_en_0; // @[package.scala 94:16:@15001.4]
  assign RetimeWrapper_94_clock = clock; // @[:@15007.4]
  assign RetimeWrapper_94_reset = reset; // @[:@15008.4]
  assign RetimeWrapper_94_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15010.4]
  assign RetimeWrapper_94_io_in = _T_1413 & io_rPort_7_en_0; // @[package.scala 94:16:@15009.4]
  assign RetimeWrapper_95_clock = clock; // @[:@15015.4]
  assign RetimeWrapper_95_reset = reset; // @[:@15016.4]
  assign RetimeWrapper_95_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15018.4]
  assign RetimeWrapper_95_io_in = _T_1505 & io_rPort_7_en_0; // @[package.scala 94:16:@15017.4]
  assign RetimeWrapper_96_clock = clock; // @[:@15071.4]
  assign RetimeWrapper_96_reset = reset; // @[:@15072.4]
  assign RetimeWrapper_96_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15074.4]
  assign RetimeWrapper_96_io_in = _T_499 & io_rPort_8_en_0; // @[package.scala 94:16:@15073.4]
  assign RetimeWrapper_97_clock = clock; // @[:@15079.4]
  assign RetimeWrapper_97_reset = reset; // @[:@15080.4]
  assign RetimeWrapper_97_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15082.4]
  assign RetimeWrapper_97_io_in = _T_591 & io_rPort_8_en_0; // @[package.scala 94:16:@15081.4]
  assign RetimeWrapper_98_clock = clock; // @[:@15087.4]
  assign RetimeWrapper_98_reset = reset; // @[:@15088.4]
  assign RetimeWrapper_98_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15090.4]
  assign RetimeWrapper_98_io_in = _T_683 & io_rPort_8_en_0; // @[package.scala 94:16:@15089.4]
  assign RetimeWrapper_99_clock = clock; // @[:@15095.4]
  assign RetimeWrapper_99_reset = reset; // @[:@15096.4]
  assign RetimeWrapper_99_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15098.4]
  assign RetimeWrapper_99_io_in = _T_775 & io_rPort_8_en_0; // @[package.scala 94:16:@15097.4]
  assign RetimeWrapper_100_clock = clock; // @[:@15103.4]
  assign RetimeWrapper_100_reset = reset; // @[:@15104.4]
  assign RetimeWrapper_100_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15106.4]
  assign RetimeWrapper_100_io_in = _T_867 & io_rPort_8_en_0; // @[package.scala 94:16:@15105.4]
  assign RetimeWrapper_101_clock = clock; // @[:@15111.4]
  assign RetimeWrapper_101_reset = reset; // @[:@15112.4]
  assign RetimeWrapper_101_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15114.4]
  assign RetimeWrapper_101_io_in = _T_959 & io_rPort_8_en_0; // @[package.scala 94:16:@15113.4]
  assign RetimeWrapper_102_clock = clock; // @[:@15119.4]
  assign RetimeWrapper_102_reset = reset; // @[:@15120.4]
  assign RetimeWrapper_102_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15122.4]
  assign RetimeWrapper_102_io_in = _T_1051 & io_rPort_8_en_0; // @[package.scala 94:16:@15121.4]
  assign RetimeWrapper_103_clock = clock; // @[:@15127.4]
  assign RetimeWrapper_103_reset = reset; // @[:@15128.4]
  assign RetimeWrapper_103_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15130.4]
  assign RetimeWrapper_103_io_in = _T_1143 & io_rPort_8_en_0; // @[package.scala 94:16:@15129.4]
  assign RetimeWrapper_104_clock = clock; // @[:@15135.4]
  assign RetimeWrapper_104_reset = reset; // @[:@15136.4]
  assign RetimeWrapper_104_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15138.4]
  assign RetimeWrapper_104_io_in = _T_1235 & io_rPort_8_en_0; // @[package.scala 94:16:@15137.4]
  assign RetimeWrapper_105_clock = clock; // @[:@15143.4]
  assign RetimeWrapper_105_reset = reset; // @[:@15144.4]
  assign RetimeWrapper_105_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15146.4]
  assign RetimeWrapper_105_io_in = _T_1327 & io_rPort_8_en_0; // @[package.scala 94:16:@15145.4]
  assign RetimeWrapper_106_clock = clock; // @[:@15151.4]
  assign RetimeWrapper_106_reset = reset; // @[:@15152.4]
  assign RetimeWrapper_106_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15154.4]
  assign RetimeWrapper_106_io_in = _T_1419 & io_rPort_8_en_0; // @[package.scala 94:16:@15153.4]
  assign RetimeWrapper_107_clock = clock; // @[:@15159.4]
  assign RetimeWrapper_107_reset = reset; // @[:@15160.4]
  assign RetimeWrapper_107_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15162.4]
  assign RetimeWrapper_107_io_in = _T_1511 & io_rPort_8_en_0; // @[package.scala 94:16:@15161.4]
endmodule
module StickySelects_13( // @[:@16462.2]
  input   clock, // @[:@16463.4]
  input   reset, // @[:@16464.4]
  input   io_ins_0, // @[:@16465.4]
  input   io_ins_1, // @[:@16465.4]
  input   io_ins_2, // @[:@16465.4]
  input   io_ins_3, // @[:@16465.4]
  output  io_outs_0, // @[:@16465.4]
  output  io_outs_1, // @[:@16465.4]
  output  io_outs_2, // @[:@16465.4]
  output  io_outs_3 // @[:@16465.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@16467.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@16468.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@16469.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@16470.4]
  reg [31:0] _RAND_3;
  wire  _T_29; // @[StickySelects.scala 47:46:@16471.4]
  wire  _T_30; // @[StickySelects.scala 47:46:@16472.4]
  wire  _T_31; // @[StickySelects.scala 49:53:@16473.4]
  wire  _T_32; // @[StickySelects.scala 49:21:@16474.4]
  wire  _T_33; // @[StickySelects.scala 47:46:@16476.4]
  wire  _T_34; // @[StickySelects.scala 47:46:@16477.4]
  wire  _T_35; // @[StickySelects.scala 49:53:@16478.4]
  wire  _T_36; // @[StickySelects.scala 49:21:@16479.4]
  wire  _T_37; // @[StickySelects.scala 47:46:@16481.4]
  wire  _T_38; // @[StickySelects.scala 47:46:@16482.4]
  wire  _T_39; // @[StickySelects.scala 49:53:@16483.4]
  wire  _T_40; // @[StickySelects.scala 49:21:@16484.4]
  wire  _T_42; // @[StickySelects.scala 47:46:@16487.4]
  wire  _T_43; // @[StickySelects.scala 49:53:@16488.4]
  wire  _T_44; // @[StickySelects.scala 49:21:@16489.4]
  assign _T_29 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@16471.4]
  assign _T_30 = _T_29 | io_ins_3; // @[StickySelects.scala 47:46:@16472.4]
  assign _T_31 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@16473.4]
  assign _T_32 = _T_30 ? io_ins_0 : _T_31; // @[StickySelects.scala 49:21:@16474.4]
  assign _T_33 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@16476.4]
  assign _T_34 = _T_33 | io_ins_3; // @[StickySelects.scala 47:46:@16477.4]
  assign _T_35 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@16478.4]
  assign _T_36 = _T_34 ? io_ins_1 : _T_35; // @[StickySelects.scala 49:21:@16479.4]
  assign _T_37 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@16481.4]
  assign _T_38 = _T_37 | io_ins_3; // @[StickySelects.scala 47:46:@16482.4]
  assign _T_39 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@16483.4]
  assign _T_40 = _T_38 ? io_ins_2 : _T_39; // @[StickySelects.scala 49:21:@16484.4]
  assign _T_42 = _T_37 | io_ins_2; // @[StickySelects.scala 47:46:@16487.4]
  assign _T_43 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@16488.4]
  assign _T_44 = _T_42 ? io_ins_3 : _T_43; // @[StickySelects.scala 49:21:@16489.4]
  assign io_outs_0 = _T_30 ? io_ins_0 : _T_31; // @[StickySelects.scala 53:57:@16491.4]
  assign io_outs_1 = _T_34 ? io_ins_1 : _T_35; // @[StickySelects.scala 53:57:@16492.4]
  assign io_outs_2 = _T_38 ? io_ins_2 : _T_39; // @[StickySelects.scala 53:57:@16493.4]
  assign io_outs_3 = _T_42 ? io_ins_3 : _T_43; // @[StickySelects.scala 53:57:@16494.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_30) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_31;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_34) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_35;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_38) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_39;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_42) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_43;
      end
    end
  end
endmodule
module x242_lb2_0( // @[:@18406.2]
  input         clock, // @[:@18407.4]
  input         reset, // @[:@18408.4]
  input  [1:0]  io_rPort_3_banks_1, // @[:@18409.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@18409.4]
  input  [9:0]  io_rPort_3_ofs_0, // @[:@18409.4]
  input         io_rPort_3_en_0, // @[:@18409.4]
  input         io_rPort_3_backpressure, // @[:@18409.4]
  output [31:0] io_rPort_3_output_0, // @[:@18409.4]
  input  [1:0]  io_rPort_2_banks_1, // @[:@18409.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@18409.4]
  input  [9:0]  io_rPort_2_ofs_0, // @[:@18409.4]
  input         io_rPort_2_en_0, // @[:@18409.4]
  input         io_rPort_2_backpressure, // @[:@18409.4]
  output [31:0] io_rPort_2_output_0, // @[:@18409.4]
  input  [1:0]  io_rPort_1_banks_1, // @[:@18409.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@18409.4]
  input  [9:0]  io_rPort_1_ofs_0, // @[:@18409.4]
  input         io_rPort_1_en_0, // @[:@18409.4]
  input         io_rPort_1_backpressure, // @[:@18409.4]
  output [31:0] io_rPort_1_output_0, // @[:@18409.4]
  input  [1:0]  io_rPort_0_banks_1, // @[:@18409.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@18409.4]
  input  [9:0]  io_rPort_0_ofs_0, // @[:@18409.4]
  input         io_rPort_0_en_0, // @[:@18409.4]
  input         io_rPort_0_backpressure, // @[:@18409.4]
  output [31:0] io_rPort_0_output_0, // @[:@18409.4]
  input  [1:0]  io_wPort_0_banks_1, // @[:@18409.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@18409.4]
  input  [9:0]  io_wPort_0_ofs_0, // @[:@18409.4]
  input  [31:0] io_wPort_0_data_0, // @[:@18409.4]
  input         io_wPort_0_en_0 // @[:@18409.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@18444.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@18444.4]
  wire [9:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18444.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18444.4]
  wire [9:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18444.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@18444.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@18444.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@18444.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@18460.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@18460.4]
  wire [9:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18460.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18460.4]
  wire [9:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18460.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@18460.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@18460.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@18460.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@18476.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@18476.4]
  wire [9:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18476.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18476.4]
  wire [9:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18476.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@18476.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@18476.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@18476.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@18492.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@18492.4]
  wire [9:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18492.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18492.4]
  wire [9:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18492.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@18492.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@18492.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@18492.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@18508.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@18508.4]
  wire [9:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18508.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18508.4]
  wire [9:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18508.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@18508.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@18508.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@18508.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@18524.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@18524.4]
  wire [9:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18524.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18524.4]
  wire [9:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18524.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@18524.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@18524.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@18524.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@18540.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@18540.4]
  wire [9:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18540.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18540.4]
  wire [9:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18540.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@18540.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@18540.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@18540.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@18556.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@18556.4]
  wire [9:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18556.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18556.4]
  wire [9:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18556.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@18556.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@18556.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@18556.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@18572.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@18572.4]
  wire [9:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18572.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18572.4]
  wire [9:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18572.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@18572.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@18572.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@18572.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@18588.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@18588.4]
  wire [9:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18588.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18588.4]
  wire [9:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18588.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@18588.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@18588.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@18588.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@18604.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@18604.4]
  wire [9:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18604.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18604.4]
  wire [9:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18604.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@18604.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@18604.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@18604.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@18620.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@18620.4]
  wire [9:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18620.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18620.4]
  wire [9:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18620.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@18620.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@18620.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@18620.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@19345.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@19345.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@19345.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@19345.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@19345.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@19353.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@19353.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@19353.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@19353.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@19353.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@19361.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@19361.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@19361.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@19361.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@19361.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@19369.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@19369.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@19369.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@19369.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@19369.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@19377.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@19377.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@19377.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@19377.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@19377.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@19385.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@19385.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@19385.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@19385.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@19385.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@19393.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@19393.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@19393.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@19393.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@19393.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@19401.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@19401.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@19401.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@19401.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@19401.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@19409.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@19409.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@19409.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@19409.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@19409.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@19417.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@19417.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@19417.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@19417.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@19417.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@19425.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@19425.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@19425.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@19425.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@19425.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@19433.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@19433.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@19433.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@19433.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@19433.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@19489.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@19489.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@19489.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@19489.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@19489.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@19497.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@19497.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@19497.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@19497.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@19497.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@19505.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@19505.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@19505.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@19505.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@19505.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@19513.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@19513.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@19513.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@19513.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@19513.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@19521.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@19521.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@19521.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@19521.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@19521.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@19529.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@19529.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@19529.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@19529.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@19529.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@19537.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@19537.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@19537.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@19537.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@19537.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@19545.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@19545.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@19545.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@19545.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@19545.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@19553.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@19553.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@19553.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@19553.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@19553.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@19561.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@19561.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@19561.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@19561.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@19561.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@19569.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@19569.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@19569.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@19569.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@19569.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@19577.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@19577.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@19577.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@19577.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@19577.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@19633.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@19633.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@19633.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@19633.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@19633.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@19641.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@19641.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@19641.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@19641.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@19641.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@19649.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@19649.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@19649.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@19649.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@19649.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@19657.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@19657.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@19657.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@19657.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@19657.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@19665.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@19665.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@19665.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@19665.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@19665.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@19673.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@19673.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@19673.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@19673.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@19673.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@19681.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@19681.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@19681.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@19681.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@19681.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@19689.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@19689.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@19689.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@19689.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@19689.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@19697.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@19697.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@19697.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@19697.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@19697.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@19705.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@19705.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@19705.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@19705.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@19705.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@19713.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@19713.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@19713.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@19713.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@19713.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@19721.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@19721.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@19721.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@19721.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@19721.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@19777.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@19777.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@19777.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@19777.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@19777.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@19785.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@19785.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@19785.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@19785.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@19785.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@19793.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@19793.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@19793.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@19793.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@19793.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@19801.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@19801.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@19801.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@19801.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@19801.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@19809.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@19809.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@19809.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@19809.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@19809.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@19817.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@19817.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@19817.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@19817.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@19817.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@19825.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@19825.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@19825.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@19825.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@19825.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@19833.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@19833.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@19833.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@19833.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@19833.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@19841.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@19841.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@19841.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@19841.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@19841.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@19849.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@19849.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@19849.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@19849.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@19849.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@19857.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@19857.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@19857.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@19857.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@19857.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@19865.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@19865.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@19865.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@19865.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@19865.4]
  wire  _T_166; // @[MemPrimitives.scala 82:210:@18636.4]
  wire  _T_168; // @[MemPrimitives.scala 82:210:@18637.4]
  wire  _T_169; // @[MemPrimitives.scala 82:228:@18638.4]
  wire  _T_170; // @[MemPrimitives.scala 83:102:@18639.4]
  wire [42:0] _T_172; // @[Cat.scala 30:58:@18641.4]
  wire  _T_179; // @[MemPrimitives.scala 82:210:@18649.4]
  wire  _T_180; // @[MemPrimitives.scala 82:228:@18650.4]
  wire  _T_181; // @[MemPrimitives.scala 83:102:@18651.4]
  wire [42:0] _T_183; // @[Cat.scala 30:58:@18653.4]
  wire  _T_190; // @[MemPrimitives.scala 82:210:@18661.4]
  wire  _T_191; // @[MemPrimitives.scala 82:228:@18662.4]
  wire  _T_192; // @[MemPrimitives.scala 83:102:@18663.4]
  wire [42:0] _T_194; // @[Cat.scala 30:58:@18665.4]
  wire  _T_199; // @[MemPrimitives.scala 82:210:@18672.4]
  wire  _T_202; // @[MemPrimitives.scala 82:228:@18674.4]
  wire  _T_203; // @[MemPrimitives.scala 83:102:@18675.4]
  wire [42:0] _T_205; // @[Cat.scala 30:58:@18677.4]
  wire  _T_213; // @[MemPrimitives.scala 82:228:@18686.4]
  wire  _T_214; // @[MemPrimitives.scala 83:102:@18687.4]
  wire [42:0] _T_216; // @[Cat.scala 30:58:@18689.4]
  wire  _T_224; // @[MemPrimitives.scala 82:228:@18698.4]
  wire  _T_225; // @[MemPrimitives.scala 83:102:@18699.4]
  wire [42:0] _T_227; // @[Cat.scala 30:58:@18701.4]
  wire  _T_232; // @[MemPrimitives.scala 82:210:@18708.4]
  wire  _T_235; // @[MemPrimitives.scala 82:228:@18710.4]
  wire  _T_236; // @[MemPrimitives.scala 83:102:@18711.4]
  wire [42:0] _T_238; // @[Cat.scala 30:58:@18713.4]
  wire  _T_246; // @[MemPrimitives.scala 82:228:@18722.4]
  wire  _T_247; // @[MemPrimitives.scala 83:102:@18723.4]
  wire [42:0] _T_249; // @[Cat.scala 30:58:@18725.4]
  wire  _T_257; // @[MemPrimitives.scala 82:228:@18734.4]
  wire  _T_258; // @[MemPrimitives.scala 83:102:@18735.4]
  wire [42:0] _T_260; // @[Cat.scala 30:58:@18737.4]
  wire  _T_265; // @[MemPrimitives.scala 82:210:@18744.4]
  wire  _T_268; // @[MemPrimitives.scala 82:228:@18746.4]
  wire  _T_269; // @[MemPrimitives.scala 83:102:@18747.4]
  wire [42:0] _T_271; // @[Cat.scala 30:58:@18749.4]
  wire  _T_279; // @[MemPrimitives.scala 82:228:@18758.4]
  wire  _T_280; // @[MemPrimitives.scala 83:102:@18759.4]
  wire [42:0] _T_282; // @[Cat.scala 30:58:@18761.4]
  wire  _T_290; // @[MemPrimitives.scala 82:228:@18770.4]
  wire  _T_291; // @[MemPrimitives.scala 83:102:@18771.4]
  wire [42:0] _T_293; // @[Cat.scala 30:58:@18773.4]
  wire  _T_298; // @[MemPrimitives.scala 110:210:@18780.4]
  wire  _T_300; // @[MemPrimitives.scala 110:210:@18781.4]
  wire  _T_301; // @[MemPrimitives.scala 110:228:@18782.4]
  wire  _T_304; // @[MemPrimitives.scala 110:210:@18784.4]
  wire  _T_306; // @[MemPrimitives.scala 110:210:@18785.4]
  wire  _T_307; // @[MemPrimitives.scala 110:228:@18786.4]
  wire  _T_310; // @[MemPrimitives.scala 110:210:@18788.4]
  wire  _T_312; // @[MemPrimitives.scala 110:210:@18789.4]
  wire  _T_313; // @[MemPrimitives.scala 110:228:@18790.4]
  wire  _T_316; // @[MemPrimitives.scala 110:210:@18792.4]
  wire  _T_318; // @[MemPrimitives.scala 110:210:@18793.4]
  wire  _T_319; // @[MemPrimitives.scala 110:228:@18794.4]
  wire  _T_321; // @[MemPrimitives.scala 126:35:@18803.4]
  wire  _T_322; // @[MemPrimitives.scala 126:35:@18804.4]
  wire  _T_323; // @[MemPrimitives.scala 126:35:@18805.4]
  wire  _T_324; // @[MemPrimitives.scala 126:35:@18806.4]
  wire [11:0] _T_326; // @[Cat.scala 30:58:@18808.4]
  wire [11:0] _T_328; // @[Cat.scala 30:58:@18810.4]
  wire [11:0] _T_330; // @[Cat.scala 30:58:@18812.4]
  wire [11:0] _T_332; // @[Cat.scala 30:58:@18814.4]
  wire [11:0] _T_333; // @[Mux.scala 31:69:@18815.4]
  wire [11:0] _T_334; // @[Mux.scala 31:69:@18816.4]
  wire [11:0] _T_335; // @[Mux.scala 31:69:@18817.4]
  wire  _T_342; // @[MemPrimitives.scala 110:210:@18825.4]
  wire  _T_343; // @[MemPrimitives.scala 110:228:@18826.4]
  wire  _T_348; // @[MemPrimitives.scala 110:210:@18829.4]
  wire  _T_349; // @[MemPrimitives.scala 110:228:@18830.4]
  wire  _T_354; // @[MemPrimitives.scala 110:210:@18833.4]
  wire  _T_355; // @[MemPrimitives.scala 110:228:@18834.4]
  wire  _T_360; // @[MemPrimitives.scala 110:210:@18837.4]
  wire  _T_361; // @[MemPrimitives.scala 110:228:@18838.4]
  wire  _T_363; // @[MemPrimitives.scala 126:35:@18847.4]
  wire  _T_364; // @[MemPrimitives.scala 126:35:@18848.4]
  wire  _T_365; // @[MemPrimitives.scala 126:35:@18849.4]
  wire  _T_366; // @[MemPrimitives.scala 126:35:@18850.4]
  wire [11:0] _T_368; // @[Cat.scala 30:58:@18852.4]
  wire [11:0] _T_370; // @[Cat.scala 30:58:@18854.4]
  wire [11:0] _T_372; // @[Cat.scala 30:58:@18856.4]
  wire [11:0] _T_374; // @[Cat.scala 30:58:@18858.4]
  wire [11:0] _T_375; // @[Mux.scala 31:69:@18859.4]
  wire [11:0] _T_376; // @[Mux.scala 31:69:@18860.4]
  wire [11:0] _T_377; // @[Mux.scala 31:69:@18861.4]
  wire  _T_384; // @[MemPrimitives.scala 110:210:@18869.4]
  wire  _T_385; // @[MemPrimitives.scala 110:228:@18870.4]
  wire  _T_390; // @[MemPrimitives.scala 110:210:@18873.4]
  wire  _T_391; // @[MemPrimitives.scala 110:228:@18874.4]
  wire  _T_396; // @[MemPrimitives.scala 110:210:@18877.4]
  wire  _T_397; // @[MemPrimitives.scala 110:228:@18878.4]
  wire  _T_402; // @[MemPrimitives.scala 110:210:@18881.4]
  wire  _T_403; // @[MemPrimitives.scala 110:228:@18882.4]
  wire  _T_405; // @[MemPrimitives.scala 126:35:@18891.4]
  wire  _T_406; // @[MemPrimitives.scala 126:35:@18892.4]
  wire  _T_407; // @[MemPrimitives.scala 126:35:@18893.4]
  wire  _T_408; // @[MemPrimitives.scala 126:35:@18894.4]
  wire [11:0] _T_410; // @[Cat.scala 30:58:@18896.4]
  wire [11:0] _T_412; // @[Cat.scala 30:58:@18898.4]
  wire [11:0] _T_414; // @[Cat.scala 30:58:@18900.4]
  wire [11:0] _T_416; // @[Cat.scala 30:58:@18902.4]
  wire [11:0] _T_417; // @[Mux.scala 31:69:@18903.4]
  wire [11:0] _T_418; // @[Mux.scala 31:69:@18904.4]
  wire [11:0] _T_419; // @[Mux.scala 31:69:@18905.4]
  wire  _T_424; // @[MemPrimitives.scala 110:210:@18912.4]
  wire  _T_427; // @[MemPrimitives.scala 110:228:@18914.4]
  wire  _T_430; // @[MemPrimitives.scala 110:210:@18916.4]
  wire  _T_433; // @[MemPrimitives.scala 110:228:@18918.4]
  wire  _T_436; // @[MemPrimitives.scala 110:210:@18920.4]
  wire  _T_439; // @[MemPrimitives.scala 110:228:@18922.4]
  wire  _T_442; // @[MemPrimitives.scala 110:210:@18924.4]
  wire  _T_445; // @[MemPrimitives.scala 110:228:@18926.4]
  wire  _T_447; // @[MemPrimitives.scala 126:35:@18935.4]
  wire  _T_448; // @[MemPrimitives.scala 126:35:@18936.4]
  wire  _T_449; // @[MemPrimitives.scala 126:35:@18937.4]
  wire  _T_450; // @[MemPrimitives.scala 126:35:@18938.4]
  wire [11:0] _T_452; // @[Cat.scala 30:58:@18940.4]
  wire [11:0] _T_454; // @[Cat.scala 30:58:@18942.4]
  wire [11:0] _T_456; // @[Cat.scala 30:58:@18944.4]
  wire [11:0] _T_458; // @[Cat.scala 30:58:@18946.4]
  wire [11:0] _T_459; // @[Mux.scala 31:69:@18947.4]
  wire [11:0] _T_460; // @[Mux.scala 31:69:@18948.4]
  wire [11:0] _T_461; // @[Mux.scala 31:69:@18949.4]
  wire  _T_469; // @[MemPrimitives.scala 110:228:@18958.4]
  wire  _T_475; // @[MemPrimitives.scala 110:228:@18962.4]
  wire  _T_481; // @[MemPrimitives.scala 110:228:@18966.4]
  wire  _T_487; // @[MemPrimitives.scala 110:228:@18970.4]
  wire  _T_489; // @[MemPrimitives.scala 126:35:@18979.4]
  wire  _T_490; // @[MemPrimitives.scala 126:35:@18980.4]
  wire  _T_491; // @[MemPrimitives.scala 126:35:@18981.4]
  wire  _T_492; // @[MemPrimitives.scala 126:35:@18982.4]
  wire [11:0] _T_494; // @[Cat.scala 30:58:@18984.4]
  wire [11:0] _T_496; // @[Cat.scala 30:58:@18986.4]
  wire [11:0] _T_498; // @[Cat.scala 30:58:@18988.4]
  wire [11:0] _T_500; // @[Cat.scala 30:58:@18990.4]
  wire [11:0] _T_501; // @[Mux.scala 31:69:@18991.4]
  wire [11:0] _T_502; // @[Mux.scala 31:69:@18992.4]
  wire [11:0] _T_503; // @[Mux.scala 31:69:@18993.4]
  wire  _T_511; // @[MemPrimitives.scala 110:228:@19002.4]
  wire  _T_517; // @[MemPrimitives.scala 110:228:@19006.4]
  wire  _T_523; // @[MemPrimitives.scala 110:228:@19010.4]
  wire  _T_529; // @[MemPrimitives.scala 110:228:@19014.4]
  wire  _T_531; // @[MemPrimitives.scala 126:35:@19023.4]
  wire  _T_532; // @[MemPrimitives.scala 126:35:@19024.4]
  wire  _T_533; // @[MemPrimitives.scala 126:35:@19025.4]
  wire  _T_534; // @[MemPrimitives.scala 126:35:@19026.4]
  wire [11:0] _T_536; // @[Cat.scala 30:58:@19028.4]
  wire [11:0] _T_538; // @[Cat.scala 30:58:@19030.4]
  wire [11:0] _T_540; // @[Cat.scala 30:58:@19032.4]
  wire [11:0] _T_542; // @[Cat.scala 30:58:@19034.4]
  wire [11:0] _T_543; // @[Mux.scala 31:69:@19035.4]
  wire [11:0] _T_544; // @[Mux.scala 31:69:@19036.4]
  wire [11:0] _T_545; // @[Mux.scala 31:69:@19037.4]
  wire  _T_550; // @[MemPrimitives.scala 110:210:@19044.4]
  wire  _T_553; // @[MemPrimitives.scala 110:228:@19046.4]
  wire  _T_556; // @[MemPrimitives.scala 110:210:@19048.4]
  wire  _T_559; // @[MemPrimitives.scala 110:228:@19050.4]
  wire  _T_562; // @[MemPrimitives.scala 110:210:@19052.4]
  wire  _T_565; // @[MemPrimitives.scala 110:228:@19054.4]
  wire  _T_568; // @[MemPrimitives.scala 110:210:@19056.4]
  wire  _T_571; // @[MemPrimitives.scala 110:228:@19058.4]
  wire  _T_573; // @[MemPrimitives.scala 126:35:@19067.4]
  wire  _T_574; // @[MemPrimitives.scala 126:35:@19068.4]
  wire  _T_575; // @[MemPrimitives.scala 126:35:@19069.4]
  wire  _T_576; // @[MemPrimitives.scala 126:35:@19070.4]
  wire [11:0] _T_578; // @[Cat.scala 30:58:@19072.4]
  wire [11:0] _T_580; // @[Cat.scala 30:58:@19074.4]
  wire [11:0] _T_582; // @[Cat.scala 30:58:@19076.4]
  wire [11:0] _T_584; // @[Cat.scala 30:58:@19078.4]
  wire [11:0] _T_585; // @[Mux.scala 31:69:@19079.4]
  wire [11:0] _T_586; // @[Mux.scala 31:69:@19080.4]
  wire [11:0] _T_587; // @[Mux.scala 31:69:@19081.4]
  wire  _T_595; // @[MemPrimitives.scala 110:228:@19090.4]
  wire  _T_601; // @[MemPrimitives.scala 110:228:@19094.4]
  wire  _T_607; // @[MemPrimitives.scala 110:228:@19098.4]
  wire  _T_613; // @[MemPrimitives.scala 110:228:@19102.4]
  wire  _T_615; // @[MemPrimitives.scala 126:35:@19111.4]
  wire  _T_616; // @[MemPrimitives.scala 126:35:@19112.4]
  wire  _T_617; // @[MemPrimitives.scala 126:35:@19113.4]
  wire  _T_618; // @[MemPrimitives.scala 126:35:@19114.4]
  wire [11:0] _T_620; // @[Cat.scala 30:58:@19116.4]
  wire [11:0] _T_622; // @[Cat.scala 30:58:@19118.4]
  wire [11:0] _T_624; // @[Cat.scala 30:58:@19120.4]
  wire [11:0] _T_626; // @[Cat.scala 30:58:@19122.4]
  wire [11:0] _T_627; // @[Mux.scala 31:69:@19123.4]
  wire [11:0] _T_628; // @[Mux.scala 31:69:@19124.4]
  wire [11:0] _T_629; // @[Mux.scala 31:69:@19125.4]
  wire  _T_637; // @[MemPrimitives.scala 110:228:@19134.4]
  wire  _T_643; // @[MemPrimitives.scala 110:228:@19138.4]
  wire  _T_649; // @[MemPrimitives.scala 110:228:@19142.4]
  wire  _T_655; // @[MemPrimitives.scala 110:228:@19146.4]
  wire  _T_657; // @[MemPrimitives.scala 126:35:@19155.4]
  wire  _T_658; // @[MemPrimitives.scala 126:35:@19156.4]
  wire  _T_659; // @[MemPrimitives.scala 126:35:@19157.4]
  wire  _T_660; // @[MemPrimitives.scala 126:35:@19158.4]
  wire [11:0] _T_662; // @[Cat.scala 30:58:@19160.4]
  wire [11:0] _T_664; // @[Cat.scala 30:58:@19162.4]
  wire [11:0] _T_666; // @[Cat.scala 30:58:@19164.4]
  wire [11:0] _T_668; // @[Cat.scala 30:58:@19166.4]
  wire [11:0] _T_669; // @[Mux.scala 31:69:@19167.4]
  wire [11:0] _T_670; // @[Mux.scala 31:69:@19168.4]
  wire [11:0] _T_671; // @[Mux.scala 31:69:@19169.4]
  wire  _T_676; // @[MemPrimitives.scala 110:210:@19176.4]
  wire  _T_679; // @[MemPrimitives.scala 110:228:@19178.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@19180.4]
  wire  _T_685; // @[MemPrimitives.scala 110:228:@19182.4]
  wire  _T_688; // @[MemPrimitives.scala 110:210:@19184.4]
  wire  _T_691; // @[MemPrimitives.scala 110:228:@19186.4]
  wire  _T_694; // @[MemPrimitives.scala 110:210:@19188.4]
  wire  _T_697; // @[MemPrimitives.scala 110:228:@19190.4]
  wire  _T_699; // @[MemPrimitives.scala 126:35:@19199.4]
  wire  _T_700; // @[MemPrimitives.scala 126:35:@19200.4]
  wire  _T_701; // @[MemPrimitives.scala 126:35:@19201.4]
  wire  _T_702; // @[MemPrimitives.scala 126:35:@19202.4]
  wire [11:0] _T_704; // @[Cat.scala 30:58:@19204.4]
  wire [11:0] _T_706; // @[Cat.scala 30:58:@19206.4]
  wire [11:0] _T_708; // @[Cat.scala 30:58:@19208.4]
  wire [11:0] _T_710; // @[Cat.scala 30:58:@19210.4]
  wire [11:0] _T_711; // @[Mux.scala 31:69:@19211.4]
  wire [11:0] _T_712; // @[Mux.scala 31:69:@19212.4]
  wire [11:0] _T_713; // @[Mux.scala 31:69:@19213.4]
  wire  _T_721; // @[MemPrimitives.scala 110:228:@19222.4]
  wire  _T_727; // @[MemPrimitives.scala 110:228:@19226.4]
  wire  _T_733; // @[MemPrimitives.scala 110:228:@19230.4]
  wire  _T_739; // @[MemPrimitives.scala 110:228:@19234.4]
  wire  _T_741; // @[MemPrimitives.scala 126:35:@19243.4]
  wire  _T_742; // @[MemPrimitives.scala 126:35:@19244.4]
  wire  _T_743; // @[MemPrimitives.scala 126:35:@19245.4]
  wire  _T_744; // @[MemPrimitives.scala 126:35:@19246.4]
  wire [11:0] _T_746; // @[Cat.scala 30:58:@19248.4]
  wire [11:0] _T_748; // @[Cat.scala 30:58:@19250.4]
  wire [11:0] _T_750; // @[Cat.scala 30:58:@19252.4]
  wire [11:0] _T_752; // @[Cat.scala 30:58:@19254.4]
  wire [11:0] _T_753; // @[Mux.scala 31:69:@19255.4]
  wire [11:0] _T_754; // @[Mux.scala 31:69:@19256.4]
  wire [11:0] _T_755; // @[Mux.scala 31:69:@19257.4]
  wire  _T_763; // @[MemPrimitives.scala 110:228:@19266.4]
  wire  _T_769; // @[MemPrimitives.scala 110:228:@19270.4]
  wire  _T_775; // @[MemPrimitives.scala 110:228:@19274.4]
  wire  _T_781; // @[MemPrimitives.scala 110:228:@19278.4]
  wire  _T_783; // @[MemPrimitives.scala 126:35:@19287.4]
  wire  _T_784; // @[MemPrimitives.scala 126:35:@19288.4]
  wire  _T_785; // @[MemPrimitives.scala 126:35:@19289.4]
  wire  _T_786; // @[MemPrimitives.scala 126:35:@19290.4]
  wire [11:0] _T_788; // @[Cat.scala 30:58:@19292.4]
  wire [11:0] _T_790; // @[Cat.scala 30:58:@19294.4]
  wire [11:0] _T_792; // @[Cat.scala 30:58:@19296.4]
  wire [11:0] _T_794; // @[Cat.scala 30:58:@19298.4]
  wire [11:0] _T_795; // @[Mux.scala 31:69:@19299.4]
  wire [11:0] _T_796; // @[Mux.scala 31:69:@19300.4]
  wire [11:0] _T_797; // @[Mux.scala 31:69:@19301.4]
  wire  _T_893; // @[package.scala 96:25:@19430.4 package.scala 96:25:@19431.4]
  wire [31:0] _T_897; // @[Mux.scala 31:69:@19440.4]
  wire  _T_890; // @[package.scala 96:25:@19422.4 package.scala 96:25:@19423.4]
  wire [31:0] _T_898; // @[Mux.scala 31:69:@19441.4]
  wire  _T_887; // @[package.scala 96:25:@19414.4 package.scala 96:25:@19415.4]
  wire [31:0] _T_899; // @[Mux.scala 31:69:@19442.4]
  wire  _T_884; // @[package.scala 96:25:@19406.4 package.scala 96:25:@19407.4]
  wire [31:0] _T_900; // @[Mux.scala 31:69:@19443.4]
  wire  _T_881; // @[package.scala 96:25:@19398.4 package.scala 96:25:@19399.4]
  wire [31:0] _T_901; // @[Mux.scala 31:69:@19444.4]
  wire  _T_878; // @[package.scala 96:25:@19390.4 package.scala 96:25:@19391.4]
  wire [31:0] _T_902; // @[Mux.scala 31:69:@19445.4]
  wire  _T_875; // @[package.scala 96:25:@19382.4 package.scala 96:25:@19383.4]
  wire [31:0] _T_903; // @[Mux.scala 31:69:@19446.4]
  wire  _T_872; // @[package.scala 96:25:@19374.4 package.scala 96:25:@19375.4]
  wire [31:0] _T_904; // @[Mux.scala 31:69:@19447.4]
  wire  _T_869; // @[package.scala 96:25:@19366.4 package.scala 96:25:@19367.4]
  wire [31:0] _T_905; // @[Mux.scala 31:69:@19448.4]
  wire  _T_866; // @[package.scala 96:25:@19358.4 package.scala 96:25:@19359.4]
  wire [31:0] _T_906; // @[Mux.scala 31:69:@19449.4]
  wire  _T_863; // @[package.scala 96:25:@19350.4 package.scala 96:25:@19351.4]
  wire  _T_1000; // @[package.scala 96:25:@19574.4 package.scala 96:25:@19575.4]
  wire [31:0] _T_1004; // @[Mux.scala 31:69:@19584.4]
  wire  _T_997; // @[package.scala 96:25:@19566.4 package.scala 96:25:@19567.4]
  wire [31:0] _T_1005; // @[Mux.scala 31:69:@19585.4]
  wire  _T_994; // @[package.scala 96:25:@19558.4 package.scala 96:25:@19559.4]
  wire [31:0] _T_1006; // @[Mux.scala 31:69:@19586.4]
  wire  _T_991; // @[package.scala 96:25:@19550.4 package.scala 96:25:@19551.4]
  wire [31:0] _T_1007; // @[Mux.scala 31:69:@19587.4]
  wire  _T_988; // @[package.scala 96:25:@19542.4 package.scala 96:25:@19543.4]
  wire [31:0] _T_1008; // @[Mux.scala 31:69:@19588.4]
  wire  _T_985; // @[package.scala 96:25:@19534.4 package.scala 96:25:@19535.4]
  wire [31:0] _T_1009; // @[Mux.scala 31:69:@19589.4]
  wire  _T_982; // @[package.scala 96:25:@19526.4 package.scala 96:25:@19527.4]
  wire [31:0] _T_1010; // @[Mux.scala 31:69:@19590.4]
  wire  _T_979; // @[package.scala 96:25:@19518.4 package.scala 96:25:@19519.4]
  wire [31:0] _T_1011; // @[Mux.scala 31:69:@19591.4]
  wire  _T_976; // @[package.scala 96:25:@19510.4 package.scala 96:25:@19511.4]
  wire [31:0] _T_1012; // @[Mux.scala 31:69:@19592.4]
  wire  _T_973; // @[package.scala 96:25:@19502.4 package.scala 96:25:@19503.4]
  wire [31:0] _T_1013; // @[Mux.scala 31:69:@19593.4]
  wire  _T_970; // @[package.scala 96:25:@19494.4 package.scala 96:25:@19495.4]
  wire  _T_1107; // @[package.scala 96:25:@19718.4 package.scala 96:25:@19719.4]
  wire [31:0] _T_1111; // @[Mux.scala 31:69:@19728.4]
  wire  _T_1104; // @[package.scala 96:25:@19710.4 package.scala 96:25:@19711.4]
  wire [31:0] _T_1112; // @[Mux.scala 31:69:@19729.4]
  wire  _T_1101; // @[package.scala 96:25:@19702.4 package.scala 96:25:@19703.4]
  wire [31:0] _T_1113; // @[Mux.scala 31:69:@19730.4]
  wire  _T_1098; // @[package.scala 96:25:@19694.4 package.scala 96:25:@19695.4]
  wire [31:0] _T_1114; // @[Mux.scala 31:69:@19731.4]
  wire  _T_1095; // @[package.scala 96:25:@19686.4 package.scala 96:25:@19687.4]
  wire [31:0] _T_1115; // @[Mux.scala 31:69:@19732.4]
  wire  _T_1092; // @[package.scala 96:25:@19678.4 package.scala 96:25:@19679.4]
  wire [31:0] _T_1116; // @[Mux.scala 31:69:@19733.4]
  wire  _T_1089; // @[package.scala 96:25:@19670.4 package.scala 96:25:@19671.4]
  wire [31:0] _T_1117; // @[Mux.scala 31:69:@19734.4]
  wire  _T_1086; // @[package.scala 96:25:@19662.4 package.scala 96:25:@19663.4]
  wire [31:0] _T_1118; // @[Mux.scala 31:69:@19735.4]
  wire  _T_1083; // @[package.scala 96:25:@19654.4 package.scala 96:25:@19655.4]
  wire [31:0] _T_1119; // @[Mux.scala 31:69:@19736.4]
  wire  _T_1080; // @[package.scala 96:25:@19646.4 package.scala 96:25:@19647.4]
  wire [31:0] _T_1120; // @[Mux.scala 31:69:@19737.4]
  wire  _T_1077; // @[package.scala 96:25:@19638.4 package.scala 96:25:@19639.4]
  wire  _T_1214; // @[package.scala 96:25:@19862.4 package.scala 96:25:@19863.4]
  wire [31:0] _T_1218; // @[Mux.scala 31:69:@19872.4]
  wire  _T_1211; // @[package.scala 96:25:@19854.4 package.scala 96:25:@19855.4]
  wire [31:0] _T_1219; // @[Mux.scala 31:69:@19873.4]
  wire  _T_1208; // @[package.scala 96:25:@19846.4 package.scala 96:25:@19847.4]
  wire [31:0] _T_1220; // @[Mux.scala 31:69:@19874.4]
  wire  _T_1205; // @[package.scala 96:25:@19838.4 package.scala 96:25:@19839.4]
  wire [31:0] _T_1221; // @[Mux.scala 31:69:@19875.4]
  wire  _T_1202; // @[package.scala 96:25:@19830.4 package.scala 96:25:@19831.4]
  wire [31:0] _T_1222; // @[Mux.scala 31:69:@19876.4]
  wire  _T_1199; // @[package.scala 96:25:@19822.4 package.scala 96:25:@19823.4]
  wire [31:0] _T_1223; // @[Mux.scala 31:69:@19877.4]
  wire  _T_1196; // @[package.scala 96:25:@19814.4 package.scala 96:25:@19815.4]
  wire [31:0] _T_1224; // @[Mux.scala 31:69:@19878.4]
  wire  _T_1193; // @[package.scala 96:25:@19806.4 package.scala 96:25:@19807.4]
  wire [31:0] _T_1225; // @[Mux.scala 31:69:@19879.4]
  wire  _T_1190; // @[package.scala 96:25:@19798.4 package.scala 96:25:@19799.4]
  wire [31:0] _T_1226; // @[Mux.scala 31:69:@19880.4]
  wire  _T_1187; // @[package.scala 96:25:@19790.4 package.scala 96:25:@19791.4]
  wire [31:0] _T_1227; // @[Mux.scala 31:69:@19881.4]
  wire  _T_1184; // @[package.scala 96:25:@19782.4 package.scala 96:25:@19783.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@18444.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@18460.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@18476.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@18492.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@18508.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@18524.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@18540.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@18556.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@18572.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@18588.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@18604.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@18620.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  StickySelects_13 StickySelects ( // @[MemPrimitives.scala 124:33:@18796.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3)
  );
  StickySelects_13 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@18840.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3)
  );
  StickySelects_13 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@18884.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3)
  );
  StickySelects_13 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@18928.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3)
  );
  StickySelects_13 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@18972.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3)
  );
  StickySelects_13 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@19016.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3)
  );
  StickySelects_13 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@19060.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3)
  );
  StickySelects_13 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@19104.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3)
  );
  StickySelects_13 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@19148.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3)
  );
  StickySelects_13 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@19192.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3)
  );
  StickySelects_13 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@19236.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3)
  );
  StickySelects_13 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@19280.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@19345.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@19353.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@19361.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@19369.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@19377.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@19385.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@19393.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@19401.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@19409.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@19417.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@19425.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@19433.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@19489.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@19497.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@19505.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@19513.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@19521.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@19529.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@19537.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@19545.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@19553.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@19561.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@19569.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@19577.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@19633.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@19641.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@19649.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@19657.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@19665.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@19673.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@19681.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@19689.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@19697.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@19705.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@19713.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@19721.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@19777.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@19785.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@19793.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@19801.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@19809.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@19817.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@19825.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@19833.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@19841.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@19849.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@19857.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@19865.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  assign _T_166 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@18636.4]
  assign _T_168 = io_wPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 82:210:@18637.4]
  assign _T_169 = _T_166 & _T_168; // @[MemPrimitives.scala 82:228:@18638.4]
  assign _T_170 = io_wPort_0_en_0 & _T_169; // @[MemPrimitives.scala 83:102:@18639.4]
  assign _T_172 = {_T_170,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18641.4]
  assign _T_179 = io_wPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 82:210:@18649.4]
  assign _T_180 = _T_166 & _T_179; // @[MemPrimitives.scala 82:228:@18650.4]
  assign _T_181 = io_wPort_0_en_0 & _T_180; // @[MemPrimitives.scala 83:102:@18651.4]
  assign _T_183 = {_T_181,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18653.4]
  assign _T_190 = io_wPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 82:210:@18661.4]
  assign _T_191 = _T_166 & _T_190; // @[MemPrimitives.scala 82:228:@18662.4]
  assign _T_192 = io_wPort_0_en_0 & _T_191; // @[MemPrimitives.scala 83:102:@18663.4]
  assign _T_194 = {_T_192,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18665.4]
  assign _T_199 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@18672.4]
  assign _T_202 = _T_199 & _T_168; // @[MemPrimitives.scala 82:228:@18674.4]
  assign _T_203 = io_wPort_0_en_0 & _T_202; // @[MemPrimitives.scala 83:102:@18675.4]
  assign _T_205 = {_T_203,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18677.4]
  assign _T_213 = _T_199 & _T_179; // @[MemPrimitives.scala 82:228:@18686.4]
  assign _T_214 = io_wPort_0_en_0 & _T_213; // @[MemPrimitives.scala 83:102:@18687.4]
  assign _T_216 = {_T_214,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18689.4]
  assign _T_224 = _T_199 & _T_190; // @[MemPrimitives.scala 82:228:@18698.4]
  assign _T_225 = io_wPort_0_en_0 & _T_224; // @[MemPrimitives.scala 83:102:@18699.4]
  assign _T_227 = {_T_225,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18701.4]
  assign _T_232 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@18708.4]
  assign _T_235 = _T_232 & _T_168; // @[MemPrimitives.scala 82:228:@18710.4]
  assign _T_236 = io_wPort_0_en_0 & _T_235; // @[MemPrimitives.scala 83:102:@18711.4]
  assign _T_238 = {_T_236,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18713.4]
  assign _T_246 = _T_232 & _T_179; // @[MemPrimitives.scala 82:228:@18722.4]
  assign _T_247 = io_wPort_0_en_0 & _T_246; // @[MemPrimitives.scala 83:102:@18723.4]
  assign _T_249 = {_T_247,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18725.4]
  assign _T_257 = _T_232 & _T_190; // @[MemPrimitives.scala 82:228:@18734.4]
  assign _T_258 = io_wPort_0_en_0 & _T_257; // @[MemPrimitives.scala 83:102:@18735.4]
  assign _T_260 = {_T_258,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18737.4]
  assign _T_265 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@18744.4]
  assign _T_268 = _T_265 & _T_168; // @[MemPrimitives.scala 82:228:@18746.4]
  assign _T_269 = io_wPort_0_en_0 & _T_268; // @[MemPrimitives.scala 83:102:@18747.4]
  assign _T_271 = {_T_269,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18749.4]
  assign _T_279 = _T_265 & _T_179; // @[MemPrimitives.scala 82:228:@18758.4]
  assign _T_280 = io_wPort_0_en_0 & _T_279; // @[MemPrimitives.scala 83:102:@18759.4]
  assign _T_282 = {_T_280,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18761.4]
  assign _T_290 = _T_265 & _T_190; // @[MemPrimitives.scala 82:228:@18770.4]
  assign _T_291 = io_wPort_0_en_0 & _T_290; // @[MemPrimitives.scala 83:102:@18771.4]
  assign _T_293 = {_T_291,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18773.4]
  assign _T_298 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@18780.4]
  assign _T_300 = io_rPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@18781.4]
  assign _T_301 = _T_298 & _T_300; // @[MemPrimitives.scala 110:228:@18782.4]
  assign _T_304 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@18784.4]
  assign _T_306 = io_rPort_1_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@18785.4]
  assign _T_307 = _T_304 & _T_306; // @[MemPrimitives.scala 110:228:@18786.4]
  assign _T_310 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@18788.4]
  assign _T_312 = io_rPort_2_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@18789.4]
  assign _T_313 = _T_310 & _T_312; // @[MemPrimitives.scala 110:228:@18790.4]
  assign _T_316 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@18792.4]
  assign _T_318 = io_rPort_3_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@18793.4]
  assign _T_319 = _T_316 & _T_318; // @[MemPrimitives.scala 110:228:@18794.4]
  assign _T_321 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@18803.4]
  assign _T_322 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@18804.4]
  assign _T_323 = StickySelects_io_outs_2; // @[MemPrimitives.scala 126:35:@18805.4]
  assign _T_324 = StickySelects_io_outs_3; // @[MemPrimitives.scala 126:35:@18806.4]
  assign _T_326 = {_T_321,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@18808.4]
  assign _T_328 = {_T_322,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@18810.4]
  assign _T_330 = {_T_323,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@18812.4]
  assign _T_332 = {_T_324,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@18814.4]
  assign _T_333 = _T_323 ? _T_330 : _T_332; // @[Mux.scala 31:69:@18815.4]
  assign _T_334 = _T_322 ? _T_328 : _T_333; // @[Mux.scala 31:69:@18816.4]
  assign _T_335 = _T_321 ? _T_326 : _T_334; // @[Mux.scala 31:69:@18817.4]
  assign _T_342 = io_rPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@18825.4]
  assign _T_343 = _T_298 & _T_342; // @[MemPrimitives.scala 110:228:@18826.4]
  assign _T_348 = io_rPort_1_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@18829.4]
  assign _T_349 = _T_304 & _T_348; // @[MemPrimitives.scala 110:228:@18830.4]
  assign _T_354 = io_rPort_2_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@18833.4]
  assign _T_355 = _T_310 & _T_354; // @[MemPrimitives.scala 110:228:@18834.4]
  assign _T_360 = io_rPort_3_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@18837.4]
  assign _T_361 = _T_316 & _T_360; // @[MemPrimitives.scala 110:228:@18838.4]
  assign _T_363 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@18847.4]
  assign _T_364 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@18848.4]
  assign _T_365 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@18849.4]
  assign _T_366 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@18850.4]
  assign _T_368 = {_T_363,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@18852.4]
  assign _T_370 = {_T_364,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@18854.4]
  assign _T_372 = {_T_365,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@18856.4]
  assign _T_374 = {_T_366,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@18858.4]
  assign _T_375 = _T_365 ? _T_372 : _T_374; // @[Mux.scala 31:69:@18859.4]
  assign _T_376 = _T_364 ? _T_370 : _T_375; // @[Mux.scala 31:69:@18860.4]
  assign _T_377 = _T_363 ? _T_368 : _T_376; // @[Mux.scala 31:69:@18861.4]
  assign _T_384 = io_rPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@18869.4]
  assign _T_385 = _T_298 & _T_384; // @[MemPrimitives.scala 110:228:@18870.4]
  assign _T_390 = io_rPort_1_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@18873.4]
  assign _T_391 = _T_304 & _T_390; // @[MemPrimitives.scala 110:228:@18874.4]
  assign _T_396 = io_rPort_2_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@18877.4]
  assign _T_397 = _T_310 & _T_396; // @[MemPrimitives.scala 110:228:@18878.4]
  assign _T_402 = io_rPort_3_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@18881.4]
  assign _T_403 = _T_316 & _T_402; // @[MemPrimitives.scala 110:228:@18882.4]
  assign _T_405 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@18891.4]
  assign _T_406 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@18892.4]
  assign _T_407 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 126:35:@18893.4]
  assign _T_408 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 126:35:@18894.4]
  assign _T_410 = {_T_405,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@18896.4]
  assign _T_412 = {_T_406,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@18898.4]
  assign _T_414 = {_T_407,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@18900.4]
  assign _T_416 = {_T_408,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@18902.4]
  assign _T_417 = _T_407 ? _T_414 : _T_416; // @[Mux.scala 31:69:@18903.4]
  assign _T_418 = _T_406 ? _T_412 : _T_417; // @[Mux.scala 31:69:@18904.4]
  assign _T_419 = _T_405 ? _T_410 : _T_418; // @[Mux.scala 31:69:@18905.4]
  assign _T_424 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@18912.4]
  assign _T_427 = _T_424 & _T_300; // @[MemPrimitives.scala 110:228:@18914.4]
  assign _T_430 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@18916.4]
  assign _T_433 = _T_430 & _T_306; // @[MemPrimitives.scala 110:228:@18918.4]
  assign _T_436 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@18920.4]
  assign _T_439 = _T_436 & _T_312; // @[MemPrimitives.scala 110:228:@18922.4]
  assign _T_442 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@18924.4]
  assign _T_445 = _T_442 & _T_318; // @[MemPrimitives.scala 110:228:@18926.4]
  assign _T_447 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@18935.4]
  assign _T_448 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@18936.4]
  assign _T_449 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@18937.4]
  assign _T_450 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@18938.4]
  assign _T_452 = {_T_447,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@18940.4]
  assign _T_454 = {_T_448,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@18942.4]
  assign _T_456 = {_T_449,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@18944.4]
  assign _T_458 = {_T_450,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@18946.4]
  assign _T_459 = _T_449 ? _T_456 : _T_458; // @[Mux.scala 31:69:@18947.4]
  assign _T_460 = _T_448 ? _T_454 : _T_459; // @[Mux.scala 31:69:@18948.4]
  assign _T_461 = _T_447 ? _T_452 : _T_460; // @[Mux.scala 31:69:@18949.4]
  assign _T_469 = _T_424 & _T_342; // @[MemPrimitives.scala 110:228:@18958.4]
  assign _T_475 = _T_430 & _T_348; // @[MemPrimitives.scala 110:228:@18962.4]
  assign _T_481 = _T_436 & _T_354; // @[MemPrimitives.scala 110:228:@18966.4]
  assign _T_487 = _T_442 & _T_360; // @[MemPrimitives.scala 110:228:@18970.4]
  assign _T_489 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@18979.4]
  assign _T_490 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@18980.4]
  assign _T_491 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 126:35:@18981.4]
  assign _T_492 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 126:35:@18982.4]
  assign _T_494 = {_T_489,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@18984.4]
  assign _T_496 = {_T_490,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@18986.4]
  assign _T_498 = {_T_491,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@18988.4]
  assign _T_500 = {_T_492,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@18990.4]
  assign _T_501 = _T_491 ? _T_498 : _T_500; // @[Mux.scala 31:69:@18991.4]
  assign _T_502 = _T_490 ? _T_496 : _T_501; // @[Mux.scala 31:69:@18992.4]
  assign _T_503 = _T_489 ? _T_494 : _T_502; // @[Mux.scala 31:69:@18993.4]
  assign _T_511 = _T_424 & _T_384; // @[MemPrimitives.scala 110:228:@19002.4]
  assign _T_517 = _T_430 & _T_390; // @[MemPrimitives.scala 110:228:@19006.4]
  assign _T_523 = _T_436 & _T_396; // @[MemPrimitives.scala 110:228:@19010.4]
  assign _T_529 = _T_442 & _T_402; // @[MemPrimitives.scala 110:228:@19014.4]
  assign _T_531 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@19023.4]
  assign _T_532 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@19024.4]
  assign _T_533 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@19025.4]
  assign _T_534 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@19026.4]
  assign _T_536 = {_T_531,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19028.4]
  assign _T_538 = {_T_532,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19030.4]
  assign _T_540 = {_T_533,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19032.4]
  assign _T_542 = {_T_534,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19034.4]
  assign _T_543 = _T_533 ? _T_540 : _T_542; // @[Mux.scala 31:69:@19035.4]
  assign _T_544 = _T_532 ? _T_538 : _T_543; // @[Mux.scala 31:69:@19036.4]
  assign _T_545 = _T_531 ? _T_536 : _T_544; // @[Mux.scala 31:69:@19037.4]
  assign _T_550 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19044.4]
  assign _T_553 = _T_550 & _T_300; // @[MemPrimitives.scala 110:228:@19046.4]
  assign _T_556 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19048.4]
  assign _T_559 = _T_556 & _T_306; // @[MemPrimitives.scala 110:228:@19050.4]
  assign _T_562 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19052.4]
  assign _T_565 = _T_562 & _T_312; // @[MemPrimitives.scala 110:228:@19054.4]
  assign _T_568 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19056.4]
  assign _T_571 = _T_568 & _T_318; // @[MemPrimitives.scala 110:228:@19058.4]
  assign _T_573 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@19067.4]
  assign _T_574 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@19068.4]
  assign _T_575 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 126:35:@19069.4]
  assign _T_576 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 126:35:@19070.4]
  assign _T_578 = {_T_573,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19072.4]
  assign _T_580 = {_T_574,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19074.4]
  assign _T_582 = {_T_575,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19076.4]
  assign _T_584 = {_T_576,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19078.4]
  assign _T_585 = _T_575 ? _T_582 : _T_584; // @[Mux.scala 31:69:@19079.4]
  assign _T_586 = _T_574 ? _T_580 : _T_585; // @[Mux.scala 31:69:@19080.4]
  assign _T_587 = _T_573 ? _T_578 : _T_586; // @[Mux.scala 31:69:@19081.4]
  assign _T_595 = _T_550 & _T_342; // @[MemPrimitives.scala 110:228:@19090.4]
  assign _T_601 = _T_556 & _T_348; // @[MemPrimitives.scala 110:228:@19094.4]
  assign _T_607 = _T_562 & _T_354; // @[MemPrimitives.scala 110:228:@19098.4]
  assign _T_613 = _T_568 & _T_360; // @[MemPrimitives.scala 110:228:@19102.4]
  assign _T_615 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@19111.4]
  assign _T_616 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@19112.4]
  assign _T_617 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@19113.4]
  assign _T_618 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@19114.4]
  assign _T_620 = {_T_615,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19116.4]
  assign _T_622 = {_T_616,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19118.4]
  assign _T_624 = {_T_617,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19120.4]
  assign _T_626 = {_T_618,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19122.4]
  assign _T_627 = _T_617 ? _T_624 : _T_626; // @[Mux.scala 31:69:@19123.4]
  assign _T_628 = _T_616 ? _T_622 : _T_627; // @[Mux.scala 31:69:@19124.4]
  assign _T_629 = _T_615 ? _T_620 : _T_628; // @[Mux.scala 31:69:@19125.4]
  assign _T_637 = _T_550 & _T_384; // @[MemPrimitives.scala 110:228:@19134.4]
  assign _T_643 = _T_556 & _T_390; // @[MemPrimitives.scala 110:228:@19138.4]
  assign _T_649 = _T_562 & _T_396; // @[MemPrimitives.scala 110:228:@19142.4]
  assign _T_655 = _T_568 & _T_402; // @[MemPrimitives.scala 110:228:@19146.4]
  assign _T_657 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@19155.4]
  assign _T_658 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@19156.4]
  assign _T_659 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 126:35:@19157.4]
  assign _T_660 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 126:35:@19158.4]
  assign _T_662 = {_T_657,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19160.4]
  assign _T_664 = {_T_658,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19162.4]
  assign _T_666 = {_T_659,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19164.4]
  assign _T_668 = {_T_660,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19166.4]
  assign _T_669 = _T_659 ? _T_666 : _T_668; // @[Mux.scala 31:69:@19167.4]
  assign _T_670 = _T_658 ? _T_664 : _T_669; // @[Mux.scala 31:69:@19168.4]
  assign _T_671 = _T_657 ? _T_662 : _T_670; // @[Mux.scala 31:69:@19169.4]
  assign _T_676 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19176.4]
  assign _T_679 = _T_676 & _T_300; // @[MemPrimitives.scala 110:228:@19178.4]
  assign _T_682 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19180.4]
  assign _T_685 = _T_682 & _T_306; // @[MemPrimitives.scala 110:228:@19182.4]
  assign _T_688 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19184.4]
  assign _T_691 = _T_688 & _T_312; // @[MemPrimitives.scala 110:228:@19186.4]
  assign _T_694 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19188.4]
  assign _T_697 = _T_694 & _T_318; // @[MemPrimitives.scala 110:228:@19190.4]
  assign _T_699 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@19199.4]
  assign _T_700 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@19200.4]
  assign _T_701 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@19201.4]
  assign _T_702 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@19202.4]
  assign _T_704 = {_T_699,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19204.4]
  assign _T_706 = {_T_700,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19206.4]
  assign _T_708 = {_T_701,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19208.4]
  assign _T_710 = {_T_702,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19210.4]
  assign _T_711 = _T_701 ? _T_708 : _T_710; // @[Mux.scala 31:69:@19211.4]
  assign _T_712 = _T_700 ? _T_706 : _T_711; // @[Mux.scala 31:69:@19212.4]
  assign _T_713 = _T_699 ? _T_704 : _T_712; // @[Mux.scala 31:69:@19213.4]
  assign _T_721 = _T_676 & _T_342; // @[MemPrimitives.scala 110:228:@19222.4]
  assign _T_727 = _T_682 & _T_348; // @[MemPrimitives.scala 110:228:@19226.4]
  assign _T_733 = _T_688 & _T_354; // @[MemPrimitives.scala 110:228:@19230.4]
  assign _T_739 = _T_694 & _T_360; // @[MemPrimitives.scala 110:228:@19234.4]
  assign _T_741 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@19243.4]
  assign _T_742 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@19244.4]
  assign _T_743 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 126:35:@19245.4]
  assign _T_744 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 126:35:@19246.4]
  assign _T_746 = {_T_741,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19248.4]
  assign _T_748 = {_T_742,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19250.4]
  assign _T_750 = {_T_743,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19252.4]
  assign _T_752 = {_T_744,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19254.4]
  assign _T_753 = _T_743 ? _T_750 : _T_752; // @[Mux.scala 31:69:@19255.4]
  assign _T_754 = _T_742 ? _T_748 : _T_753; // @[Mux.scala 31:69:@19256.4]
  assign _T_755 = _T_741 ? _T_746 : _T_754; // @[Mux.scala 31:69:@19257.4]
  assign _T_763 = _T_676 & _T_384; // @[MemPrimitives.scala 110:228:@19266.4]
  assign _T_769 = _T_682 & _T_390; // @[MemPrimitives.scala 110:228:@19270.4]
  assign _T_775 = _T_688 & _T_396; // @[MemPrimitives.scala 110:228:@19274.4]
  assign _T_781 = _T_694 & _T_402; // @[MemPrimitives.scala 110:228:@19278.4]
  assign _T_783 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@19287.4]
  assign _T_784 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@19288.4]
  assign _T_785 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@19289.4]
  assign _T_786 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@19290.4]
  assign _T_788 = {_T_783,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19292.4]
  assign _T_790 = {_T_784,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19294.4]
  assign _T_792 = {_T_785,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19296.4]
  assign _T_794 = {_T_786,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19298.4]
  assign _T_795 = _T_785 ? _T_792 : _T_794; // @[Mux.scala 31:69:@19299.4]
  assign _T_796 = _T_784 ? _T_790 : _T_795; // @[Mux.scala 31:69:@19300.4]
  assign _T_797 = _T_783 ? _T_788 : _T_796; // @[Mux.scala 31:69:@19301.4]
  assign _T_893 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@19430.4 package.scala 96:25:@19431.4]
  assign _T_897 = _T_893 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@19440.4]
  assign _T_890 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@19422.4 package.scala 96:25:@19423.4]
  assign _T_898 = _T_890 ? Mem1D_9_io_output : _T_897; // @[Mux.scala 31:69:@19441.4]
  assign _T_887 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@19414.4 package.scala 96:25:@19415.4]
  assign _T_899 = _T_887 ? Mem1D_8_io_output : _T_898; // @[Mux.scala 31:69:@19442.4]
  assign _T_884 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@19406.4 package.scala 96:25:@19407.4]
  assign _T_900 = _T_884 ? Mem1D_7_io_output : _T_899; // @[Mux.scala 31:69:@19443.4]
  assign _T_881 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@19398.4 package.scala 96:25:@19399.4]
  assign _T_901 = _T_881 ? Mem1D_6_io_output : _T_900; // @[Mux.scala 31:69:@19444.4]
  assign _T_878 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@19390.4 package.scala 96:25:@19391.4]
  assign _T_902 = _T_878 ? Mem1D_5_io_output : _T_901; // @[Mux.scala 31:69:@19445.4]
  assign _T_875 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@19382.4 package.scala 96:25:@19383.4]
  assign _T_903 = _T_875 ? Mem1D_4_io_output : _T_902; // @[Mux.scala 31:69:@19446.4]
  assign _T_872 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@19374.4 package.scala 96:25:@19375.4]
  assign _T_904 = _T_872 ? Mem1D_3_io_output : _T_903; // @[Mux.scala 31:69:@19447.4]
  assign _T_869 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@19366.4 package.scala 96:25:@19367.4]
  assign _T_905 = _T_869 ? Mem1D_2_io_output : _T_904; // @[Mux.scala 31:69:@19448.4]
  assign _T_866 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@19358.4 package.scala 96:25:@19359.4]
  assign _T_906 = _T_866 ? Mem1D_1_io_output : _T_905; // @[Mux.scala 31:69:@19449.4]
  assign _T_863 = RetimeWrapper_io_out; // @[package.scala 96:25:@19350.4 package.scala 96:25:@19351.4]
  assign _T_1000 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@19574.4 package.scala 96:25:@19575.4]
  assign _T_1004 = _T_1000 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@19584.4]
  assign _T_997 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@19566.4 package.scala 96:25:@19567.4]
  assign _T_1005 = _T_997 ? Mem1D_9_io_output : _T_1004; // @[Mux.scala 31:69:@19585.4]
  assign _T_994 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@19558.4 package.scala 96:25:@19559.4]
  assign _T_1006 = _T_994 ? Mem1D_8_io_output : _T_1005; // @[Mux.scala 31:69:@19586.4]
  assign _T_991 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@19550.4 package.scala 96:25:@19551.4]
  assign _T_1007 = _T_991 ? Mem1D_7_io_output : _T_1006; // @[Mux.scala 31:69:@19587.4]
  assign _T_988 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@19542.4 package.scala 96:25:@19543.4]
  assign _T_1008 = _T_988 ? Mem1D_6_io_output : _T_1007; // @[Mux.scala 31:69:@19588.4]
  assign _T_985 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@19534.4 package.scala 96:25:@19535.4]
  assign _T_1009 = _T_985 ? Mem1D_5_io_output : _T_1008; // @[Mux.scala 31:69:@19589.4]
  assign _T_982 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@19526.4 package.scala 96:25:@19527.4]
  assign _T_1010 = _T_982 ? Mem1D_4_io_output : _T_1009; // @[Mux.scala 31:69:@19590.4]
  assign _T_979 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@19518.4 package.scala 96:25:@19519.4]
  assign _T_1011 = _T_979 ? Mem1D_3_io_output : _T_1010; // @[Mux.scala 31:69:@19591.4]
  assign _T_976 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@19510.4 package.scala 96:25:@19511.4]
  assign _T_1012 = _T_976 ? Mem1D_2_io_output : _T_1011; // @[Mux.scala 31:69:@19592.4]
  assign _T_973 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@19502.4 package.scala 96:25:@19503.4]
  assign _T_1013 = _T_973 ? Mem1D_1_io_output : _T_1012; // @[Mux.scala 31:69:@19593.4]
  assign _T_970 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@19494.4 package.scala 96:25:@19495.4]
  assign _T_1107 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@19718.4 package.scala 96:25:@19719.4]
  assign _T_1111 = _T_1107 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@19728.4]
  assign _T_1104 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@19710.4 package.scala 96:25:@19711.4]
  assign _T_1112 = _T_1104 ? Mem1D_9_io_output : _T_1111; // @[Mux.scala 31:69:@19729.4]
  assign _T_1101 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@19702.4 package.scala 96:25:@19703.4]
  assign _T_1113 = _T_1101 ? Mem1D_8_io_output : _T_1112; // @[Mux.scala 31:69:@19730.4]
  assign _T_1098 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@19694.4 package.scala 96:25:@19695.4]
  assign _T_1114 = _T_1098 ? Mem1D_7_io_output : _T_1113; // @[Mux.scala 31:69:@19731.4]
  assign _T_1095 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@19686.4 package.scala 96:25:@19687.4]
  assign _T_1115 = _T_1095 ? Mem1D_6_io_output : _T_1114; // @[Mux.scala 31:69:@19732.4]
  assign _T_1092 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@19678.4 package.scala 96:25:@19679.4]
  assign _T_1116 = _T_1092 ? Mem1D_5_io_output : _T_1115; // @[Mux.scala 31:69:@19733.4]
  assign _T_1089 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@19670.4 package.scala 96:25:@19671.4]
  assign _T_1117 = _T_1089 ? Mem1D_4_io_output : _T_1116; // @[Mux.scala 31:69:@19734.4]
  assign _T_1086 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@19662.4 package.scala 96:25:@19663.4]
  assign _T_1118 = _T_1086 ? Mem1D_3_io_output : _T_1117; // @[Mux.scala 31:69:@19735.4]
  assign _T_1083 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@19654.4 package.scala 96:25:@19655.4]
  assign _T_1119 = _T_1083 ? Mem1D_2_io_output : _T_1118; // @[Mux.scala 31:69:@19736.4]
  assign _T_1080 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@19646.4 package.scala 96:25:@19647.4]
  assign _T_1120 = _T_1080 ? Mem1D_1_io_output : _T_1119; // @[Mux.scala 31:69:@19737.4]
  assign _T_1077 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@19638.4 package.scala 96:25:@19639.4]
  assign _T_1214 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@19862.4 package.scala 96:25:@19863.4]
  assign _T_1218 = _T_1214 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@19872.4]
  assign _T_1211 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@19854.4 package.scala 96:25:@19855.4]
  assign _T_1219 = _T_1211 ? Mem1D_9_io_output : _T_1218; // @[Mux.scala 31:69:@19873.4]
  assign _T_1208 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@19846.4 package.scala 96:25:@19847.4]
  assign _T_1220 = _T_1208 ? Mem1D_8_io_output : _T_1219; // @[Mux.scala 31:69:@19874.4]
  assign _T_1205 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@19838.4 package.scala 96:25:@19839.4]
  assign _T_1221 = _T_1205 ? Mem1D_7_io_output : _T_1220; // @[Mux.scala 31:69:@19875.4]
  assign _T_1202 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@19830.4 package.scala 96:25:@19831.4]
  assign _T_1222 = _T_1202 ? Mem1D_6_io_output : _T_1221; // @[Mux.scala 31:69:@19876.4]
  assign _T_1199 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@19822.4 package.scala 96:25:@19823.4]
  assign _T_1223 = _T_1199 ? Mem1D_5_io_output : _T_1222; // @[Mux.scala 31:69:@19877.4]
  assign _T_1196 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@19814.4 package.scala 96:25:@19815.4]
  assign _T_1224 = _T_1196 ? Mem1D_4_io_output : _T_1223; // @[Mux.scala 31:69:@19878.4]
  assign _T_1193 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@19806.4 package.scala 96:25:@19807.4]
  assign _T_1225 = _T_1193 ? Mem1D_3_io_output : _T_1224; // @[Mux.scala 31:69:@19879.4]
  assign _T_1190 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@19798.4 package.scala 96:25:@19799.4]
  assign _T_1226 = _T_1190 ? Mem1D_2_io_output : _T_1225; // @[Mux.scala 31:69:@19880.4]
  assign _T_1187 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@19790.4 package.scala 96:25:@19791.4]
  assign _T_1227 = _T_1187 ? Mem1D_1_io_output : _T_1226; // @[Mux.scala 31:69:@19881.4]
  assign _T_1184 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@19782.4 package.scala 96:25:@19783.4]
  assign io_rPort_3_output_0 = _T_1184 ? Mem1D_io_output : _T_1227; // @[MemPrimitives.scala 152:13:@19883.4]
  assign io_rPort_2_output_0 = _T_1077 ? Mem1D_io_output : _T_1120; // @[MemPrimitives.scala 152:13:@19739.4]
  assign io_rPort_1_output_0 = _T_970 ? Mem1D_io_output : _T_1013; // @[MemPrimitives.scala 152:13:@19595.4]
  assign io_rPort_0_output_0 = _T_863 ? Mem1D_io_output : _T_906; // @[MemPrimitives.scala 152:13:@19451.4]
  assign Mem1D_clock = clock; // @[:@18445.4]
  assign Mem1D_reset = reset; // @[:@18446.4]
  assign Mem1D_io_r_ofs_0 = _T_335[9:0]; // @[MemPrimitives.scala 131:28:@18821.4]
  assign Mem1D_io_r_backpressure = _T_335[10]; // @[MemPrimitives.scala 132:32:@18822.4]
  assign Mem1D_io_w_ofs_0 = _T_172[9:0]; // @[MemPrimitives.scala 94:28:@18645.4]
  assign Mem1D_io_w_data_0 = _T_172[41:10]; // @[MemPrimitives.scala 95:29:@18646.4]
  assign Mem1D_io_w_en_0 = _T_172[42]; // @[MemPrimitives.scala 96:27:@18647.4]
  assign Mem1D_1_clock = clock; // @[:@18461.4]
  assign Mem1D_1_reset = reset; // @[:@18462.4]
  assign Mem1D_1_io_r_ofs_0 = _T_377[9:0]; // @[MemPrimitives.scala 131:28:@18865.4]
  assign Mem1D_1_io_r_backpressure = _T_377[10]; // @[MemPrimitives.scala 132:32:@18866.4]
  assign Mem1D_1_io_w_ofs_0 = _T_183[9:0]; // @[MemPrimitives.scala 94:28:@18657.4]
  assign Mem1D_1_io_w_data_0 = _T_183[41:10]; // @[MemPrimitives.scala 95:29:@18658.4]
  assign Mem1D_1_io_w_en_0 = _T_183[42]; // @[MemPrimitives.scala 96:27:@18659.4]
  assign Mem1D_2_clock = clock; // @[:@18477.4]
  assign Mem1D_2_reset = reset; // @[:@18478.4]
  assign Mem1D_2_io_r_ofs_0 = _T_419[9:0]; // @[MemPrimitives.scala 131:28:@18909.4]
  assign Mem1D_2_io_r_backpressure = _T_419[10]; // @[MemPrimitives.scala 132:32:@18910.4]
  assign Mem1D_2_io_w_ofs_0 = _T_194[9:0]; // @[MemPrimitives.scala 94:28:@18669.4]
  assign Mem1D_2_io_w_data_0 = _T_194[41:10]; // @[MemPrimitives.scala 95:29:@18670.4]
  assign Mem1D_2_io_w_en_0 = _T_194[42]; // @[MemPrimitives.scala 96:27:@18671.4]
  assign Mem1D_3_clock = clock; // @[:@18493.4]
  assign Mem1D_3_reset = reset; // @[:@18494.4]
  assign Mem1D_3_io_r_ofs_0 = _T_461[9:0]; // @[MemPrimitives.scala 131:28:@18953.4]
  assign Mem1D_3_io_r_backpressure = _T_461[10]; // @[MemPrimitives.scala 132:32:@18954.4]
  assign Mem1D_3_io_w_ofs_0 = _T_205[9:0]; // @[MemPrimitives.scala 94:28:@18681.4]
  assign Mem1D_3_io_w_data_0 = _T_205[41:10]; // @[MemPrimitives.scala 95:29:@18682.4]
  assign Mem1D_3_io_w_en_0 = _T_205[42]; // @[MemPrimitives.scala 96:27:@18683.4]
  assign Mem1D_4_clock = clock; // @[:@18509.4]
  assign Mem1D_4_reset = reset; // @[:@18510.4]
  assign Mem1D_4_io_r_ofs_0 = _T_503[9:0]; // @[MemPrimitives.scala 131:28:@18997.4]
  assign Mem1D_4_io_r_backpressure = _T_503[10]; // @[MemPrimitives.scala 132:32:@18998.4]
  assign Mem1D_4_io_w_ofs_0 = _T_216[9:0]; // @[MemPrimitives.scala 94:28:@18693.4]
  assign Mem1D_4_io_w_data_0 = _T_216[41:10]; // @[MemPrimitives.scala 95:29:@18694.4]
  assign Mem1D_4_io_w_en_0 = _T_216[42]; // @[MemPrimitives.scala 96:27:@18695.4]
  assign Mem1D_5_clock = clock; // @[:@18525.4]
  assign Mem1D_5_reset = reset; // @[:@18526.4]
  assign Mem1D_5_io_r_ofs_0 = _T_545[9:0]; // @[MemPrimitives.scala 131:28:@19041.4]
  assign Mem1D_5_io_r_backpressure = _T_545[10]; // @[MemPrimitives.scala 132:32:@19042.4]
  assign Mem1D_5_io_w_ofs_0 = _T_227[9:0]; // @[MemPrimitives.scala 94:28:@18705.4]
  assign Mem1D_5_io_w_data_0 = _T_227[41:10]; // @[MemPrimitives.scala 95:29:@18706.4]
  assign Mem1D_5_io_w_en_0 = _T_227[42]; // @[MemPrimitives.scala 96:27:@18707.4]
  assign Mem1D_6_clock = clock; // @[:@18541.4]
  assign Mem1D_6_reset = reset; // @[:@18542.4]
  assign Mem1D_6_io_r_ofs_0 = _T_587[9:0]; // @[MemPrimitives.scala 131:28:@19085.4]
  assign Mem1D_6_io_r_backpressure = _T_587[10]; // @[MemPrimitives.scala 132:32:@19086.4]
  assign Mem1D_6_io_w_ofs_0 = _T_238[9:0]; // @[MemPrimitives.scala 94:28:@18717.4]
  assign Mem1D_6_io_w_data_0 = _T_238[41:10]; // @[MemPrimitives.scala 95:29:@18718.4]
  assign Mem1D_6_io_w_en_0 = _T_238[42]; // @[MemPrimitives.scala 96:27:@18719.4]
  assign Mem1D_7_clock = clock; // @[:@18557.4]
  assign Mem1D_7_reset = reset; // @[:@18558.4]
  assign Mem1D_7_io_r_ofs_0 = _T_629[9:0]; // @[MemPrimitives.scala 131:28:@19129.4]
  assign Mem1D_7_io_r_backpressure = _T_629[10]; // @[MemPrimitives.scala 132:32:@19130.4]
  assign Mem1D_7_io_w_ofs_0 = _T_249[9:0]; // @[MemPrimitives.scala 94:28:@18729.4]
  assign Mem1D_7_io_w_data_0 = _T_249[41:10]; // @[MemPrimitives.scala 95:29:@18730.4]
  assign Mem1D_7_io_w_en_0 = _T_249[42]; // @[MemPrimitives.scala 96:27:@18731.4]
  assign Mem1D_8_clock = clock; // @[:@18573.4]
  assign Mem1D_8_reset = reset; // @[:@18574.4]
  assign Mem1D_8_io_r_ofs_0 = _T_671[9:0]; // @[MemPrimitives.scala 131:28:@19173.4]
  assign Mem1D_8_io_r_backpressure = _T_671[10]; // @[MemPrimitives.scala 132:32:@19174.4]
  assign Mem1D_8_io_w_ofs_0 = _T_260[9:0]; // @[MemPrimitives.scala 94:28:@18741.4]
  assign Mem1D_8_io_w_data_0 = _T_260[41:10]; // @[MemPrimitives.scala 95:29:@18742.4]
  assign Mem1D_8_io_w_en_0 = _T_260[42]; // @[MemPrimitives.scala 96:27:@18743.4]
  assign Mem1D_9_clock = clock; // @[:@18589.4]
  assign Mem1D_9_reset = reset; // @[:@18590.4]
  assign Mem1D_9_io_r_ofs_0 = _T_713[9:0]; // @[MemPrimitives.scala 131:28:@19217.4]
  assign Mem1D_9_io_r_backpressure = _T_713[10]; // @[MemPrimitives.scala 132:32:@19218.4]
  assign Mem1D_9_io_w_ofs_0 = _T_271[9:0]; // @[MemPrimitives.scala 94:28:@18753.4]
  assign Mem1D_9_io_w_data_0 = _T_271[41:10]; // @[MemPrimitives.scala 95:29:@18754.4]
  assign Mem1D_9_io_w_en_0 = _T_271[42]; // @[MemPrimitives.scala 96:27:@18755.4]
  assign Mem1D_10_clock = clock; // @[:@18605.4]
  assign Mem1D_10_reset = reset; // @[:@18606.4]
  assign Mem1D_10_io_r_ofs_0 = _T_755[9:0]; // @[MemPrimitives.scala 131:28:@19261.4]
  assign Mem1D_10_io_r_backpressure = _T_755[10]; // @[MemPrimitives.scala 132:32:@19262.4]
  assign Mem1D_10_io_w_ofs_0 = _T_282[9:0]; // @[MemPrimitives.scala 94:28:@18765.4]
  assign Mem1D_10_io_w_data_0 = _T_282[41:10]; // @[MemPrimitives.scala 95:29:@18766.4]
  assign Mem1D_10_io_w_en_0 = _T_282[42]; // @[MemPrimitives.scala 96:27:@18767.4]
  assign Mem1D_11_clock = clock; // @[:@18621.4]
  assign Mem1D_11_reset = reset; // @[:@18622.4]
  assign Mem1D_11_io_r_ofs_0 = _T_797[9:0]; // @[MemPrimitives.scala 131:28:@19305.4]
  assign Mem1D_11_io_r_backpressure = _T_797[10]; // @[MemPrimitives.scala 132:32:@19306.4]
  assign Mem1D_11_io_w_ofs_0 = _T_293[9:0]; // @[MemPrimitives.scala 94:28:@18777.4]
  assign Mem1D_11_io_w_data_0 = _T_293[41:10]; // @[MemPrimitives.scala 95:29:@18778.4]
  assign Mem1D_11_io_w_en_0 = _T_293[42]; // @[MemPrimitives.scala 96:27:@18779.4]
  assign StickySelects_clock = clock; // @[:@18797.4]
  assign StickySelects_reset = reset; // @[:@18798.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_301; // @[MemPrimitives.scala 125:64:@18799.4]
  assign StickySelects_io_ins_1 = io_rPort_1_en_0 & _T_307; // @[MemPrimitives.scala 125:64:@18800.4]
  assign StickySelects_io_ins_2 = io_rPort_2_en_0 & _T_313; // @[MemPrimitives.scala 125:64:@18801.4]
  assign StickySelects_io_ins_3 = io_rPort_3_en_0 & _T_319; // @[MemPrimitives.scala 125:64:@18802.4]
  assign StickySelects_1_clock = clock; // @[:@18841.4]
  assign StickySelects_1_reset = reset; // @[:@18842.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_343; // @[MemPrimitives.scala 125:64:@18843.4]
  assign StickySelects_1_io_ins_1 = io_rPort_1_en_0 & _T_349; // @[MemPrimitives.scala 125:64:@18844.4]
  assign StickySelects_1_io_ins_2 = io_rPort_2_en_0 & _T_355; // @[MemPrimitives.scala 125:64:@18845.4]
  assign StickySelects_1_io_ins_3 = io_rPort_3_en_0 & _T_361; // @[MemPrimitives.scala 125:64:@18846.4]
  assign StickySelects_2_clock = clock; // @[:@18885.4]
  assign StickySelects_2_reset = reset; // @[:@18886.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_385; // @[MemPrimitives.scala 125:64:@18887.4]
  assign StickySelects_2_io_ins_1 = io_rPort_1_en_0 & _T_391; // @[MemPrimitives.scala 125:64:@18888.4]
  assign StickySelects_2_io_ins_2 = io_rPort_2_en_0 & _T_397; // @[MemPrimitives.scala 125:64:@18889.4]
  assign StickySelects_2_io_ins_3 = io_rPort_3_en_0 & _T_403; // @[MemPrimitives.scala 125:64:@18890.4]
  assign StickySelects_3_clock = clock; // @[:@18929.4]
  assign StickySelects_3_reset = reset; // @[:@18930.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_427; // @[MemPrimitives.scala 125:64:@18931.4]
  assign StickySelects_3_io_ins_1 = io_rPort_1_en_0 & _T_433; // @[MemPrimitives.scala 125:64:@18932.4]
  assign StickySelects_3_io_ins_2 = io_rPort_2_en_0 & _T_439; // @[MemPrimitives.scala 125:64:@18933.4]
  assign StickySelects_3_io_ins_3 = io_rPort_3_en_0 & _T_445; // @[MemPrimitives.scala 125:64:@18934.4]
  assign StickySelects_4_clock = clock; // @[:@18973.4]
  assign StickySelects_4_reset = reset; // @[:@18974.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_469; // @[MemPrimitives.scala 125:64:@18975.4]
  assign StickySelects_4_io_ins_1 = io_rPort_1_en_0 & _T_475; // @[MemPrimitives.scala 125:64:@18976.4]
  assign StickySelects_4_io_ins_2 = io_rPort_2_en_0 & _T_481; // @[MemPrimitives.scala 125:64:@18977.4]
  assign StickySelects_4_io_ins_3 = io_rPort_3_en_0 & _T_487; // @[MemPrimitives.scala 125:64:@18978.4]
  assign StickySelects_5_clock = clock; // @[:@19017.4]
  assign StickySelects_5_reset = reset; // @[:@19018.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_511; // @[MemPrimitives.scala 125:64:@19019.4]
  assign StickySelects_5_io_ins_1 = io_rPort_1_en_0 & _T_517; // @[MemPrimitives.scala 125:64:@19020.4]
  assign StickySelects_5_io_ins_2 = io_rPort_2_en_0 & _T_523; // @[MemPrimitives.scala 125:64:@19021.4]
  assign StickySelects_5_io_ins_3 = io_rPort_3_en_0 & _T_529; // @[MemPrimitives.scala 125:64:@19022.4]
  assign StickySelects_6_clock = clock; // @[:@19061.4]
  assign StickySelects_6_reset = reset; // @[:@19062.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_553; // @[MemPrimitives.scala 125:64:@19063.4]
  assign StickySelects_6_io_ins_1 = io_rPort_1_en_0 & _T_559; // @[MemPrimitives.scala 125:64:@19064.4]
  assign StickySelects_6_io_ins_2 = io_rPort_2_en_0 & _T_565; // @[MemPrimitives.scala 125:64:@19065.4]
  assign StickySelects_6_io_ins_3 = io_rPort_3_en_0 & _T_571; // @[MemPrimitives.scala 125:64:@19066.4]
  assign StickySelects_7_clock = clock; // @[:@19105.4]
  assign StickySelects_7_reset = reset; // @[:@19106.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_595; // @[MemPrimitives.scala 125:64:@19107.4]
  assign StickySelects_7_io_ins_1 = io_rPort_1_en_0 & _T_601; // @[MemPrimitives.scala 125:64:@19108.4]
  assign StickySelects_7_io_ins_2 = io_rPort_2_en_0 & _T_607; // @[MemPrimitives.scala 125:64:@19109.4]
  assign StickySelects_7_io_ins_3 = io_rPort_3_en_0 & _T_613; // @[MemPrimitives.scala 125:64:@19110.4]
  assign StickySelects_8_clock = clock; // @[:@19149.4]
  assign StickySelects_8_reset = reset; // @[:@19150.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_637; // @[MemPrimitives.scala 125:64:@19151.4]
  assign StickySelects_8_io_ins_1 = io_rPort_1_en_0 & _T_643; // @[MemPrimitives.scala 125:64:@19152.4]
  assign StickySelects_8_io_ins_2 = io_rPort_2_en_0 & _T_649; // @[MemPrimitives.scala 125:64:@19153.4]
  assign StickySelects_8_io_ins_3 = io_rPort_3_en_0 & _T_655; // @[MemPrimitives.scala 125:64:@19154.4]
  assign StickySelects_9_clock = clock; // @[:@19193.4]
  assign StickySelects_9_reset = reset; // @[:@19194.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_679; // @[MemPrimitives.scala 125:64:@19195.4]
  assign StickySelects_9_io_ins_1 = io_rPort_1_en_0 & _T_685; // @[MemPrimitives.scala 125:64:@19196.4]
  assign StickySelects_9_io_ins_2 = io_rPort_2_en_0 & _T_691; // @[MemPrimitives.scala 125:64:@19197.4]
  assign StickySelects_9_io_ins_3 = io_rPort_3_en_0 & _T_697; // @[MemPrimitives.scala 125:64:@19198.4]
  assign StickySelects_10_clock = clock; // @[:@19237.4]
  assign StickySelects_10_reset = reset; // @[:@19238.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_721; // @[MemPrimitives.scala 125:64:@19239.4]
  assign StickySelects_10_io_ins_1 = io_rPort_1_en_0 & _T_727; // @[MemPrimitives.scala 125:64:@19240.4]
  assign StickySelects_10_io_ins_2 = io_rPort_2_en_0 & _T_733; // @[MemPrimitives.scala 125:64:@19241.4]
  assign StickySelects_10_io_ins_3 = io_rPort_3_en_0 & _T_739; // @[MemPrimitives.scala 125:64:@19242.4]
  assign StickySelects_11_clock = clock; // @[:@19281.4]
  assign StickySelects_11_reset = reset; // @[:@19282.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_763; // @[MemPrimitives.scala 125:64:@19283.4]
  assign StickySelects_11_io_ins_1 = io_rPort_1_en_0 & _T_769; // @[MemPrimitives.scala 125:64:@19284.4]
  assign StickySelects_11_io_ins_2 = io_rPort_2_en_0 & _T_775; // @[MemPrimitives.scala 125:64:@19285.4]
  assign StickySelects_11_io_ins_3 = io_rPort_3_en_0 & _T_781; // @[MemPrimitives.scala 125:64:@19286.4]
  assign RetimeWrapper_clock = clock; // @[:@19346.4]
  assign RetimeWrapper_reset = reset; // @[:@19347.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19349.4]
  assign RetimeWrapper_io_in = _T_301 & io_rPort_0_en_0; // @[package.scala 94:16:@19348.4]
  assign RetimeWrapper_1_clock = clock; // @[:@19354.4]
  assign RetimeWrapper_1_reset = reset; // @[:@19355.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19357.4]
  assign RetimeWrapper_1_io_in = _T_343 & io_rPort_0_en_0; // @[package.scala 94:16:@19356.4]
  assign RetimeWrapper_2_clock = clock; // @[:@19362.4]
  assign RetimeWrapper_2_reset = reset; // @[:@19363.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19365.4]
  assign RetimeWrapper_2_io_in = _T_385 & io_rPort_0_en_0; // @[package.scala 94:16:@19364.4]
  assign RetimeWrapper_3_clock = clock; // @[:@19370.4]
  assign RetimeWrapper_3_reset = reset; // @[:@19371.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19373.4]
  assign RetimeWrapper_3_io_in = _T_427 & io_rPort_0_en_0; // @[package.scala 94:16:@19372.4]
  assign RetimeWrapper_4_clock = clock; // @[:@19378.4]
  assign RetimeWrapper_4_reset = reset; // @[:@19379.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19381.4]
  assign RetimeWrapper_4_io_in = _T_469 & io_rPort_0_en_0; // @[package.scala 94:16:@19380.4]
  assign RetimeWrapper_5_clock = clock; // @[:@19386.4]
  assign RetimeWrapper_5_reset = reset; // @[:@19387.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19389.4]
  assign RetimeWrapper_5_io_in = _T_511 & io_rPort_0_en_0; // @[package.scala 94:16:@19388.4]
  assign RetimeWrapper_6_clock = clock; // @[:@19394.4]
  assign RetimeWrapper_6_reset = reset; // @[:@19395.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19397.4]
  assign RetimeWrapper_6_io_in = _T_553 & io_rPort_0_en_0; // @[package.scala 94:16:@19396.4]
  assign RetimeWrapper_7_clock = clock; // @[:@19402.4]
  assign RetimeWrapper_7_reset = reset; // @[:@19403.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19405.4]
  assign RetimeWrapper_7_io_in = _T_595 & io_rPort_0_en_0; // @[package.scala 94:16:@19404.4]
  assign RetimeWrapper_8_clock = clock; // @[:@19410.4]
  assign RetimeWrapper_8_reset = reset; // @[:@19411.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19413.4]
  assign RetimeWrapper_8_io_in = _T_637 & io_rPort_0_en_0; // @[package.scala 94:16:@19412.4]
  assign RetimeWrapper_9_clock = clock; // @[:@19418.4]
  assign RetimeWrapper_9_reset = reset; // @[:@19419.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19421.4]
  assign RetimeWrapper_9_io_in = _T_679 & io_rPort_0_en_0; // @[package.scala 94:16:@19420.4]
  assign RetimeWrapper_10_clock = clock; // @[:@19426.4]
  assign RetimeWrapper_10_reset = reset; // @[:@19427.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19429.4]
  assign RetimeWrapper_10_io_in = _T_721 & io_rPort_0_en_0; // @[package.scala 94:16:@19428.4]
  assign RetimeWrapper_11_clock = clock; // @[:@19434.4]
  assign RetimeWrapper_11_reset = reset; // @[:@19435.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19437.4]
  assign RetimeWrapper_11_io_in = _T_763 & io_rPort_0_en_0; // @[package.scala 94:16:@19436.4]
  assign RetimeWrapper_12_clock = clock; // @[:@19490.4]
  assign RetimeWrapper_12_reset = reset; // @[:@19491.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19493.4]
  assign RetimeWrapper_12_io_in = _T_307 & io_rPort_1_en_0; // @[package.scala 94:16:@19492.4]
  assign RetimeWrapper_13_clock = clock; // @[:@19498.4]
  assign RetimeWrapper_13_reset = reset; // @[:@19499.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19501.4]
  assign RetimeWrapper_13_io_in = _T_349 & io_rPort_1_en_0; // @[package.scala 94:16:@19500.4]
  assign RetimeWrapper_14_clock = clock; // @[:@19506.4]
  assign RetimeWrapper_14_reset = reset; // @[:@19507.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19509.4]
  assign RetimeWrapper_14_io_in = _T_391 & io_rPort_1_en_0; // @[package.scala 94:16:@19508.4]
  assign RetimeWrapper_15_clock = clock; // @[:@19514.4]
  assign RetimeWrapper_15_reset = reset; // @[:@19515.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19517.4]
  assign RetimeWrapper_15_io_in = _T_433 & io_rPort_1_en_0; // @[package.scala 94:16:@19516.4]
  assign RetimeWrapper_16_clock = clock; // @[:@19522.4]
  assign RetimeWrapper_16_reset = reset; // @[:@19523.4]
  assign RetimeWrapper_16_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19525.4]
  assign RetimeWrapper_16_io_in = _T_475 & io_rPort_1_en_0; // @[package.scala 94:16:@19524.4]
  assign RetimeWrapper_17_clock = clock; // @[:@19530.4]
  assign RetimeWrapper_17_reset = reset; // @[:@19531.4]
  assign RetimeWrapper_17_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19533.4]
  assign RetimeWrapper_17_io_in = _T_517 & io_rPort_1_en_0; // @[package.scala 94:16:@19532.4]
  assign RetimeWrapper_18_clock = clock; // @[:@19538.4]
  assign RetimeWrapper_18_reset = reset; // @[:@19539.4]
  assign RetimeWrapper_18_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19541.4]
  assign RetimeWrapper_18_io_in = _T_559 & io_rPort_1_en_0; // @[package.scala 94:16:@19540.4]
  assign RetimeWrapper_19_clock = clock; // @[:@19546.4]
  assign RetimeWrapper_19_reset = reset; // @[:@19547.4]
  assign RetimeWrapper_19_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19549.4]
  assign RetimeWrapper_19_io_in = _T_601 & io_rPort_1_en_0; // @[package.scala 94:16:@19548.4]
  assign RetimeWrapper_20_clock = clock; // @[:@19554.4]
  assign RetimeWrapper_20_reset = reset; // @[:@19555.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19557.4]
  assign RetimeWrapper_20_io_in = _T_643 & io_rPort_1_en_0; // @[package.scala 94:16:@19556.4]
  assign RetimeWrapper_21_clock = clock; // @[:@19562.4]
  assign RetimeWrapper_21_reset = reset; // @[:@19563.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19565.4]
  assign RetimeWrapper_21_io_in = _T_685 & io_rPort_1_en_0; // @[package.scala 94:16:@19564.4]
  assign RetimeWrapper_22_clock = clock; // @[:@19570.4]
  assign RetimeWrapper_22_reset = reset; // @[:@19571.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19573.4]
  assign RetimeWrapper_22_io_in = _T_727 & io_rPort_1_en_0; // @[package.scala 94:16:@19572.4]
  assign RetimeWrapper_23_clock = clock; // @[:@19578.4]
  assign RetimeWrapper_23_reset = reset; // @[:@19579.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19581.4]
  assign RetimeWrapper_23_io_in = _T_769 & io_rPort_1_en_0; // @[package.scala 94:16:@19580.4]
  assign RetimeWrapper_24_clock = clock; // @[:@19634.4]
  assign RetimeWrapper_24_reset = reset; // @[:@19635.4]
  assign RetimeWrapper_24_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19637.4]
  assign RetimeWrapper_24_io_in = _T_313 & io_rPort_2_en_0; // @[package.scala 94:16:@19636.4]
  assign RetimeWrapper_25_clock = clock; // @[:@19642.4]
  assign RetimeWrapper_25_reset = reset; // @[:@19643.4]
  assign RetimeWrapper_25_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19645.4]
  assign RetimeWrapper_25_io_in = _T_355 & io_rPort_2_en_0; // @[package.scala 94:16:@19644.4]
  assign RetimeWrapper_26_clock = clock; // @[:@19650.4]
  assign RetimeWrapper_26_reset = reset; // @[:@19651.4]
  assign RetimeWrapper_26_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19653.4]
  assign RetimeWrapper_26_io_in = _T_397 & io_rPort_2_en_0; // @[package.scala 94:16:@19652.4]
  assign RetimeWrapper_27_clock = clock; // @[:@19658.4]
  assign RetimeWrapper_27_reset = reset; // @[:@19659.4]
  assign RetimeWrapper_27_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19661.4]
  assign RetimeWrapper_27_io_in = _T_439 & io_rPort_2_en_0; // @[package.scala 94:16:@19660.4]
  assign RetimeWrapper_28_clock = clock; // @[:@19666.4]
  assign RetimeWrapper_28_reset = reset; // @[:@19667.4]
  assign RetimeWrapper_28_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19669.4]
  assign RetimeWrapper_28_io_in = _T_481 & io_rPort_2_en_0; // @[package.scala 94:16:@19668.4]
  assign RetimeWrapper_29_clock = clock; // @[:@19674.4]
  assign RetimeWrapper_29_reset = reset; // @[:@19675.4]
  assign RetimeWrapper_29_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19677.4]
  assign RetimeWrapper_29_io_in = _T_523 & io_rPort_2_en_0; // @[package.scala 94:16:@19676.4]
  assign RetimeWrapper_30_clock = clock; // @[:@19682.4]
  assign RetimeWrapper_30_reset = reset; // @[:@19683.4]
  assign RetimeWrapper_30_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19685.4]
  assign RetimeWrapper_30_io_in = _T_565 & io_rPort_2_en_0; // @[package.scala 94:16:@19684.4]
  assign RetimeWrapper_31_clock = clock; // @[:@19690.4]
  assign RetimeWrapper_31_reset = reset; // @[:@19691.4]
  assign RetimeWrapper_31_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19693.4]
  assign RetimeWrapper_31_io_in = _T_607 & io_rPort_2_en_0; // @[package.scala 94:16:@19692.4]
  assign RetimeWrapper_32_clock = clock; // @[:@19698.4]
  assign RetimeWrapper_32_reset = reset; // @[:@19699.4]
  assign RetimeWrapper_32_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19701.4]
  assign RetimeWrapper_32_io_in = _T_649 & io_rPort_2_en_0; // @[package.scala 94:16:@19700.4]
  assign RetimeWrapper_33_clock = clock; // @[:@19706.4]
  assign RetimeWrapper_33_reset = reset; // @[:@19707.4]
  assign RetimeWrapper_33_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19709.4]
  assign RetimeWrapper_33_io_in = _T_691 & io_rPort_2_en_0; // @[package.scala 94:16:@19708.4]
  assign RetimeWrapper_34_clock = clock; // @[:@19714.4]
  assign RetimeWrapper_34_reset = reset; // @[:@19715.4]
  assign RetimeWrapper_34_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19717.4]
  assign RetimeWrapper_34_io_in = _T_733 & io_rPort_2_en_0; // @[package.scala 94:16:@19716.4]
  assign RetimeWrapper_35_clock = clock; // @[:@19722.4]
  assign RetimeWrapper_35_reset = reset; // @[:@19723.4]
  assign RetimeWrapper_35_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19725.4]
  assign RetimeWrapper_35_io_in = _T_775 & io_rPort_2_en_0; // @[package.scala 94:16:@19724.4]
  assign RetimeWrapper_36_clock = clock; // @[:@19778.4]
  assign RetimeWrapper_36_reset = reset; // @[:@19779.4]
  assign RetimeWrapper_36_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19781.4]
  assign RetimeWrapper_36_io_in = _T_319 & io_rPort_3_en_0; // @[package.scala 94:16:@19780.4]
  assign RetimeWrapper_37_clock = clock; // @[:@19786.4]
  assign RetimeWrapper_37_reset = reset; // @[:@19787.4]
  assign RetimeWrapper_37_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19789.4]
  assign RetimeWrapper_37_io_in = _T_361 & io_rPort_3_en_0; // @[package.scala 94:16:@19788.4]
  assign RetimeWrapper_38_clock = clock; // @[:@19794.4]
  assign RetimeWrapper_38_reset = reset; // @[:@19795.4]
  assign RetimeWrapper_38_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19797.4]
  assign RetimeWrapper_38_io_in = _T_403 & io_rPort_3_en_0; // @[package.scala 94:16:@19796.4]
  assign RetimeWrapper_39_clock = clock; // @[:@19802.4]
  assign RetimeWrapper_39_reset = reset; // @[:@19803.4]
  assign RetimeWrapper_39_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19805.4]
  assign RetimeWrapper_39_io_in = _T_445 & io_rPort_3_en_0; // @[package.scala 94:16:@19804.4]
  assign RetimeWrapper_40_clock = clock; // @[:@19810.4]
  assign RetimeWrapper_40_reset = reset; // @[:@19811.4]
  assign RetimeWrapper_40_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19813.4]
  assign RetimeWrapper_40_io_in = _T_487 & io_rPort_3_en_0; // @[package.scala 94:16:@19812.4]
  assign RetimeWrapper_41_clock = clock; // @[:@19818.4]
  assign RetimeWrapper_41_reset = reset; // @[:@19819.4]
  assign RetimeWrapper_41_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19821.4]
  assign RetimeWrapper_41_io_in = _T_529 & io_rPort_3_en_0; // @[package.scala 94:16:@19820.4]
  assign RetimeWrapper_42_clock = clock; // @[:@19826.4]
  assign RetimeWrapper_42_reset = reset; // @[:@19827.4]
  assign RetimeWrapper_42_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19829.4]
  assign RetimeWrapper_42_io_in = _T_571 & io_rPort_3_en_0; // @[package.scala 94:16:@19828.4]
  assign RetimeWrapper_43_clock = clock; // @[:@19834.4]
  assign RetimeWrapper_43_reset = reset; // @[:@19835.4]
  assign RetimeWrapper_43_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19837.4]
  assign RetimeWrapper_43_io_in = _T_613 & io_rPort_3_en_0; // @[package.scala 94:16:@19836.4]
  assign RetimeWrapper_44_clock = clock; // @[:@19842.4]
  assign RetimeWrapper_44_reset = reset; // @[:@19843.4]
  assign RetimeWrapper_44_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19845.4]
  assign RetimeWrapper_44_io_in = _T_655 & io_rPort_3_en_0; // @[package.scala 94:16:@19844.4]
  assign RetimeWrapper_45_clock = clock; // @[:@19850.4]
  assign RetimeWrapper_45_reset = reset; // @[:@19851.4]
  assign RetimeWrapper_45_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19853.4]
  assign RetimeWrapper_45_io_in = _T_697 & io_rPort_3_en_0; // @[package.scala 94:16:@19852.4]
  assign RetimeWrapper_46_clock = clock; // @[:@19858.4]
  assign RetimeWrapper_46_reset = reset; // @[:@19859.4]
  assign RetimeWrapper_46_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19861.4]
  assign RetimeWrapper_46_io_in = _T_739 & io_rPort_3_en_0; // @[package.scala 94:16:@19860.4]
  assign RetimeWrapper_47_clock = clock; // @[:@19866.4]
  assign RetimeWrapper_47_reset = reset; // @[:@19867.4]
  assign RetimeWrapper_47_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19869.4]
  assign RetimeWrapper_47_io_in = _T_781 & io_rPort_3_en_0; // @[package.scala 94:16:@19868.4]
endmodule
module Divider( // @[:@21491.2]
  input         clock, // @[:@21492.4]
  input         io_flow, // @[:@21494.4]
  input  [31:0] io_dividend, // @[:@21494.4]
  input  [31:0] io_divisor, // @[:@21494.4]
  output [31:0] io_out // @[:@21494.4]
);
  wire [31:0] m_m_axis_dout_tdata; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire  m_m_axis_dout_tvalid; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire [31:0] m_s_axis_divisor_tdata; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire  m_s_axis_divisor_tvalid; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire [31:0] m_s_axis_dividend_tdata; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire  m_s_axis_dividend_tvalid; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire  m_aclken; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire  m_aclk; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire [29:0] _T_15; // @[ZynqBlackBoxes.scala 34:37:@21512.4]
  div_32_32_20_Signed_Fractional m ( // @[ZynqBlackBoxes.scala 26:19:@21496.4]
    .m_axis_dout_tdata(m_m_axis_dout_tdata),
    .m_axis_dout_tvalid(m_m_axis_dout_tvalid),
    .s_axis_divisor_tdata(m_s_axis_divisor_tdata),
    .s_axis_divisor_tvalid(m_s_axis_divisor_tvalid),
    .s_axis_dividend_tdata(m_s_axis_dividend_tdata),
    .s_axis_dividend_tvalid(m_s_axis_dividend_tvalid),
    .aclken(m_aclken),
    .aclk(m_aclk)
  );
  assign _T_15 = m_m_axis_dout_tdata[31:2]; // @[ZynqBlackBoxes.scala 34:37:@21512.4]
  assign io_out = {{2'd0}, _T_15}; // @[ZynqBlackBoxes.scala 34:12:@21513.4]
  assign m_s_axis_divisor_tdata = io_divisor; // @[ZynqBlackBoxes.scala 32:31:@21510.4]
  assign m_s_axis_divisor_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 31:32:@21509.4]
  assign m_s_axis_dividend_tdata = io_dividend; // @[ZynqBlackBoxes.scala 30:32:@21508.4]
  assign m_s_axis_dividend_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 29:33:@21507.4]
  assign m_aclken = io_flow; // @[ZynqBlackBoxes.scala 28:17:@21506.4 ZynqBlackBoxes.scala 33:17:@21511.4]
  assign m_aclk = clock; // @[ZynqBlackBoxes.scala 27:15:@21505.4]
endmodule
module x250_div( // @[:@21551.2]
  input         clock, // @[:@21552.4]
  input  [31:0] io_a, // @[:@21554.4]
  input         io_flow, // @[:@21554.4]
  output [31:0] io_result // @[:@21554.4]
);
  wire  x250_div_clock; // @[BigIPZynq.scala 25:21:@21562.4]
  wire  x250_div_io_flow; // @[BigIPZynq.scala 25:21:@21562.4]
  wire [31:0] x250_div_io_dividend; // @[BigIPZynq.scala 25:21:@21562.4]
  wire [31:0] x250_div_io_divisor; // @[BigIPZynq.scala 25:21:@21562.4]
  wire [31:0] x250_div_io_out; // @[BigIPZynq.scala 25:21:@21562.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@21575.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@21575.4]
  wire [31:0] _T_15; // @[FixedPoint.scala 24:59:@21560.4]
  wire [31:0] _T_19; // @[BigIPZynq.scala 29:16:@21570.4]
  Divider x250_div ( // @[BigIPZynq.scala 25:21:@21562.4]
    .clock(x250_div_clock),
    .io_flow(x250_div_io_flow),
    .io_dividend(x250_div_io_dividend),
    .io_divisor(x250_div_io_divisor),
    .io_out(x250_div_io_out)
  );
  _ _ ( // @[Math.scala 720:24:@21575.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign _T_15 = $signed(io_a); // @[FixedPoint.scala 24:59:@21560.4]
  assign _T_19 = $signed(x250_div_io_out); // @[BigIPZynq.scala 29:16:@21570.4]
  assign io_result = __io_result; // @[Math.scala 290:34:@21583.4]
  assign x250_div_clock = clock; // @[:@21563.4]
  assign x250_div_io_flow = io_flow; // @[BigIPZynq.scala 28:17:@21569.4]
  assign x250_div_io_dividend = $unsigned(_T_15); // @[BigIPZynq.scala 26:21:@21566.4]
  assign x250_div_io_divisor = 32'h3; // @[BigIPZynq.scala 27:20:@21568.4]
  assign __io_b = $unsigned(_T_19); // @[Math.scala 721:17:@21578.4]
endmodule
module RetimeWrapper_243( // @[:@21597.2]
  input         clock, // @[:@21598.4]
  input         reset, // @[:@21599.4]
  input         io_flow, // @[:@21600.4]
  input  [31:0] io_in, // @[:@21600.4]
  output [31:0] io_out // @[:@21600.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21602.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21602.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21602.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21602.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21602.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21602.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(19)) sr ( // @[RetimeShiftRegister.scala 15:20:@21602.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21615.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21614.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21613.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21612.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21611.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21609.4]
endmodule
module RetimeWrapper_245( // @[:@21808.2]
  input   clock, // @[:@21809.4]
  input   reset, // @[:@21810.4]
  input   io_flow, // @[:@21811.4]
  input   io_in, // @[:@21811.4]
  output  io_out // @[:@21811.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@21813.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@21813.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@21813.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21813.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21813.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21813.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@21813.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21826.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21825.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@21824.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21823.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21822.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21820.4]
endmodule
module RetimeWrapper_246( // @[:@21840.2]
  input         clock, // @[:@21841.4]
  input         reset, // @[:@21842.4]
  input         io_flow, // @[:@21843.4]
  input  [31:0] io_in, // @[:@21843.4]
  output [31:0] io_out // @[:@21843.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21845.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21845.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21845.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21845.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21845.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21845.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(13)) sr ( // @[RetimeShiftRegister.scala 15:20:@21845.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21858.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21857.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21856.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21855.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21854.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21852.4]
endmodule
module RetimeWrapper_248( // @[:@21904.2]
  input         clock, // @[:@21905.4]
  input         reset, // @[:@21906.4]
  input         io_flow, // @[:@21907.4]
  input  [31:0] io_in, // @[:@21907.4]
  output [31:0] io_out // @[:@21907.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21909.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21909.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21909.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21909.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21909.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21909.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@21909.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21922.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21921.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21920.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21919.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21918.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21916.4]
endmodule
module RetimeWrapper_249( // @[:@21936.2]
  input         clock, // @[:@21937.4]
  input         reset, // @[:@21938.4]
  input         io_flow, // @[:@21939.4]
  input  [31:0] io_in, // @[:@21939.4]
  output [31:0] io_out // @[:@21939.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21941.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21941.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21941.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21941.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21941.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21941.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@21941.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21954.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21953.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21952.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21951.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21950.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21948.4]
endmodule
module RetimeWrapper_251( // @[:@22000.2]
  input         clock, // @[:@22001.4]
  input         reset, // @[:@22002.4]
  input         io_flow, // @[:@22003.4]
  input  [31:0] io_in, // @[:@22003.4]
  output [31:0] io_out // @[:@22003.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22005.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22005.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22005.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22005.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22005.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22005.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@22005.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22018.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22017.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22016.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22015.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22014.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22012.4]
endmodule
module RetimeWrapper_256( // @[:@22160.2]
  input   clock, // @[:@22161.4]
  input   reset, // @[:@22162.4]
  input   io_flow, // @[:@22163.4]
  input   io_in, // @[:@22163.4]
  output  io_out // @[:@22163.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@22165.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@22165.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@22165.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22165.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22165.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22165.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(45)) sr ( // @[RetimeShiftRegister.scala 15:20:@22165.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22178.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22177.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@22176.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22175.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22174.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22172.4]
endmodule
module RetimeWrapper_257( // @[:@22192.2]
  input         clock, // @[:@22193.4]
  input         reset, // @[:@22194.4]
  input         io_flow, // @[:@22195.4]
  input  [31:0] io_in, // @[:@22195.4]
  output [31:0] io_out // @[:@22195.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22197.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22197.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22197.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22197.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22197.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22197.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(37)) sr ( // @[RetimeShiftRegister.scala 15:20:@22197.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22210.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22209.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22208.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22207.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22206.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22204.4]
endmodule
module RetimeWrapper_259( // @[:@22256.2]
  input         clock, // @[:@22257.4]
  input         reset, // @[:@22258.4]
  input         io_flow, // @[:@22259.4]
  input  [31:0] io_in, // @[:@22259.4]
  output [31:0] io_out // @[:@22259.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22261.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22261.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22261.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22261.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22261.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22261.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(45)) sr ( // @[RetimeShiftRegister.scala 15:20:@22261.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22274.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22273.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22272.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22271.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22270.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22268.4]
endmodule
module RetimeWrapper_260( // @[:@22288.2]
  input         clock, // @[:@22289.4]
  input         reset, // @[:@22290.4]
  input         io_flow, // @[:@22291.4]
  input  [31:0] io_in, // @[:@22291.4]
  output [31:0] io_out // @[:@22291.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22293.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22293.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22293.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22293.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22293.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22293.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@22293.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22306.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22305.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22304.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22303.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22302.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22300.4]
endmodule
module RetimeWrapper_277( // @[:@24117.2]
  input         clock, // @[:@24118.4]
  input         reset, // @[:@24119.4]
  input         io_flow, // @[:@24120.4]
  input  [31:0] io_in, // @[:@24120.4]
  output [31:0] io_out // @[:@24120.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@24122.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@24122.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@24122.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24122.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24122.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24122.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(43)) sr ( // @[RetimeShiftRegister.scala 15:20:@24122.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24135.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24134.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@24133.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24132.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24131.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24129.4]
endmodule
module RetimeWrapper_280( // @[:@24360.2]
  input   clock, // @[:@24361.4]
  input   reset, // @[:@24362.4]
  input   io_flow, // @[:@24363.4]
  input   io_in, // @[:@24363.4]
  output  io_out // @[:@24363.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@24365.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@24365.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@24365.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24365.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24365.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24365.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@24365.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24378.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24377.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@24376.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24375.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24374.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24372.4]
endmodule
module RetimeWrapper_307( // @[:@26951.2]
  input         clock, // @[:@26952.4]
  input         reset, // @[:@26953.4]
  input         io_flow, // @[:@26954.4]
  input  [31:0] io_in, // @[:@26954.4]
  output [31:0] io_out // @[:@26954.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26956.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26956.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26956.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26956.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26956.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26956.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(17)) sr ( // @[RetimeShiftRegister.scala 15:20:@26956.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26969.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26968.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26967.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26966.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26965.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26963.4]
endmodule
module RetimeWrapper_313( // @[:@27290.2]
  input         clock, // @[:@27291.4]
  input         reset, // @[:@27292.4]
  input         io_flow, // @[:@27293.4]
  input  [31:0] io_in, // @[:@27293.4]
  output [31:0] io_out // @[:@27293.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@27295.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@27295.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@27295.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@27295.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@27295.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@27295.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@27295.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@27308.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@27307.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@27306.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@27305.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@27304.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@27302.4]
endmodule
module fix2fixBox_128( // @[:@29108.2]
  input  [31:0] io_a, // @[:@29111.4]
  output [32:0] io_b // @[:@29111.4]
);
  assign io_b = {1'h0,io_a}; // @[Converter.scala 95:38:@29125.4]
endmodule
module __87( // @[:@29127.2]
  input  [31:0] io_b, // @[:@29130.4]
  output [32:0] io_result // @[:@29130.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@29135.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@29135.4]
  fix2fixBox_128 fix2fixBox ( // @[BigIPZynq.scala 219:30:@29135.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@29143.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@29138.4]
endmodule
module x325_x7( // @[:@29239.2]
  input         clock, // @[:@29240.4]
  input         reset, // @[:@29241.4]
  input  [31:0] io_a, // @[:@29242.4]
  input  [31:0] io_b, // @[:@29242.4]
  input         io_flow, // @[:@29242.4]
  output [31:0] io_result // @[:@29242.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@29250.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@29250.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@29257.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@29257.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@29267.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@29267.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@29267.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@29267.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@29267.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@29255.4 Math.scala 724:14:@29256.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@29262.4 Math.scala 724:14:@29263.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@29264.4]
  __87 _ ( // @[Math.scala 720:24:@29250.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __87 __1 ( // @[Math.scala 720:24:@29257.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@29267.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@29255.4 Math.scala 724:14:@29256.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@29262.4 Math.scala 724:14:@29263.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@29264.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@29275.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@29253.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@29260.4]
  assign fix2fixBox_clock = clock; // @[:@29268.4]
  assign fix2fixBox_reset = reset; // @[:@29269.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@29270.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@29273.4]
endmodule
module RetimeWrapper_345( // @[:@30303.2]
  input         clock, // @[:@30304.4]
  input         reset, // @[:@30305.4]
  input         io_flow, // @[:@30306.4]
  input  [31:0] io_in, // @[:@30306.4]
  output [31:0] io_out // @[:@30306.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30308.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30308.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30308.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30308.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30308.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30308.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@30308.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30321.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30320.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30319.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30318.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30317.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30315.4]
endmodule
module fix2fixBox_152( // @[:@30492.2]
  input  [31:0] io_a, // @[:@30495.4]
  output [31:0] io_b // @[:@30495.4]
);
  wire [24:0] new_dec; // @[Converter.scala 63:26:@30505.4]
  assign new_dec = io_a[24:0]; // @[Converter.scala 63:26:@30505.4]
  assign io_b = {new_dec,7'h0}; // @[Converter.scala 94:38:@30508.4]
endmodule
module x333( // @[:@30510.2]
  input  [31:0] io_b, // @[:@30513.4]
  output [31:0] io_result // @[:@30513.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@30518.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@30518.4]
  fix2fixBox_152 fix2fixBox ( // @[BigIPZynq.scala 219:30:@30518.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@30526.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@30521.4]
endmodule
module Multiplier( // @[:@30538.2]
  input         clock, // @[:@30539.4]
  input         io_flow, // @[:@30541.4]
  input  [38:0] io_a, // @[:@30541.4]
  input  [38:0] io_b, // @[:@30541.4]
  output [38:0] io_out // @[:@30541.4]
);
  wire [38:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@30543.4]
  wire [38:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@30543.4]
  wire [38:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@30543.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@30543.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@30543.4]
  mul_39_39_39_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@30543.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@30553.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@30551.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@30550.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@30552.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@30549.4]
endmodule
module fix2fixBox_153( // @[:@30555.2]
  input  [38:0] io_a, // @[:@30558.4]
  output [31:0] io_b // @[:@30558.4]
);
  wire [6:0] tmp_frac; // @[Converter.scala 38:42:@30566.4]
  wire [24:0] new_dec; // @[Converter.scala 88:34:@30569.4]
  assign tmp_frac = io_a[13:7]; // @[Converter.scala 38:42:@30566.4]
  assign new_dec = io_a[38:14]; // @[Converter.scala 88:34:@30569.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@30572.4]
endmodule
module x334_mul( // @[:@30574.2]
  input         clock, // @[:@30575.4]
  input  [31:0] io_a, // @[:@30577.4]
  input  [31:0] io_b, // @[:@30577.4]
  input         io_flow, // @[:@30577.4]
  output [31:0] io_result // @[:@30577.4]
);
  wire  x334_mul_clock; // @[BigIPZynq.scala 63:21:@30592.4]
  wire  x334_mul_io_flow; // @[BigIPZynq.scala 63:21:@30592.4]
  wire [38:0] x334_mul_io_a; // @[BigIPZynq.scala 63:21:@30592.4]
  wire [38:0] x334_mul_io_b; // @[BigIPZynq.scala 63:21:@30592.4]
  wire [38:0] x334_mul_io_out; // @[BigIPZynq.scala 63:21:@30592.4]
  wire [38:0] fix2fixBox_io_a; // @[Math.scala 253:30:@30600.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@30600.4]
  wire  _T_16; // @[FixedPoint.scala 50:25:@30584.4]
  wire [6:0] _T_20; // @[Bitwise.scala 72:12:@30586.4]
  wire  _T_22; // @[FixedPoint.scala 50:25:@30588.4]
  wire [6:0] _T_26; // @[Bitwise.scala 72:12:@30590.4]
  Multiplier x334_mul ( // @[BigIPZynq.scala 63:21:@30592.4]
    .clock(x334_mul_clock),
    .io_flow(x334_mul_io_flow),
    .io_a(x334_mul_io_a),
    .io_b(x334_mul_io_b),
    .io_out(x334_mul_io_out)
  );
  fix2fixBox_153 fix2fixBox ( // @[Math.scala 253:30:@30600.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_16 = io_a[31]; // @[FixedPoint.scala 50:25:@30584.4]
  assign _T_20 = _T_16 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@30586.4]
  assign _T_22 = io_b[31]; // @[FixedPoint.scala 50:25:@30588.4]
  assign _T_26 = _T_22 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@30590.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@30608.4]
  assign x334_mul_clock = clock; // @[:@30593.4]
  assign x334_mul_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@30597.4]
  assign x334_mul_io_a = {_T_20,io_a}; // @[BigIPZynq.scala 64:14:@30595.4]
  assign x334_mul_io_b = {_T_26,io_b}; // @[BigIPZynq.scala 65:14:@30596.4]
  assign fix2fixBox_io_a = x334_mul_io_out; // @[Math.scala 254:23:@30603.4]
endmodule
module fix2fixBox_154( // @[:@30610.2]
  input  [31:0] io_a, // @[:@30613.4]
  output [31:0] io_b // @[:@30613.4]
);
  wire [24:0] _T_25; // @[Converter.scala 84:75:@30625.4]
  assign _T_25 = io_a[31:7]; // @[Converter.scala 84:75:@30625.4]
  assign io_b = {7'h0,_T_25}; // @[Converter.scala 95:38:@30628.4]
endmodule
module x335( // @[:@30630.2]
  input  [31:0] io_b, // @[:@30633.4]
  output [31:0] io_result // @[:@30633.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@30638.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@30638.4]
  fix2fixBox_154 fix2fixBox ( // @[BigIPZynq.scala 219:30:@30638.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@30646.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@30641.4]
endmodule
module RetimeWrapper_347( // @[:@30660.2]
  input   clock, // @[:@30661.4]
  input   reset, // @[:@30662.4]
  input   io_flow, // @[:@30663.4]
  input   io_in, // @[:@30663.4]
  output  io_out // @[:@30663.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@30665.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@30665.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@30665.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30665.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30665.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30665.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(58)) sr ( // @[RetimeShiftRegister.scala 15:20:@30665.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30678.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30677.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@30676.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30675.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30674.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30672.4]
endmodule
module RetimeWrapper_348( // @[:@30692.2]
  input         clock, // @[:@30693.4]
  input         reset, // @[:@30694.4]
  input         io_flow, // @[:@30695.4]
  input  [31:0] io_in, // @[:@30695.4]
  output [31:0] io_out // @[:@30695.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30697.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30697.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30697.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30697.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30697.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30697.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(50)) sr ( // @[RetimeShiftRegister.scala 15:20:@30697.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30710.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30709.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30708.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30707.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30706.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30704.4]
endmodule
module RetimeWrapper_350( // @[:@30756.2]
  input         clock, // @[:@30757.4]
  input         reset, // @[:@30758.4]
  input         io_flow, // @[:@30759.4]
  input  [31:0] io_in, // @[:@30759.4]
  output [31:0] io_out // @[:@30759.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30761.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30761.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30761.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30761.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30761.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30761.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(58)) sr ( // @[RetimeShiftRegister.scala 15:20:@30761.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30774.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30773.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30772.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30771.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30770.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30768.4]
endmodule
module RetimeWrapper_354( // @[:@30884.2]
  input   clock, // @[:@30885.4]
  input   reset, // @[:@30886.4]
  input   io_flow, // @[:@30887.4]
  input   io_in, // @[:@30887.4]
  output  io_out // @[:@30887.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@30889.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@30889.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@30889.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30889.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30889.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30889.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(35)) sr ( // @[RetimeShiftRegister.scala 15:20:@30889.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30902.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30901.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@30900.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30899.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30898.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30896.4]
endmodule
module RetimeWrapper_355( // @[:@30916.2]
  input   clock, // @[:@30917.4]
  input   reset, // @[:@30918.4]
  input   io_flow, // @[:@30919.4]
  input   io_in, // @[:@30919.4]
  output  io_out // @[:@30919.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@30921.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@30921.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@30921.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30921.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30921.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30921.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(59)) sr ( // @[RetimeShiftRegister.scala 15:20:@30921.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30934.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30933.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@30932.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30931.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30930.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30928.4]
endmodule
module RetimeWrapper_356( // @[:@30948.2]
  input         clock, // @[:@30949.4]
  input         reset, // @[:@30950.4]
  input         io_flow, // @[:@30951.4]
  input  [31:0] io_in, // @[:@30951.4]
  output [31:0] io_out // @[:@30951.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30953.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30953.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30953.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30953.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30953.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30953.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(51)) sr ( // @[RetimeShiftRegister.scala 15:20:@30953.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30966.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30965.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30964.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30963.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30962.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30960.4]
endmodule
module RetimeWrapper_358( // @[:@31012.2]
  input         clock, // @[:@31013.4]
  input         reset, // @[:@31014.4]
  input         io_flow, // @[:@31015.4]
  input  [31:0] io_in, // @[:@31015.4]
  output [31:0] io_out // @[:@31015.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31017.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31017.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31017.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31017.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31017.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31017.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(59)) sr ( // @[RetimeShiftRegister.scala 15:20:@31017.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31030.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31029.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31028.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31027.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31026.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31024.4]
endmodule
module RetimeWrapper_359( // @[:@31044.2]
  input         clock, // @[:@31045.4]
  input         reset, // @[:@31046.4]
  input         io_flow, // @[:@31047.4]
  input  [31:0] io_in, // @[:@31047.4]
  output [31:0] io_out // @[:@31047.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31049.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31049.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31049.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31049.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31049.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31049.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(38)) sr ( // @[RetimeShiftRegister.scala 15:20:@31049.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31062.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31061.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31060.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31059.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31058.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31056.4]
endmodule
module RetimeWrapper_361( // @[:@31108.2]
  input         clock, // @[:@31109.4]
  input         reset, // @[:@31110.4]
  input         io_flow, // @[:@31111.4]
  input  [31:0] io_in, // @[:@31111.4]
  output [31:0] io_out // @[:@31111.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31113.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31113.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31113.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31113.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31113.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31113.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(27)) sr ( // @[RetimeShiftRegister.scala 15:20:@31113.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31126.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31125.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31124.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31123.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31122.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31120.4]
endmodule
module RetimeWrapper_362( // @[:@31140.2]
  input         clock, // @[:@31141.4]
  input         reset, // @[:@31142.4]
  input         io_flow, // @[:@31143.4]
  input  [31:0] io_in, // @[:@31143.4]
  output [31:0] io_out // @[:@31143.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31145.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31145.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31145.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31145.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31145.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31145.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(14)) sr ( // @[RetimeShiftRegister.scala 15:20:@31145.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31158.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31157.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31156.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31155.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31154.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31152.4]
endmodule
module RetimeWrapper_363( // @[:@31172.2]
  input   clock, // @[:@31173.4]
  input   reset, // @[:@31174.4]
  input   io_flow, // @[:@31175.4]
  input   io_in, // @[:@31175.4]
  output  io_out // @[:@31175.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@31177.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@31177.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@31177.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31177.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31177.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31177.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(34)) sr ( // @[RetimeShiftRegister.scala 15:20:@31177.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31190.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31189.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@31188.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31187.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31186.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31184.4]
endmodule
module RetimeWrapper_365( // @[:@31236.2]
  input         clock, // @[:@31237.4]
  input         reset, // @[:@31238.4]
  input         io_flow, // @[:@31239.4]
  input  [31:0] io_in, // @[:@31239.4]
  output [31:0] io_out // @[:@31239.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31241.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31241.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31241.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31241.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31241.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31241.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(34)) sr ( // @[RetimeShiftRegister.scala 15:20:@31241.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31254.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31253.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31252.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31251.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31250.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31248.4]
endmodule
module RetimeWrapper_366( // @[:@31268.2]
  input         clock, // @[:@31269.4]
  input         reset, // @[:@31270.4]
  input         io_flow, // @[:@31271.4]
  input  [31:0] io_in, // @[:@31271.4]
  output [31:0] io_out // @[:@31271.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31273.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31273.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31273.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31273.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31273.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31273.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(15)) sr ( // @[RetimeShiftRegister.scala 15:20:@31273.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31286.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31285.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31284.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31283.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31282.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31280.4]
endmodule
module RetimeWrapper_372( // @[:@31460.2]
  input         clock, // @[:@31461.4]
  input         reset, // @[:@31462.4]
  input         io_flow, // @[:@31463.4]
  input  [32:0] io_in, // @[:@31463.4]
  output [32:0] io_out // @[:@31463.4]
);
  wire [32:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31465.4]
  wire [32:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31465.4]
  wire [32:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31465.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31465.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31465.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31465.4]
  RetimeShiftRegister #(.WIDTH(33), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@31465.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31478.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31477.4]
  assign sr_init = 33'h0; // @[RetimeShiftRegister.scala 19:16:@31476.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31475.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31474.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31472.4]
endmodule
module RetimeWrapper_373( // @[:@31492.2]
  input         clock, // @[:@31493.4]
  input         reset, // @[:@31494.4]
  input         io_flow, // @[:@31495.4]
  input  [33:0] io_in, // @[:@31495.4]
  output [33:0] io_out // @[:@31495.4]
);
  wire [33:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31497.4]
  wire [33:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31497.4]
  wire [33:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31497.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31497.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31497.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31497.4]
  RetimeShiftRegister #(.WIDTH(34), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@31497.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31510.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31509.4]
  assign sr_init = 34'h0; // @[RetimeShiftRegister.scala 19:16:@31508.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31507.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31506.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31504.4]
endmodule
module RetimeWrapper_380( // @[:@32283.2]
  input   clock, // @[:@32284.4]
  input   reset, // @[:@32285.4]
  input   io_flow, // @[:@32286.4]
  input   io_in, // @[:@32286.4]
  output  io_out // @[:@32286.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@32288.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@32288.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@32288.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@32288.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@32288.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@32288.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(73)) sr ( // @[RetimeShiftRegister.scala 15:20:@32288.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@32301.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@32300.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@32299.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@32298.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@32297.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@32295.4]
endmodule
module x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@32367.2]
  input          clock, // @[:@32368.4]
  input          reset, // @[:@32369.4]
  output         io_in_x209_TREADY, // @[:@32370.4]
  input  [255:0] io_in_x209_TDATA, // @[:@32370.4]
  input  [7:0]   io_in_x209_TID, // @[:@32370.4]
  input  [7:0]   io_in_x209_TDEST, // @[:@32370.4]
  output         io_in_x210_TVALID, // @[:@32370.4]
  input          io_in_x210_TREADY, // @[:@32370.4]
  output [255:0] io_in_x210_TDATA, // @[:@32370.4]
  input          io_sigsIn_backpressure, // @[:@32370.4]
  input          io_sigsIn_datapathEn, // @[:@32370.4]
  input          io_sigsIn_break, // @[:@32370.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@32370.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@32370.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@32370.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@32370.4]
  input          io_rr // @[:@32370.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@32384.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@32384.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@32396.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@32396.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32419.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32419.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32419.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@32419.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@32419.4]
  wire  x241_lb_0_clock; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_reset; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [1:0] x241_lb_0_io_rPort_8_banks_1; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [2:0] x241_lb_0_io_rPort_8_banks_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [9:0] x241_lb_0_io_rPort_8_ofs_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_8_en_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_8_backpressure; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [31:0] x241_lb_0_io_rPort_8_output_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [1:0] x241_lb_0_io_rPort_7_banks_1; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [2:0] x241_lb_0_io_rPort_7_banks_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [9:0] x241_lb_0_io_rPort_7_ofs_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_7_en_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_7_backpressure; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [31:0] x241_lb_0_io_rPort_7_output_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [1:0] x241_lb_0_io_rPort_6_banks_1; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [2:0] x241_lb_0_io_rPort_6_banks_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [9:0] x241_lb_0_io_rPort_6_ofs_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_6_en_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_6_backpressure; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [31:0] x241_lb_0_io_rPort_6_output_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [1:0] x241_lb_0_io_rPort_5_banks_1; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [2:0] x241_lb_0_io_rPort_5_banks_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [9:0] x241_lb_0_io_rPort_5_ofs_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_5_en_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_5_backpressure; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [31:0] x241_lb_0_io_rPort_5_output_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [1:0] x241_lb_0_io_rPort_4_banks_1; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [2:0] x241_lb_0_io_rPort_4_banks_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [9:0] x241_lb_0_io_rPort_4_ofs_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_4_en_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_4_backpressure; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [31:0] x241_lb_0_io_rPort_4_output_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [1:0] x241_lb_0_io_rPort_3_banks_1; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [2:0] x241_lb_0_io_rPort_3_banks_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [9:0] x241_lb_0_io_rPort_3_ofs_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_3_en_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_3_backpressure; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [31:0] x241_lb_0_io_rPort_3_output_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [1:0] x241_lb_0_io_rPort_2_banks_1; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [2:0] x241_lb_0_io_rPort_2_banks_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [9:0] x241_lb_0_io_rPort_2_ofs_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_2_en_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_2_backpressure; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [31:0] x241_lb_0_io_rPort_2_output_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [1:0] x241_lb_0_io_rPort_1_banks_1; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [2:0] x241_lb_0_io_rPort_1_banks_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [9:0] x241_lb_0_io_rPort_1_ofs_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_1_en_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_1_backpressure; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [31:0] x241_lb_0_io_rPort_1_output_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [1:0] x241_lb_0_io_rPort_0_banks_1; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [2:0] x241_lb_0_io_rPort_0_banks_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [9:0] x241_lb_0_io_rPort_0_ofs_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_0_en_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_rPort_0_backpressure; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [31:0] x241_lb_0_io_rPort_0_output_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [1:0] x241_lb_0_io_wPort_0_banks_1; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [2:0] x241_lb_0_io_wPort_0_banks_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [9:0] x241_lb_0_io_wPort_0_ofs_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire [31:0] x241_lb_0_io_wPort_0_data_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x241_lb_0_io_wPort_0_en_0; // @[m_x241_lb_0.scala 35:17:@32429.4]
  wire  x242_lb2_0_clock; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire  x242_lb2_0_reset; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [1:0] x242_lb2_0_io_rPort_3_banks_1; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [2:0] x242_lb2_0_io_rPort_3_banks_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [9:0] x242_lb2_0_io_rPort_3_ofs_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire  x242_lb2_0_io_rPort_3_en_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire  x242_lb2_0_io_rPort_3_backpressure; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [31:0] x242_lb2_0_io_rPort_3_output_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [1:0] x242_lb2_0_io_rPort_2_banks_1; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [2:0] x242_lb2_0_io_rPort_2_banks_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [9:0] x242_lb2_0_io_rPort_2_ofs_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire  x242_lb2_0_io_rPort_2_en_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire  x242_lb2_0_io_rPort_2_backpressure; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [31:0] x242_lb2_0_io_rPort_2_output_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [1:0] x242_lb2_0_io_rPort_1_banks_1; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [2:0] x242_lb2_0_io_rPort_1_banks_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [9:0] x242_lb2_0_io_rPort_1_ofs_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire  x242_lb2_0_io_rPort_1_en_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire  x242_lb2_0_io_rPort_1_backpressure; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [31:0] x242_lb2_0_io_rPort_1_output_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [1:0] x242_lb2_0_io_rPort_0_banks_1; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [2:0] x242_lb2_0_io_rPort_0_banks_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [9:0] x242_lb2_0_io_rPort_0_ofs_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire  x242_lb2_0_io_rPort_0_en_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire  x242_lb2_0_io_rPort_0_backpressure; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [31:0] x242_lb2_0_io_rPort_0_output_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [1:0] x242_lb2_0_io_wPort_0_banks_1; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [2:0] x242_lb2_0_io_wPort_0_banks_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [9:0] x242_lb2_0_io_wPort_0_ofs_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire [31:0] x242_lb2_0_io_wPort_0_data_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire  x242_lb2_0_io_wPort_0_en_0; // @[m_x242_lb2_0.scala 30:17:@32496.4]
  wire  x416_sum_1_clock; // @[Math.scala 150:24:@32591.4]
  wire  x416_sum_1_reset; // @[Math.scala 150:24:@32591.4]
  wire [31:0] x416_sum_1_io_a; // @[Math.scala 150:24:@32591.4]
  wire [31:0] x416_sum_1_io_b; // @[Math.scala 150:24:@32591.4]
  wire  x416_sum_1_io_flow; // @[Math.scala 150:24:@32591.4]
  wire [31:0] x416_sum_1_io_result; // @[Math.scala 150:24:@32591.4]
  wire  x419_sum_1_clock; // @[Math.scala 150:24:@32629.4]
  wire  x419_sum_1_reset; // @[Math.scala 150:24:@32629.4]
  wire [31:0] x419_sum_1_io_a; // @[Math.scala 150:24:@32629.4]
  wire [31:0] x419_sum_1_io_b; // @[Math.scala 150:24:@32629.4]
  wire  x419_sum_1_io_flow; // @[Math.scala 150:24:@32629.4]
  wire [31:0] x419_sum_1_io_result; // @[Math.scala 150:24:@32629.4]
  wire  x422_sum_1_clock; // @[Math.scala 150:24:@32667.4]
  wire  x422_sum_1_reset; // @[Math.scala 150:24:@32667.4]
  wire [31:0] x422_sum_1_io_a; // @[Math.scala 150:24:@32667.4]
  wire [31:0] x422_sum_1_io_b; // @[Math.scala 150:24:@32667.4]
  wire  x422_sum_1_io_flow; // @[Math.scala 150:24:@32667.4]
  wire [31:0] x422_sum_1_io_result; // @[Math.scala 150:24:@32667.4]
  wire  x425_sum_1_clock; // @[Math.scala 150:24:@32705.4]
  wire  x425_sum_1_reset; // @[Math.scala 150:24:@32705.4]
  wire [31:0] x425_sum_1_io_a; // @[Math.scala 150:24:@32705.4]
  wire [31:0] x425_sum_1_io_b; // @[Math.scala 150:24:@32705.4]
  wire  x425_sum_1_io_flow; // @[Math.scala 150:24:@32705.4]
  wire [31:0] x425_sum_1_io_result; // @[Math.scala 150:24:@32705.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32728.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32728.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32728.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@32728.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@32728.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@32746.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@32746.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@32746.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@32746.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@32746.4]
  wire  x428_sum_1_clock; // @[Math.scala 150:24:@32759.4]
  wire  x428_sum_1_reset; // @[Math.scala 150:24:@32759.4]
  wire [31:0] x428_sum_1_io_a; // @[Math.scala 150:24:@32759.4]
  wire [31:0] x428_sum_1_io_b; // @[Math.scala 150:24:@32759.4]
  wire  x428_sum_1_io_flow; // @[Math.scala 150:24:@32759.4]
  wire [31:0] x428_sum_1_io_result; // @[Math.scala 150:24:@32759.4]
  wire  x431_sum_1_clock; // @[Math.scala 150:24:@32797.4]
  wire  x431_sum_1_reset; // @[Math.scala 150:24:@32797.4]
  wire [31:0] x431_sum_1_io_a; // @[Math.scala 150:24:@32797.4]
  wire [31:0] x431_sum_1_io_b; // @[Math.scala 150:24:@32797.4]
  wire  x431_sum_1_io_flow; // @[Math.scala 150:24:@32797.4]
  wire [31:0] x431_sum_1_io_result; // @[Math.scala 150:24:@32797.4]
  wire  x434_sub_1_clock; // @[Math.scala 191:24:@32823.4]
  wire  x434_sub_1_reset; // @[Math.scala 191:24:@32823.4]
  wire [31:0] x434_sub_1_io_a; // @[Math.scala 191:24:@32823.4]
  wire [31:0] x434_sub_1_io_b; // @[Math.scala 191:24:@32823.4]
  wire  x434_sub_1_io_flow; // @[Math.scala 191:24:@32823.4]
  wire [31:0] x434_sub_1_io_result; // @[Math.scala 191:24:@32823.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@32833.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@32833.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@32833.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@32833.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@32833.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@32842.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@32842.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@32842.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@32842.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@32842.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@32851.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@32851.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@32851.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@32851.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@32851.4]
  wire  x438_sum_1_clock; // @[Math.scala 150:24:@32890.4]
  wire  x438_sum_1_reset; // @[Math.scala 150:24:@32890.4]
  wire [31:0] x438_sum_1_io_a; // @[Math.scala 150:24:@32890.4]
  wire [31:0] x438_sum_1_io_b; // @[Math.scala 150:24:@32890.4]
  wire  x438_sum_1_io_flow; // @[Math.scala 150:24:@32890.4]
  wire [31:0] x438_sum_1_io_result; // @[Math.scala 150:24:@32890.4]
  wire  x250_div_1_clock; // @[Math.scala 327:24:@32902.4]
  wire [31:0] x250_div_1_io_a; // @[Math.scala 327:24:@32902.4]
  wire  x250_div_1_io_flow; // @[Math.scala 327:24:@32902.4]
  wire [31:0] x250_div_1_io_result; // @[Math.scala 327:24:@32902.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@32912.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@32912.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@32912.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@32912.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@32912.4]
  wire  x251_sum_1_clock; // @[Math.scala 150:24:@32921.4]
  wire  x251_sum_1_reset; // @[Math.scala 150:24:@32921.4]
  wire [31:0] x251_sum_1_io_a; // @[Math.scala 150:24:@32921.4]
  wire [31:0] x251_sum_1_io_b; // @[Math.scala 150:24:@32921.4]
  wire  x251_sum_1_io_flow; // @[Math.scala 150:24:@32921.4]
  wire [31:0] x251_sum_1_io_result; // @[Math.scala 150:24:@32921.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@32931.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@32931.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@32931.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@32931.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@32931.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@32940.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@32940.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@32940.4]
  wire [31:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@32940.4]
  wire [31:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@32940.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@32949.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@32949.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@32949.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@32949.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@32949.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@32958.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@32958.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@32958.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@32958.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@32958.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@32967.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@32967.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@32967.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@32967.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@32967.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@32978.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@32978.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@32978.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@32978.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@32978.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@32999.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@32999.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@32999.4]
  wire [31:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@32999.4]
  wire [31:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@32999.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@33015.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@33015.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@33015.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@33015.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@33015.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@33024.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@33024.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@33024.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@33024.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@33024.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@33038.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@33038.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@33038.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@33038.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@33038.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@33053.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@33053.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@33053.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@33053.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@33053.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@33062.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@33062.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@33062.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@33062.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@33062.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@33071.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@33071.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@33071.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@33071.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@33071.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@33080.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@33080.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@33080.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@33080.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@33080.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@33089.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@33089.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@33089.4]
  wire [31:0] RetimeWrapper_21_io_in; // @[package.scala 93:22:@33089.4]
  wire [31:0] RetimeWrapper_21_io_out; // @[package.scala 93:22:@33089.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@33098.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@33098.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@33098.4]
  wire [31:0] RetimeWrapper_22_io_in; // @[package.scala 93:22:@33098.4]
  wire [31:0] RetimeWrapper_22_io_out; // @[package.scala 93:22:@33098.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@33110.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@33110.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@33110.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@33110.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@33110.4]
  wire  x260_rdcol_1_clock; // @[Math.scala 191:24:@33133.4]
  wire  x260_rdcol_1_reset; // @[Math.scala 191:24:@33133.4]
  wire [31:0] x260_rdcol_1_io_a; // @[Math.scala 191:24:@33133.4]
  wire [31:0] x260_rdcol_1_io_b; // @[Math.scala 191:24:@33133.4]
  wire  x260_rdcol_1_io_flow; // @[Math.scala 191:24:@33133.4]
  wire [31:0] x260_rdcol_1_io_result; // @[Math.scala 191:24:@33133.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@33148.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@33148.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@33148.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@33148.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@33148.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@33157.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@33157.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@33157.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@33157.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@33157.4]
  wire  x441_sum_1_clock; // @[Math.scala 150:24:@33200.4]
  wire  x441_sum_1_reset; // @[Math.scala 150:24:@33200.4]
  wire [31:0] x441_sum_1_io_a; // @[Math.scala 150:24:@33200.4]
  wire [31:0] x441_sum_1_io_b; // @[Math.scala 150:24:@33200.4]
  wire  x441_sum_1_io_flow; // @[Math.scala 150:24:@33200.4]
  wire [31:0] x441_sum_1_io_result; // @[Math.scala 150:24:@33200.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@33223.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@33223.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@33223.4]
  wire [31:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@33223.4]
  wire [31:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@33223.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@33241.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@33241.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@33241.4]
  wire [31:0] RetimeWrapper_27_io_in; // @[package.scala 93:22:@33241.4]
  wire [31:0] RetimeWrapper_27_io_out; // @[package.scala 93:22:@33241.4]
  wire  x444_sum_1_clock; // @[Math.scala 150:24:@33254.4]
  wire  x444_sum_1_reset; // @[Math.scala 150:24:@33254.4]
  wire [31:0] x444_sum_1_io_a; // @[Math.scala 150:24:@33254.4]
  wire [31:0] x444_sum_1_io_b; // @[Math.scala 150:24:@33254.4]
  wire  x444_sum_1_io_flow; // @[Math.scala 150:24:@33254.4]
  wire [31:0] x444_sum_1_io_result; // @[Math.scala 150:24:@33254.4]
  wire  x447_sum_1_clock; // @[Math.scala 150:24:@33292.4]
  wire  x447_sum_1_reset; // @[Math.scala 150:24:@33292.4]
  wire [31:0] x447_sum_1_io_a; // @[Math.scala 150:24:@33292.4]
  wire [31:0] x447_sum_1_io_b; // @[Math.scala 150:24:@33292.4]
  wire  x447_sum_1_io_flow; // @[Math.scala 150:24:@33292.4]
  wire [31:0] x447_sum_1_io_result; // @[Math.scala 150:24:@33292.4]
  wire  x450_sum_1_clock; // @[Math.scala 150:24:@33330.4]
  wire  x450_sum_1_reset; // @[Math.scala 150:24:@33330.4]
  wire [31:0] x450_sum_1_io_a; // @[Math.scala 150:24:@33330.4]
  wire [31:0] x450_sum_1_io_b; // @[Math.scala 150:24:@33330.4]
  wire  x450_sum_1_io_flow; // @[Math.scala 150:24:@33330.4]
  wire [31:0] x450_sum_1_io_result; // @[Math.scala 150:24:@33330.4]
  wire  x453_sum_1_clock; // @[Math.scala 150:24:@33368.4]
  wire  x453_sum_1_reset; // @[Math.scala 150:24:@33368.4]
  wire [31:0] x453_sum_1_io_a; // @[Math.scala 150:24:@33368.4]
  wire [31:0] x453_sum_1_io_b; // @[Math.scala 150:24:@33368.4]
  wire  x453_sum_1_io_flow; // @[Math.scala 150:24:@33368.4]
  wire [31:0] x453_sum_1_io_result; // @[Math.scala 150:24:@33368.4]
  wire  x456_sum_1_clock; // @[Math.scala 150:24:@33406.4]
  wire  x456_sum_1_reset; // @[Math.scala 150:24:@33406.4]
  wire [31:0] x456_sum_1_io_a; // @[Math.scala 150:24:@33406.4]
  wire [31:0] x456_sum_1_io_b; // @[Math.scala 150:24:@33406.4]
  wire  x456_sum_1_io_flow; // @[Math.scala 150:24:@33406.4]
  wire [31:0] x456_sum_1_io_result; // @[Math.scala 150:24:@33406.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@33421.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@33421.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@33421.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@33421.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@33421.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@33435.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@33435.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@33435.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@33435.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@33435.4]
  wire  x459_sub_1_clock; // @[Math.scala 191:24:@33446.4]
  wire  x459_sub_1_reset; // @[Math.scala 191:24:@33446.4]
  wire [31:0] x459_sub_1_io_a; // @[Math.scala 191:24:@33446.4]
  wire [31:0] x459_sub_1_io_b; // @[Math.scala 191:24:@33446.4]
  wire  x459_sub_1_io_flow; // @[Math.scala 191:24:@33446.4]
  wire [31:0] x459_sub_1_io_result; // @[Math.scala 191:24:@33446.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@33456.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@33456.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@33456.4]
  wire [31:0] RetimeWrapper_30_io_in; // @[package.scala 93:22:@33456.4]
  wire [31:0] RetimeWrapper_30_io_out; // @[package.scala 93:22:@33456.4]
  wire  x265_div_1_clock; // @[Math.scala 327:24:@33470.4]
  wire [31:0] x265_div_1_io_a; // @[Math.scala 327:24:@33470.4]
  wire  x265_div_1_io_flow; // @[Math.scala 327:24:@33470.4]
  wire [31:0] x265_div_1_io_result; // @[Math.scala 327:24:@33470.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@33480.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@33480.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@33480.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@33480.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@33480.4]
  wire  x266_sum_1_clock; // @[Math.scala 150:24:@33489.4]
  wire  x266_sum_1_reset; // @[Math.scala 150:24:@33489.4]
  wire [31:0] x266_sum_1_io_a; // @[Math.scala 150:24:@33489.4]
  wire [31:0] x266_sum_1_io_b; // @[Math.scala 150:24:@33489.4]
  wire  x266_sum_1_io_flow; // @[Math.scala 150:24:@33489.4]
  wire [31:0] x266_sum_1_io_result; // @[Math.scala 150:24:@33489.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@33499.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@33499.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@33499.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@33499.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@33499.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@33508.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@33508.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@33508.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@33508.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@33508.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@33520.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@33520.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@33520.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@33520.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@33520.4]
  wire  x269_rdcol_1_clock; // @[Math.scala 191:24:@33543.4]
  wire  x269_rdcol_1_reset; // @[Math.scala 191:24:@33543.4]
  wire [31:0] x269_rdcol_1_io_a; // @[Math.scala 191:24:@33543.4]
  wire [31:0] x269_rdcol_1_io_b; // @[Math.scala 191:24:@33543.4]
  wire  x269_rdcol_1_io_flow; // @[Math.scala 191:24:@33543.4]
  wire [31:0] x269_rdcol_1_io_result; // @[Math.scala 191:24:@33543.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@33560.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@33560.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@33560.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@33560.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@33560.4]
  wire  x463_sum_1_clock; // @[Math.scala 150:24:@33603.4]
  wire  x463_sum_1_reset; // @[Math.scala 150:24:@33603.4]
  wire [31:0] x463_sum_1_io_a; // @[Math.scala 150:24:@33603.4]
  wire [31:0] x463_sum_1_io_b; // @[Math.scala 150:24:@33603.4]
  wire  x463_sum_1_io_flow; // @[Math.scala 150:24:@33603.4]
  wire [31:0] x463_sum_1_io_result; // @[Math.scala 150:24:@33603.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@33626.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@33626.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@33626.4]
  wire [31:0] RetimeWrapper_36_io_in; // @[package.scala 93:22:@33626.4]
  wire [31:0] RetimeWrapper_36_io_out; // @[package.scala 93:22:@33626.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@33644.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@33644.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@33644.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@33644.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@33644.4]
  wire  x466_sum_1_clock; // @[Math.scala 150:24:@33657.4]
  wire  x466_sum_1_reset; // @[Math.scala 150:24:@33657.4]
  wire [31:0] x466_sum_1_io_a; // @[Math.scala 150:24:@33657.4]
  wire [31:0] x466_sum_1_io_b; // @[Math.scala 150:24:@33657.4]
  wire  x466_sum_1_io_flow; // @[Math.scala 150:24:@33657.4]
  wire [31:0] x466_sum_1_io_result; // @[Math.scala 150:24:@33657.4]
  wire  x469_sum_1_clock; // @[Math.scala 150:24:@33695.4]
  wire  x469_sum_1_reset; // @[Math.scala 150:24:@33695.4]
  wire [31:0] x469_sum_1_io_a; // @[Math.scala 150:24:@33695.4]
  wire [31:0] x469_sum_1_io_b; // @[Math.scala 150:24:@33695.4]
  wire  x469_sum_1_io_flow; // @[Math.scala 150:24:@33695.4]
  wire [31:0] x469_sum_1_io_result; // @[Math.scala 150:24:@33695.4]
  wire  x472_sum_1_clock; // @[Math.scala 150:24:@33733.4]
  wire  x472_sum_1_reset; // @[Math.scala 150:24:@33733.4]
  wire [31:0] x472_sum_1_io_a; // @[Math.scala 150:24:@33733.4]
  wire [31:0] x472_sum_1_io_b; // @[Math.scala 150:24:@33733.4]
  wire  x472_sum_1_io_flow; // @[Math.scala 150:24:@33733.4]
  wire [31:0] x472_sum_1_io_result; // @[Math.scala 150:24:@33733.4]
  wire  x475_sum_1_clock; // @[Math.scala 150:24:@33771.4]
  wire  x475_sum_1_reset; // @[Math.scala 150:24:@33771.4]
  wire [31:0] x475_sum_1_io_a; // @[Math.scala 150:24:@33771.4]
  wire [31:0] x475_sum_1_io_b; // @[Math.scala 150:24:@33771.4]
  wire  x475_sum_1_io_flow; // @[Math.scala 150:24:@33771.4]
  wire [31:0] x475_sum_1_io_result; // @[Math.scala 150:24:@33771.4]
  wire  x478_sum_1_clock; // @[Math.scala 150:24:@33809.4]
  wire  x478_sum_1_reset; // @[Math.scala 150:24:@33809.4]
  wire [31:0] x478_sum_1_io_a; // @[Math.scala 150:24:@33809.4]
  wire [31:0] x478_sum_1_io_b; // @[Math.scala 150:24:@33809.4]
  wire  x478_sum_1_io_flow; // @[Math.scala 150:24:@33809.4]
  wire [31:0] x478_sum_1_io_result; // @[Math.scala 150:24:@33809.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@33824.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@33824.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@33824.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@33824.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@33824.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@33838.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@33838.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@33838.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@33838.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@33838.4]
  wire  x481_sub_1_clock; // @[Math.scala 191:24:@33849.4]
  wire  x481_sub_1_reset; // @[Math.scala 191:24:@33849.4]
  wire [31:0] x481_sub_1_io_a; // @[Math.scala 191:24:@33849.4]
  wire [31:0] x481_sub_1_io_b; // @[Math.scala 191:24:@33849.4]
  wire  x481_sub_1_io_flow; // @[Math.scala 191:24:@33849.4]
  wire [31:0] x481_sub_1_io_result; // @[Math.scala 191:24:@33849.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@33859.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@33859.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@33859.4]
  wire [31:0] RetimeWrapper_40_io_in; // @[package.scala 93:22:@33859.4]
  wire [31:0] RetimeWrapper_40_io_out; // @[package.scala 93:22:@33859.4]
  wire  x274_div_1_clock; // @[Math.scala 327:24:@33873.4]
  wire [31:0] x274_div_1_io_a; // @[Math.scala 327:24:@33873.4]
  wire  x274_div_1_io_flow; // @[Math.scala 327:24:@33873.4]
  wire [31:0] x274_div_1_io_result; // @[Math.scala 327:24:@33873.4]
  wire  x275_sum_1_clock; // @[Math.scala 150:24:@33883.4]
  wire  x275_sum_1_reset; // @[Math.scala 150:24:@33883.4]
  wire [31:0] x275_sum_1_io_a; // @[Math.scala 150:24:@33883.4]
  wire [31:0] x275_sum_1_io_b; // @[Math.scala 150:24:@33883.4]
  wire  x275_sum_1_io_flow; // @[Math.scala 150:24:@33883.4]
  wire [31:0] x275_sum_1_io_result; // @[Math.scala 150:24:@33883.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@33893.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@33893.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@33893.4]
  wire [31:0] RetimeWrapper_41_io_in; // @[package.scala 93:22:@33893.4]
  wire [31:0] RetimeWrapper_41_io_out; // @[package.scala 93:22:@33893.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@33902.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@33902.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@33902.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@33902.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@33902.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@33914.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@33914.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@33914.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@33914.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@33914.4]
  wire  x278_rdrow_1_clock; // @[Math.scala 191:24:@33937.4]
  wire  x278_rdrow_1_reset; // @[Math.scala 191:24:@33937.4]
  wire [31:0] x278_rdrow_1_io_a; // @[Math.scala 191:24:@33937.4]
  wire [31:0] x278_rdrow_1_io_b; // @[Math.scala 191:24:@33937.4]
  wire  x278_rdrow_1_io_flow; // @[Math.scala 191:24:@33937.4]
  wire [31:0] x278_rdrow_1_io_result; // @[Math.scala 191:24:@33937.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@33963.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@33963.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@33963.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@33963.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@33963.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@33972.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@33972.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@33972.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@33972.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@33972.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@33994.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@33994.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@33994.4]
  wire [31:0] RetimeWrapper_46_io_in; // @[package.scala 93:22:@33994.4]
  wire [31:0] RetimeWrapper_46_io_out; // @[package.scala 93:22:@33994.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@34020.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@34020.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@34020.4]
  wire [31:0] RetimeWrapper_47_io_in; // @[package.scala 93:22:@34020.4]
  wire [31:0] RetimeWrapper_47_io_out; // @[package.scala 93:22:@34020.4]
  wire  x487_sum_1_clock; // @[Math.scala 150:24:@34041.4]
  wire  x487_sum_1_reset; // @[Math.scala 150:24:@34041.4]
  wire [31:0] x487_sum_1_io_a; // @[Math.scala 150:24:@34041.4]
  wire [31:0] x487_sum_1_io_b; // @[Math.scala 150:24:@34041.4]
  wire  x487_sum_1_io_flow; // @[Math.scala 150:24:@34041.4]
  wire [31:0] x487_sum_1_io_result; // @[Math.scala 150:24:@34041.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@34051.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@34051.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@34051.4]
  wire [31:0] RetimeWrapper_48_io_in; // @[package.scala 93:22:@34051.4]
  wire [31:0] RetimeWrapper_48_io_out; // @[package.scala 93:22:@34051.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@34060.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@34060.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@34060.4]
  wire [31:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@34060.4]
  wire [31:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@34060.4]
  wire  x286_sum_1_clock; // @[Math.scala 150:24:@34069.4]
  wire  x286_sum_1_reset; // @[Math.scala 150:24:@34069.4]
  wire [31:0] x286_sum_1_io_a; // @[Math.scala 150:24:@34069.4]
  wire [31:0] x286_sum_1_io_b; // @[Math.scala 150:24:@34069.4]
  wire  x286_sum_1_io_flow; // @[Math.scala 150:24:@34069.4]
  wire [31:0] x286_sum_1_io_result; // @[Math.scala 150:24:@34069.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@34079.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@34079.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@34079.4]
  wire [31:0] RetimeWrapper_50_io_in; // @[package.scala 93:22:@34079.4]
  wire [31:0] RetimeWrapper_50_io_out; // @[package.scala 93:22:@34079.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@34088.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@34088.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@34088.4]
  wire [31:0] RetimeWrapper_51_io_in; // @[package.scala 93:22:@34088.4]
  wire [31:0] RetimeWrapper_51_io_out; // @[package.scala 93:22:@34088.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@34097.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@34097.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@34097.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@34097.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@34097.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@34109.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@34109.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@34109.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@34109.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@34109.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@34136.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@34136.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@34136.4]
  wire [31:0] RetimeWrapper_54_io_in; // @[package.scala 93:22:@34136.4]
  wire [31:0] RetimeWrapper_54_io_out; // @[package.scala 93:22:@34136.4]
  wire  x291_sum_1_clock; // @[Math.scala 150:24:@34147.4]
  wire  x291_sum_1_reset; // @[Math.scala 150:24:@34147.4]
  wire [31:0] x291_sum_1_io_a; // @[Math.scala 150:24:@34147.4]
  wire [31:0] x291_sum_1_io_b; // @[Math.scala 150:24:@34147.4]
  wire  x291_sum_1_io_flow; // @[Math.scala 150:24:@34147.4]
  wire [31:0] x291_sum_1_io_result; // @[Math.scala 150:24:@34147.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@34157.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@34157.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@34157.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@34157.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@34157.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@34169.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@34169.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@34169.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@34169.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@34169.4]
  wire  x296_sum_1_clock; // @[Math.scala 150:24:@34196.4]
  wire  x296_sum_1_reset; // @[Math.scala 150:24:@34196.4]
  wire [31:0] x296_sum_1_io_a; // @[Math.scala 150:24:@34196.4]
  wire [31:0] x296_sum_1_io_b; // @[Math.scala 150:24:@34196.4]
  wire  x296_sum_1_io_flow; // @[Math.scala 150:24:@34196.4]
  wire [31:0] x296_sum_1_io_result; // @[Math.scala 150:24:@34196.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@34206.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@34206.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@34206.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@34206.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@34206.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@34218.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@34218.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@34218.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@34218.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@34218.4]
  wire  x299_rdrow_1_clock; // @[Math.scala 191:24:@34241.4]
  wire  x299_rdrow_1_reset; // @[Math.scala 191:24:@34241.4]
  wire [31:0] x299_rdrow_1_io_a; // @[Math.scala 191:24:@34241.4]
  wire [31:0] x299_rdrow_1_io_b; // @[Math.scala 191:24:@34241.4]
  wire  x299_rdrow_1_io_flow; // @[Math.scala 191:24:@34241.4]
  wire [31:0] x299_rdrow_1_io_result; // @[Math.scala 191:24:@34241.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@34267.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@34267.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@34267.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@34267.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@34267.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@34289.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@34289.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@34289.4]
  wire [31:0] RetimeWrapper_60_io_in; // @[package.scala 93:22:@34289.4]
  wire [31:0] RetimeWrapper_60_io_out; // @[package.scala 93:22:@34289.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@34315.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@34315.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@34315.4]
  wire [31:0] RetimeWrapper_61_io_in; // @[package.scala 93:22:@34315.4]
  wire [31:0] RetimeWrapper_61_io_out; // @[package.scala 93:22:@34315.4]
  wire  x492_sum_1_clock; // @[Math.scala 150:24:@34336.4]
  wire  x492_sum_1_reset; // @[Math.scala 150:24:@34336.4]
  wire [31:0] x492_sum_1_io_a; // @[Math.scala 150:24:@34336.4]
  wire [31:0] x492_sum_1_io_b; // @[Math.scala 150:24:@34336.4]
  wire  x492_sum_1_io_flow; // @[Math.scala 150:24:@34336.4]
  wire [31:0] x492_sum_1_io_result; // @[Math.scala 150:24:@34336.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@34346.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@34346.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@34346.4]
  wire [31:0] RetimeWrapper_62_io_in; // @[package.scala 93:22:@34346.4]
  wire [31:0] RetimeWrapper_62_io_out; // @[package.scala 93:22:@34346.4]
  wire  x307_sum_1_clock; // @[Math.scala 150:24:@34355.4]
  wire  x307_sum_1_reset; // @[Math.scala 150:24:@34355.4]
  wire [31:0] x307_sum_1_io_a; // @[Math.scala 150:24:@34355.4]
  wire [31:0] x307_sum_1_io_b; // @[Math.scala 150:24:@34355.4]
  wire  x307_sum_1_io_flow; // @[Math.scala 150:24:@34355.4]
  wire [31:0] x307_sum_1_io_result; // @[Math.scala 150:24:@34355.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@34365.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@34365.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@34365.4]
  wire [31:0] RetimeWrapper_63_io_in; // @[package.scala 93:22:@34365.4]
  wire [31:0] RetimeWrapper_63_io_out; // @[package.scala 93:22:@34365.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@34374.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@34374.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@34374.4]
  wire [31:0] RetimeWrapper_64_io_in; // @[package.scala 93:22:@34374.4]
  wire [31:0] RetimeWrapper_64_io_out; // @[package.scala 93:22:@34374.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@34383.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@34383.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@34383.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@34383.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@34383.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@34395.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@34395.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@34395.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@34395.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@34395.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@34422.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@34422.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@34422.4]
  wire [31:0] RetimeWrapper_67_io_in; // @[package.scala 93:22:@34422.4]
  wire [31:0] RetimeWrapper_67_io_out; // @[package.scala 93:22:@34422.4]
  wire  x312_sum_1_clock; // @[Math.scala 150:24:@34431.4]
  wire  x312_sum_1_reset; // @[Math.scala 150:24:@34431.4]
  wire [31:0] x312_sum_1_io_a; // @[Math.scala 150:24:@34431.4]
  wire [31:0] x312_sum_1_io_b; // @[Math.scala 150:24:@34431.4]
  wire  x312_sum_1_io_flow; // @[Math.scala 150:24:@34431.4]
  wire [31:0] x312_sum_1_io_result; // @[Math.scala 150:24:@34431.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@34441.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@34441.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@34441.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@34441.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@34441.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@34453.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@34453.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@34453.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@34453.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@34453.4]
  wire  x317_sum_1_clock; // @[Math.scala 150:24:@34480.4]
  wire  x317_sum_1_reset; // @[Math.scala 150:24:@34480.4]
  wire [31:0] x317_sum_1_io_a; // @[Math.scala 150:24:@34480.4]
  wire [31:0] x317_sum_1_io_b; // @[Math.scala 150:24:@34480.4]
  wire  x317_sum_1_io_flow; // @[Math.scala 150:24:@34480.4]
  wire [31:0] x317_sum_1_io_result; // @[Math.scala 150:24:@34480.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@34490.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@34490.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@34490.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@34490.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@34490.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@34502.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@34502.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@34502.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@34502.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@34502.4]
  wire  x325_x7_1_clock; // @[Math.scala 150:24:@34550.4]
  wire  x325_x7_1_reset; // @[Math.scala 150:24:@34550.4]
  wire [31:0] x325_x7_1_io_a; // @[Math.scala 150:24:@34550.4]
  wire [31:0] x325_x7_1_io_b; // @[Math.scala 150:24:@34550.4]
  wire  x325_x7_1_io_flow; // @[Math.scala 150:24:@34550.4]
  wire [31:0] x325_x7_1_io_result; // @[Math.scala 150:24:@34550.4]
  wire  x326_x8_1_clock; // @[Math.scala 150:24:@34560.4]
  wire  x326_x8_1_reset; // @[Math.scala 150:24:@34560.4]
  wire [31:0] x326_x8_1_io_a; // @[Math.scala 150:24:@34560.4]
  wire [31:0] x326_x8_1_io_b; // @[Math.scala 150:24:@34560.4]
  wire  x326_x8_1_io_flow; // @[Math.scala 150:24:@34560.4]
  wire [31:0] x326_x8_1_io_result; // @[Math.scala 150:24:@34560.4]
  wire  x327_x7_1_clock; // @[Math.scala 150:24:@34570.4]
  wire  x327_x7_1_reset; // @[Math.scala 150:24:@34570.4]
  wire [31:0] x327_x7_1_io_a; // @[Math.scala 150:24:@34570.4]
  wire [31:0] x327_x7_1_io_b; // @[Math.scala 150:24:@34570.4]
  wire  x327_x7_1_io_flow; // @[Math.scala 150:24:@34570.4]
  wire [31:0] x327_x7_1_io_result; // @[Math.scala 150:24:@34570.4]
  wire  x328_x8_1_clock; // @[Math.scala 150:24:@34580.4]
  wire  x328_x8_1_reset; // @[Math.scala 150:24:@34580.4]
  wire [31:0] x328_x8_1_io_a; // @[Math.scala 150:24:@34580.4]
  wire [31:0] x328_x8_1_io_b; // @[Math.scala 150:24:@34580.4]
  wire  x328_x8_1_io_flow; // @[Math.scala 150:24:@34580.4]
  wire [31:0] x328_x8_1_io_result; // @[Math.scala 150:24:@34580.4]
  wire  x329_x7_1_clock; // @[Math.scala 150:24:@34590.4]
  wire  x329_x7_1_reset; // @[Math.scala 150:24:@34590.4]
  wire [31:0] x329_x7_1_io_a; // @[Math.scala 150:24:@34590.4]
  wire [31:0] x329_x7_1_io_b; // @[Math.scala 150:24:@34590.4]
  wire  x329_x7_1_io_flow; // @[Math.scala 150:24:@34590.4]
  wire [31:0] x329_x7_1_io_result; // @[Math.scala 150:24:@34590.4]
  wire  x330_x8_1_clock; // @[Math.scala 150:24:@34600.4]
  wire  x330_x8_1_reset; // @[Math.scala 150:24:@34600.4]
  wire [31:0] x330_x8_1_io_a; // @[Math.scala 150:24:@34600.4]
  wire [31:0] x330_x8_1_io_b; // @[Math.scala 150:24:@34600.4]
  wire  x330_x8_1_io_flow; // @[Math.scala 150:24:@34600.4]
  wire [31:0] x330_x8_1_io_result; // @[Math.scala 150:24:@34600.4]
  wire  x331_x7_1_clock; // @[Math.scala 150:24:@34610.4]
  wire  x331_x7_1_reset; // @[Math.scala 150:24:@34610.4]
  wire [31:0] x331_x7_1_io_a; // @[Math.scala 150:24:@34610.4]
  wire [31:0] x331_x7_1_io_b; // @[Math.scala 150:24:@34610.4]
  wire  x331_x7_1_io_flow; // @[Math.scala 150:24:@34610.4]
  wire [31:0] x331_x7_1_io_result; // @[Math.scala 150:24:@34610.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@34620.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@34620.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@34620.4]
  wire [31:0] RetimeWrapper_72_io_in; // @[package.scala 93:22:@34620.4]
  wire [31:0] RetimeWrapper_72_io_out; // @[package.scala 93:22:@34620.4]
  wire  x332_sum_1_clock; // @[Math.scala 150:24:@34629.4]
  wire  x332_sum_1_reset; // @[Math.scala 150:24:@34629.4]
  wire [31:0] x332_sum_1_io_a; // @[Math.scala 150:24:@34629.4]
  wire [31:0] x332_sum_1_io_b; // @[Math.scala 150:24:@34629.4]
  wire  x332_sum_1_io_flow; // @[Math.scala 150:24:@34629.4]
  wire [31:0] x332_sum_1_io_result; // @[Math.scala 150:24:@34629.4]
  wire [31:0] x333_1_io_b; // @[Math.scala 720:24:@34639.4]
  wire [31:0] x333_1_io_result; // @[Math.scala 720:24:@34639.4]
  wire  x334_mul_1_clock; // @[Math.scala 262:24:@34650.4]
  wire [31:0] x334_mul_1_io_a; // @[Math.scala 262:24:@34650.4]
  wire [31:0] x334_mul_1_io_b; // @[Math.scala 262:24:@34650.4]
  wire  x334_mul_1_io_flow; // @[Math.scala 262:24:@34650.4]
  wire [31:0] x334_mul_1_io_result; // @[Math.scala 262:24:@34650.4]
  wire [31:0] x335_1_io_b; // @[Math.scala 720:24:@34660.4]
  wire [31:0] x335_1_io_result; // @[Math.scala 720:24:@34660.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@34669.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@34669.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@34669.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@34669.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@34669.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@34678.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@34678.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@34678.4]
  wire [31:0] RetimeWrapper_74_io_in; // @[package.scala 93:22:@34678.4]
  wire [31:0] RetimeWrapper_74_io_out; // @[package.scala 93:22:@34678.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@34687.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@34687.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@34687.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@34687.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@34687.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@34696.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@34696.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@34696.4]
  wire [31:0] RetimeWrapper_76_io_in; // @[package.scala 93:22:@34696.4]
  wire [31:0] RetimeWrapper_76_io_out; // @[package.scala 93:22:@34696.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@34705.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@34705.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@34705.4]
  wire [31:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@34705.4]
  wire [31:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@34705.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@34714.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@34714.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@34714.4]
  wire [31:0] RetimeWrapper_78_io_in; // @[package.scala 93:22:@34714.4]
  wire [31:0] RetimeWrapper_78_io_out; // @[package.scala 93:22:@34714.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@34725.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@34725.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@34725.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@34725.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@34725.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@34746.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@34746.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@34746.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@34746.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@34746.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@34755.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@34755.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@34755.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@34755.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@34755.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@34764.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@34764.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@34764.4]
  wire [31:0] RetimeWrapper_82_io_in; // @[package.scala 93:22:@34764.4]
  wire [31:0] RetimeWrapper_82_io_out; // @[package.scala 93:22:@34764.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@34773.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@34773.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@34773.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@34773.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@34773.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@34782.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@34782.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@34782.4]
  wire [31:0] RetimeWrapper_84_io_in; // @[package.scala 93:22:@34782.4]
  wire [31:0] RetimeWrapper_84_io_out; // @[package.scala 93:22:@34782.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@34791.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@34791.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@34791.4]
  wire [31:0] RetimeWrapper_85_io_in; // @[package.scala 93:22:@34791.4]
  wire [31:0] RetimeWrapper_85_io_out; // @[package.scala 93:22:@34791.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@34803.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@34803.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@34803.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@34803.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@34803.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@34824.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@34824.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@34824.4]
  wire [31:0] RetimeWrapper_87_io_in; // @[package.scala 93:22:@34824.4]
  wire [31:0] RetimeWrapper_87_io_out; // @[package.scala 93:22:@34824.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@34833.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@34833.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@34833.4]
  wire [31:0] RetimeWrapper_88_io_in; // @[package.scala 93:22:@34833.4]
  wire [31:0] RetimeWrapper_88_io_out; // @[package.scala 93:22:@34833.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@34842.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@34842.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@34842.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@34842.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@34842.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@34854.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@34854.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@34854.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@34854.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@34854.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@34875.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@34875.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@34875.4]
  wire [31:0] RetimeWrapper_91_io_in; // @[package.scala 93:22:@34875.4]
  wire [31:0] RetimeWrapper_91_io_out; // @[package.scala 93:22:@34875.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@34884.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@34884.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@34884.4]
  wire [31:0] RetimeWrapper_92_io_in; // @[package.scala 93:22:@34884.4]
  wire [31:0] RetimeWrapper_92_io_out; // @[package.scala 93:22:@34884.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@34893.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@34893.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@34893.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@34893.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@34893.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@34905.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@34905.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@34905.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@34905.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@34905.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@34926.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@34926.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@34926.4]
  wire [31:0] RetimeWrapper_95_io_in; // @[package.scala 93:22:@34926.4]
  wire [31:0] RetimeWrapper_95_io_out; // @[package.scala 93:22:@34926.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@34935.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@34935.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@34935.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@34935.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@34935.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@34947.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@34947.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@34947.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@34947.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@34947.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@34970.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@34970.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@34970.4]
  wire [32:0] RetimeWrapper_98_io_in; // @[package.scala 93:22:@34970.4]
  wire [32:0] RetimeWrapper_98_io_out; // @[package.scala 93:22:@34970.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@34982.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@34982.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@34982.4]
  wire [33:0] RetimeWrapper_99_io_in; // @[package.scala 93:22:@34982.4]
  wire [33:0] RetimeWrapper_99_io_out; // @[package.scala 93:22:@34982.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@34992.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@34992.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@34992.4]
  wire [31:0] RetimeWrapper_100_io_in; // @[package.scala 93:22:@34992.4]
  wire [31:0] RetimeWrapper_100_io_out; // @[package.scala 93:22:@34992.4]
  wire  x349_x9_1_clock; // @[Math.scala 150:24:@35001.4]
  wire  x349_x9_1_reset; // @[Math.scala 150:24:@35001.4]
  wire [31:0] x349_x9_1_io_a; // @[Math.scala 150:24:@35001.4]
  wire [31:0] x349_x9_1_io_b; // @[Math.scala 150:24:@35001.4]
  wire  x349_x9_1_io_flow; // @[Math.scala 150:24:@35001.4]
  wire [31:0] x349_x9_1_io_result; // @[Math.scala 150:24:@35001.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@35011.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@35011.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@35011.4]
  wire [31:0] RetimeWrapper_101_io_in; // @[package.scala 93:22:@35011.4]
  wire [31:0] RetimeWrapper_101_io_out; // @[package.scala 93:22:@35011.4]
  wire  x350_x10_1_clock; // @[Math.scala 150:24:@35022.4]
  wire  x350_x10_1_reset; // @[Math.scala 150:24:@35022.4]
  wire [31:0] x350_x10_1_io_a; // @[Math.scala 150:24:@35022.4]
  wire [31:0] x350_x10_1_io_b; // @[Math.scala 150:24:@35022.4]
  wire  x350_x10_1_io_flow; // @[Math.scala 150:24:@35022.4]
  wire [31:0] x350_x10_1_io_result; // @[Math.scala 150:24:@35022.4]
  wire  x351_sum_1_clock; // @[Math.scala 150:24:@35032.4]
  wire  x351_sum_1_reset; // @[Math.scala 150:24:@35032.4]
  wire [31:0] x351_sum_1_io_a; // @[Math.scala 150:24:@35032.4]
  wire [31:0] x351_sum_1_io_b; // @[Math.scala 150:24:@35032.4]
  wire  x351_sum_1_io_flow; // @[Math.scala 150:24:@35032.4]
  wire [31:0] x351_sum_1_io_result; // @[Math.scala 150:24:@35032.4]
  wire [31:0] x352_1_io_b; // @[Math.scala 720:24:@35042.4]
  wire [31:0] x352_1_io_result; // @[Math.scala 720:24:@35042.4]
  wire  x353_mul_1_clock; // @[Math.scala 262:24:@35053.4]
  wire [31:0] x353_mul_1_io_a; // @[Math.scala 262:24:@35053.4]
  wire [31:0] x353_mul_1_io_b; // @[Math.scala 262:24:@35053.4]
  wire  x353_mul_1_io_flow; // @[Math.scala 262:24:@35053.4]
  wire [31:0] x353_mul_1_io_result; // @[Math.scala 262:24:@35053.4]
  wire [31:0] x354_1_io_b; // @[Math.scala 720:24:@35063.4]
  wire [31:0] x354_1_io_result; // @[Math.scala 720:24:@35063.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@35076.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@35076.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@35076.4]
  wire [31:0] RetimeWrapper_102_io_in; // @[package.scala 93:22:@35076.4]
  wire [31:0] RetimeWrapper_102_io_out; // @[package.scala 93:22:@35076.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@35085.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@35085.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@35085.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@35085.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@35085.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@35094.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@35094.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@35094.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@35094.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@35094.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@35103.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@35103.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@35103.4]
  wire  RetimeWrapper_105_io_in; // @[package.scala 93:22:@35103.4]
  wire  RetimeWrapper_105_io_out; // @[package.scala 93:22:@35103.4]
  wire  b237; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 62:18:@32404.4]
  wire  b238; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 63:18:@32405.4]
  wire  _T_205; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 67:30:@32407.4]
  wire  _T_206; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 67:37:@32408.4]
  wire  _T_210; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 69:76:@32413.4]
  wire  _T_211; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 69:62:@32414.4]
  wire  _T_213; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 69:101:@32415.4]
  wire [31:0] b235_number; // @[Math.scala 723:22:@32389.4 Math.scala 724:14:@32390.4]
  wire [31:0] _T_242; // @[Math.scala 406:49:@32542.4]
  wire [31:0] _T_244; // @[Math.scala 406:56:@32544.4]
  wire [31:0] _T_245; // @[Math.scala 406:56:@32545.4]
  wire [31:0] x412_number; // @[implicits.scala 133:21:@32546.4]
  wire [31:0] _T_255; // @[Math.scala 406:49:@32555.4]
  wire [31:0] _T_257; // @[Math.scala 406:56:@32557.4]
  wire [31:0] _T_258; // @[Math.scala 406:56:@32558.4]
  wire [31:0] b236_number; // @[Math.scala 723:22:@32401.4 Math.scala 724:14:@32402.4]
  wire  _T_262; // @[FixedPoint.scala 50:25:@32564.4]
  wire [15:0] _T_266; // @[Bitwise.scala 72:12:@32566.4]
  wire [15:0] _T_267; // @[FixedPoint.scala 18:52:@32567.4]
  wire  _T_273; // @[Math.scala 451:55:@32569.4]
  wire [15:0] _T_274; // @[FixedPoint.scala 18:52:@32570.4]
  wire  _T_280; // @[Math.scala 451:110:@32572.4]
  wire  _T_281; // @[Math.scala 451:94:@32573.4]
  wire [31:0] _T_283; // @[Cat.scala 30:58:@32575.4]
  wire [31:0] _T_293; // @[Math.scala 406:49:@32583.4]
  wire [31:0] _T_295; // @[Math.scala 406:56:@32585.4]
  wire [31:0] _T_296; // @[Math.scala 406:56:@32586.4]
  wire [31:0] x416_sum_number; // @[Math.scala 154:22:@32597.4 Math.scala 155:14:@32598.4]
  wire  _T_303; // @[FixedPoint.scala 50:25:@32602.4]
  wire [7:0] _T_307; // @[Bitwise.scala 72:12:@32604.4]
  wire [23:0] _T_308; // @[FixedPoint.scala 18:52:@32605.4]
  wire  _T_314; // @[Math.scala 451:55:@32607.4]
  wire [7:0] _T_315; // @[FixedPoint.scala 18:52:@32608.4]
  wire  _T_321; // @[Math.scala 451:110:@32610.4]
  wire  _T_322; // @[Math.scala 451:94:@32611.4]
  wire [31:0] _T_324; // @[Cat.scala 30:58:@32613.4]
  wire [31:0] _T_334; // @[Math.scala 406:49:@32621.4]
  wire [31:0] _T_336; // @[Math.scala 406:56:@32623.4]
  wire [31:0] _T_337; // @[Math.scala 406:56:@32624.4]
  wire [31:0] x419_sum_number; // @[Math.scala 154:22:@32635.4 Math.scala 155:14:@32636.4]
  wire  _T_344; // @[FixedPoint.scala 50:25:@32640.4]
  wire [3:0] _T_348; // @[Bitwise.scala 72:12:@32642.4]
  wire [27:0] _T_349; // @[FixedPoint.scala 18:52:@32643.4]
  wire  _T_355; // @[Math.scala 451:55:@32645.4]
  wire [3:0] _T_356; // @[FixedPoint.scala 18:52:@32646.4]
  wire  _T_362; // @[Math.scala 451:110:@32648.4]
  wire  _T_363; // @[Math.scala 451:94:@32649.4]
  wire [31:0] _T_365; // @[Cat.scala 30:58:@32651.4]
  wire [31:0] _T_375; // @[Math.scala 406:49:@32659.4]
  wire [31:0] _T_377; // @[Math.scala 406:56:@32661.4]
  wire [31:0] _T_378; // @[Math.scala 406:56:@32662.4]
  wire [31:0] x422_sum_number; // @[Math.scala 154:22:@32673.4 Math.scala 155:14:@32674.4]
  wire  _T_385; // @[FixedPoint.scala 50:25:@32678.4]
  wire [1:0] _T_389; // @[Bitwise.scala 72:12:@32680.4]
  wire [29:0] _T_390; // @[FixedPoint.scala 18:52:@32681.4]
  wire  _T_396; // @[Math.scala 451:55:@32683.4]
  wire [1:0] _T_397; // @[FixedPoint.scala 18:52:@32684.4]
  wire  _T_403; // @[Math.scala 451:110:@32686.4]
  wire  _T_404; // @[Math.scala 451:94:@32687.4]
  wire [31:0] _T_406; // @[Cat.scala 30:58:@32689.4]
  wire [31:0] _T_416; // @[Math.scala 406:49:@32697.4]
  wire [31:0] _T_418; // @[Math.scala 406:56:@32699.4]
  wire [31:0] _T_419; // @[Math.scala 406:56:@32700.4]
  wire [31:0] x425_sum_number; // @[Math.scala 154:22:@32711.4 Math.scala 155:14:@32712.4]
  wire  _T_426; // @[FixedPoint.scala 50:25:@32716.4]
  wire [1:0] _T_430; // @[Bitwise.scala 72:12:@32718.4]
  wire [29:0] _T_431; // @[FixedPoint.scala 18:52:@32719.4]
  wire  _T_437; // @[Math.scala 451:55:@32721.4]
  wire [1:0] _T_438; // @[FixedPoint.scala 18:52:@32722.4]
  wire  _T_444; // @[Math.scala 451:110:@32724.4]
  wire  _T_445; // @[Math.scala 451:94:@32725.4]
  wire [31:0] _T_449; // @[package.scala 96:25:@32733.4 package.scala 96:25:@32734.4]
  wire [31:0] _T_459; // @[Math.scala 406:49:@32742.4]
  wire [31:0] _T_461; // @[Math.scala 406:56:@32744.4]
  wire [31:0] _T_462; // @[Math.scala 406:56:@32745.4]
  wire [31:0] _T_466; // @[package.scala 96:25:@32753.4]
  wire [31:0] x428_sum_number; // @[Math.scala 154:22:@32765.4 Math.scala 155:14:@32766.4]
  wire  _T_473; // @[FixedPoint.scala 50:25:@32770.4]
  wire [1:0] _T_477; // @[Bitwise.scala 72:12:@32772.4]
  wire [29:0] _T_478; // @[FixedPoint.scala 18:52:@32773.4]
  wire  _T_484; // @[Math.scala 451:55:@32775.4]
  wire [1:0] _T_485; // @[FixedPoint.scala 18:52:@32776.4]
  wire  _T_491; // @[Math.scala 451:110:@32778.4]
  wire  _T_492; // @[Math.scala 451:94:@32779.4]
  wire [31:0] _T_494; // @[Cat.scala 30:58:@32781.4]
  wire [31:0] _T_504; // @[Math.scala 406:49:@32789.4]
  wire [31:0] _T_506; // @[Math.scala 406:56:@32791.4]
  wire [31:0] _T_507; // @[Math.scala 406:56:@32792.4]
  wire [31:0] x431_sum_number; // @[Math.scala 154:22:@32803.4 Math.scala 155:14:@32804.4]
  wire [31:0] _T_517; // @[Math.scala 476:37:@32809.4]
  wire  x499_x432_D1; // @[package.scala 96:25:@32838.4 package.scala 96:25:@32839.4]
  wire [31:0] x501_x431_sum_D1_number; // @[package.scala 96:25:@32856.4 package.scala 96:25:@32857.4]
  wire [31:0] x434_sub_number; // @[Math.scala 195:22:@32829.4 Math.scala 196:14:@32830.4]
  wire  _T_548; // @[FixedPoint.scala 50:25:@32864.4]
  wire [1:0] _T_552; // @[Bitwise.scala 72:12:@32866.4]
  wire [29:0] _T_553; // @[FixedPoint.scala 18:52:@32867.4]
  wire  _T_559; // @[Math.scala 451:55:@32869.4]
  wire [1:0] _T_560; // @[FixedPoint.scala 18:52:@32870.4]
  wire  _T_566; // @[Math.scala 451:110:@32872.4]
  wire  _T_567; // @[Math.scala 451:94:@32873.4]
  wire [31:0] _T_569; // @[Cat.scala 30:58:@32875.4]
  wire [31:0] x248_1_number; // @[Math.scala 454:20:@32876.4]
  wire [40:0] _GEN_0; // @[Math.scala 461:32:@32881.4]
  wire [40:0] _T_574; // @[Math.scala 461:32:@32881.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@32886.4]
  wire [38:0] _T_577; // @[Math.scala 461:32:@32886.4]
  wire  _T_610; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 164:101:@32975.4]
  wire  _T_614; // @[package.scala 96:25:@32983.4 package.scala 96:25:@32984.4]
  wire  _T_616; // @[implicits.scala 55:10:@32985.4]
  wire  _T_617; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 164:118:@32986.4]
  wire  _T_619; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 164:207:@32988.4]
  wire  _T_620; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 164:226:@32989.4]
  wire  x505_b237_D21; // @[package.scala 96:25:@32954.4 package.scala 96:25:@32955.4]
  wire  _T_621; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 164:252:@32990.4]
  wire  x503_b238_D21; // @[package.scala 96:25:@32936.4 package.scala 96:25:@32937.4]
  wire [31:0] x508_b235_D23_number; // @[package.scala 96:25:@33004.4 package.scala 96:25:@33005.4]
  wire [31:0] _T_633; // @[Math.scala 476:37:@33012.4]
  wire [31:0] x509_b236_D23_number; // @[package.scala 96:25:@33029.4 package.scala 96:25:@33030.4]
  wire [31:0] _T_646; // @[Math.scala 476:37:@33035.4]
  wire  x254; // @[package.scala 96:25:@33020.4 package.scala 96:25:@33021.4]
  wire  x255; // @[package.scala 96:25:@33043.4 package.scala 96:25:@33044.4]
  wire  x256; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 183:24:@33047.4]
  wire  _T_684; // @[package.scala 96:25:@33115.4 package.scala 96:25:@33116.4]
  wire  _T_686; // @[implicits.scala 55:10:@33117.4]
  wire  _T_687; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 202:194:@33118.4]
  wire  x510_x257_D21; // @[package.scala 96:25:@33058.4 package.scala 96:25:@33059.4]
  wire  _T_688; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 202:283:@33119.4]
  wire  x513_b237_D45; // @[package.scala 96:25:@33085.4 package.scala 96:25:@33086.4]
  wire  _T_689; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 202:291:@33120.4]
  wire  x511_b238_D45; // @[package.scala 96:25:@33067.4 package.scala 96:25:@33068.4]
  wire [31:0] x260_rdcol_number; // @[Math.scala 195:22:@33139.4 Math.scala 196:14:@33140.4]
  wire [31:0] _T_704; // @[Math.scala 476:37:@33145.4]
  wire  x516_x254_D1; // @[package.scala 96:25:@33162.4 package.scala 96:25:@33163.4]
  wire  x261; // @[package.scala 96:25:@33153.4 package.scala 96:25:@33154.4]
  wire  x262; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 212:24:@33166.4]
  wire  _T_718; // @[FixedPoint.scala 50:25:@33173.4]
  wire [15:0] _T_722; // @[Bitwise.scala 72:12:@33175.4]
  wire [15:0] _T_723; // @[FixedPoint.scala 18:52:@33176.4]
  wire  _T_729; // @[Math.scala 451:55:@33178.4]
  wire [15:0] _T_730; // @[FixedPoint.scala 18:52:@33179.4]
  wire  _T_736; // @[Math.scala 451:110:@33181.4]
  wire  _T_737; // @[Math.scala 451:94:@33182.4]
  wire [31:0] _T_739; // @[Cat.scala 30:58:@33184.4]
  wire [31:0] _T_751; // @[Math.scala 406:56:@33194.4]
  wire [31:0] _T_752; // @[Math.scala 406:56:@33195.4]
  wire [31:0] x441_sum_number; // @[Math.scala 154:22:@33206.4 Math.scala 155:14:@33207.4]
  wire  _T_759; // @[FixedPoint.scala 50:25:@33211.4]
  wire [7:0] _T_763; // @[Bitwise.scala 72:12:@33213.4]
  wire [23:0] _T_764; // @[FixedPoint.scala 18:52:@33214.4]
  wire  _T_770; // @[Math.scala 451:55:@33216.4]
  wire [7:0] _T_771; // @[FixedPoint.scala 18:52:@33217.4]
  wire  _T_777; // @[Math.scala 451:110:@33219.4]
  wire  _T_778; // @[Math.scala 451:94:@33220.4]
  wire [31:0] _T_782; // @[package.scala 96:25:@33228.4 package.scala 96:25:@33229.4]
  wire [31:0] _T_792; // @[Math.scala 406:49:@33237.4]
  wire [31:0] _T_794; // @[Math.scala 406:56:@33239.4]
  wire [31:0] _T_795; // @[Math.scala 406:56:@33240.4]
  wire [31:0] _T_799; // @[package.scala 96:25:@33248.4]
  wire [31:0] x444_sum_number; // @[Math.scala 154:22:@33260.4 Math.scala 155:14:@33261.4]
  wire  _T_806; // @[FixedPoint.scala 50:25:@33265.4]
  wire [3:0] _T_810; // @[Bitwise.scala 72:12:@33267.4]
  wire [27:0] _T_811; // @[FixedPoint.scala 18:52:@33268.4]
  wire  _T_817; // @[Math.scala 451:55:@33270.4]
  wire [3:0] _T_818; // @[FixedPoint.scala 18:52:@33271.4]
  wire  _T_824; // @[Math.scala 451:110:@33273.4]
  wire  _T_825; // @[Math.scala 451:94:@33274.4]
  wire [31:0] _T_827; // @[Cat.scala 30:58:@33276.4]
  wire [31:0] _T_837; // @[Math.scala 406:49:@33284.4]
  wire [31:0] _T_839; // @[Math.scala 406:56:@33286.4]
  wire [31:0] _T_840; // @[Math.scala 406:56:@33287.4]
  wire [31:0] x447_sum_number; // @[Math.scala 154:22:@33298.4 Math.scala 155:14:@33299.4]
  wire  _T_847; // @[FixedPoint.scala 50:25:@33303.4]
  wire [1:0] _T_851; // @[Bitwise.scala 72:12:@33305.4]
  wire [29:0] _T_852; // @[FixedPoint.scala 18:52:@33306.4]
  wire  _T_858; // @[Math.scala 451:55:@33308.4]
  wire [1:0] _T_859; // @[FixedPoint.scala 18:52:@33309.4]
  wire  _T_865; // @[Math.scala 451:110:@33311.4]
  wire  _T_866; // @[Math.scala 451:94:@33312.4]
  wire [31:0] _T_868; // @[Cat.scala 30:58:@33314.4]
  wire [31:0] _T_878; // @[Math.scala 406:49:@33322.4]
  wire [31:0] _T_880; // @[Math.scala 406:56:@33324.4]
  wire [31:0] _T_881; // @[Math.scala 406:56:@33325.4]
  wire [31:0] x450_sum_number; // @[Math.scala 154:22:@33336.4 Math.scala 155:14:@33337.4]
  wire  _T_888; // @[FixedPoint.scala 50:25:@33341.4]
  wire [1:0] _T_892; // @[Bitwise.scala 72:12:@33343.4]
  wire [29:0] _T_893; // @[FixedPoint.scala 18:52:@33344.4]
  wire  _T_899; // @[Math.scala 451:55:@33346.4]
  wire [1:0] _T_900; // @[FixedPoint.scala 18:52:@33347.4]
  wire  _T_906; // @[Math.scala 451:110:@33349.4]
  wire  _T_907; // @[Math.scala 451:94:@33350.4]
  wire [31:0] _T_909; // @[Cat.scala 30:58:@33352.4]
  wire [31:0] _T_919; // @[Math.scala 406:49:@33360.4]
  wire [31:0] _T_921; // @[Math.scala 406:56:@33362.4]
  wire [31:0] _T_922; // @[Math.scala 406:56:@33363.4]
  wire [31:0] x453_sum_number; // @[Math.scala 154:22:@33374.4 Math.scala 155:14:@33375.4]
  wire  _T_929; // @[FixedPoint.scala 50:25:@33379.4]
  wire [1:0] _T_933; // @[Bitwise.scala 72:12:@33381.4]
  wire [29:0] _T_934; // @[FixedPoint.scala 18:52:@33382.4]
  wire  _T_940; // @[Math.scala 451:55:@33384.4]
  wire [1:0] _T_941; // @[FixedPoint.scala 18:52:@33385.4]
  wire  _T_947; // @[Math.scala 451:110:@33387.4]
  wire  _T_948; // @[Math.scala 451:94:@33388.4]
  wire [31:0] _T_950; // @[Cat.scala 30:58:@33390.4]
  wire [31:0] _T_960; // @[Math.scala 406:49:@33398.4]
  wire [31:0] _T_962; // @[Math.scala 406:56:@33400.4]
  wire [31:0] _T_963; // @[Math.scala 406:56:@33401.4]
  wire [31:0] x456_sum_number; // @[Math.scala 154:22:@33412.4 Math.scala 155:14:@33413.4]
  wire [31:0] _T_973; // @[Math.scala 476:37:@33418.4]
  wire  x457; // @[package.scala 96:25:@33426.4 package.scala 96:25:@33427.4]
  wire [31:0] x517_x456_sum_D1_number; // @[package.scala 96:25:@33461.4 package.scala 96:25:@33462.4]
  wire [31:0] x459_sub_number; // @[Math.scala 195:22:@33452.4 Math.scala 196:14:@33453.4]
  wire  _T_1030; // @[package.scala 96:25:@33525.4 package.scala 96:25:@33526.4]
  wire  _T_1032; // @[implicits.scala 55:10:@33527.4]
  wire  _T_1033; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 275:194:@33528.4]
  wire  x520_x263_D20; // @[package.scala 96:25:@33513.4 package.scala 96:25:@33514.4]
  wire  _T_1034; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 275:283:@33529.4]
  wire  _T_1035; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 275:291:@33530.4]
  wire [31:0] x269_rdcol_number; // @[Math.scala 195:22:@33549.4 Math.scala 196:14:@33550.4]
  wire [31:0] _T_1052; // @[Math.scala 476:37:@33557.4]
  wire  x270; // @[package.scala 96:25:@33565.4 package.scala 96:25:@33566.4]
  wire  x271; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 291:59:@33569.4]
  wire  _T_1063; // @[FixedPoint.scala 50:25:@33576.4]
  wire [15:0] _T_1067; // @[Bitwise.scala 72:12:@33578.4]
  wire [15:0] _T_1068; // @[FixedPoint.scala 18:52:@33579.4]
  wire  _T_1074; // @[Math.scala 451:55:@33581.4]
  wire [15:0] _T_1075; // @[FixedPoint.scala 18:52:@33582.4]
  wire  _T_1081; // @[Math.scala 451:110:@33584.4]
  wire  _T_1082; // @[Math.scala 451:94:@33585.4]
  wire [31:0] _T_1084; // @[Cat.scala 30:58:@33587.4]
  wire [31:0] _T_1096; // @[Math.scala 406:56:@33597.4]
  wire [31:0] _T_1097; // @[Math.scala 406:56:@33598.4]
  wire [31:0] x463_sum_number; // @[Math.scala 154:22:@33609.4 Math.scala 155:14:@33610.4]
  wire  _T_1104; // @[FixedPoint.scala 50:25:@33614.4]
  wire [7:0] _T_1108; // @[Bitwise.scala 72:12:@33616.4]
  wire [23:0] _T_1109; // @[FixedPoint.scala 18:52:@33617.4]
  wire  _T_1115; // @[Math.scala 451:55:@33619.4]
  wire [7:0] _T_1116; // @[FixedPoint.scala 18:52:@33620.4]
  wire  _T_1122; // @[Math.scala 451:110:@33622.4]
  wire  _T_1123; // @[Math.scala 451:94:@33623.4]
  wire [31:0] _T_1127; // @[package.scala 96:25:@33631.4 package.scala 96:25:@33632.4]
  wire [31:0] _T_1137; // @[Math.scala 406:49:@33640.4]
  wire [31:0] _T_1139; // @[Math.scala 406:56:@33642.4]
  wire [31:0] _T_1140; // @[Math.scala 406:56:@33643.4]
  wire [31:0] _T_1144; // @[package.scala 96:25:@33651.4]
  wire [31:0] x466_sum_number; // @[Math.scala 154:22:@33663.4 Math.scala 155:14:@33664.4]
  wire  _T_1151; // @[FixedPoint.scala 50:25:@33668.4]
  wire [3:0] _T_1155; // @[Bitwise.scala 72:12:@33670.4]
  wire [27:0] _T_1156; // @[FixedPoint.scala 18:52:@33671.4]
  wire  _T_1162; // @[Math.scala 451:55:@33673.4]
  wire [3:0] _T_1163; // @[FixedPoint.scala 18:52:@33674.4]
  wire  _T_1169; // @[Math.scala 451:110:@33676.4]
  wire  _T_1170; // @[Math.scala 451:94:@33677.4]
  wire [31:0] _T_1172; // @[Cat.scala 30:58:@33679.4]
  wire [31:0] _T_1182; // @[Math.scala 406:49:@33687.4]
  wire [31:0] _T_1184; // @[Math.scala 406:56:@33689.4]
  wire [31:0] _T_1185; // @[Math.scala 406:56:@33690.4]
  wire [31:0] x469_sum_number; // @[Math.scala 154:22:@33701.4 Math.scala 155:14:@33702.4]
  wire  _T_1192; // @[FixedPoint.scala 50:25:@33706.4]
  wire [1:0] _T_1196; // @[Bitwise.scala 72:12:@33708.4]
  wire [29:0] _T_1197; // @[FixedPoint.scala 18:52:@33709.4]
  wire  _T_1203; // @[Math.scala 451:55:@33711.4]
  wire [1:0] _T_1204; // @[FixedPoint.scala 18:52:@33712.4]
  wire  _T_1210; // @[Math.scala 451:110:@33714.4]
  wire  _T_1211; // @[Math.scala 451:94:@33715.4]
  wire [31:0] _T_1213; // @[Cat.scala 30:58:@33717.4]
  wire [31:0] _T_1223; // @[Math.scala 406:49:@33725.4]
  wire [31:0] _T_1225; // @[Math.scala 406:56:@33727.4]
  wire [31:0] _T_1226; // @[Math.scala 406:56:@33728.4]
  wire [31:0] x472_sum_number; // @[Math.scala 154:22:@33739.4 Math.scala 155:14:@33740.4]
  wire  _T_1233; // @[FixedPoint.scala 50:25:@33744.4]
  wire [1:0] _T_1237; // @[Bitwise.scala 72:12:@33746.4]
  wire [29:0] _T_1238; // @[FixedPoint.scala 18:52:@33747.4]
  wire  _T_1244; // @[Math.scala 451:55:@33749.4]
  wire [1:0] _T_1245; // @[FixedPoint.scala 18:52:@33750.4]
  wire  _T_1251; // @[Math.scala 451:110:@33752.4]
  wire  _T_1252; // @[Math.scala 451:94:@33753.4]
  wire [31:0] _T_1254; // @[Cat.scala 30:58:@33755.4]
  wire [31:0] _T_1264; // @[Math.scala 406:49:@33763.4]
  wire [31:0] _T_1266; // @[Math.scala 406:56:@33765.4]
  wire [31:0] _T_1267; // @[Math.scala 406:56:@33766.4]
  wire [31:0] x475_sum_number; // @[Math.scala 154:22:@33777.4 Math.scala 155:14:@33778.4]
  wire  _T_1274; // @[FixedPoint.scala 50:25:@33782.4]
  wire [1:0] _T_1278; // @[Bitwise.scala 72:12:@33784.4]
  wire [29:0] _T_1279; // @[FixedPoint.scala 18:52:@33785.4]
  wire  _T_1285; // @[Math.scala 451:55:@33787.4]
  wire [1:0] _T_1286; // @[FixedPoint.scala 18:52:@33788.4]
  wire  _T_1292; // @[Math.scala 451:110:@33790.4]
  wire  _T_1293; // @[Math.scala 451:94:@33791.4]
  wire [31:0] _T_1295; // @[Cat.scala 30:58:@33793.4]
  wire [31:0] _T_1305; // @[Math.scala 406:49:@33801.4]
  wire [31:0] _T_1307; // @[Math.scala 406:56:@33803.4]
  wire [31:0] _T_1308; // @[Math.scala 406:56:@33804.4]
  wire [31:0] x478_sum_number; // @[Math.scala 154:22:@33815.4 Math.scala 155:14:@33816.4]
  wire [31:0] _T_1318; // @[Math.scala 476:37:@33821.4]
  wire  x479; // @[package.scala 96:25:@33829.4 package.scala 96:25:@33830.4]
  wire [31:0] x521_x478_sum_D1_number; // @[package.scala 96:25:@33864.4 package.scala 96:25:@33865.4]
  wire [31:0] x481_sub_number; // @[Math.scala 195:22:@33855.4 Math.scala 196:14:@33856.4]
  wire  _T_1372; // @[package.scala 96:25:@33919.4 package.scala 96:25:@33920.4]
  wire  _T_1374; // @[implicits.scala 55:10:@33921.4]
  wire  _T_1375; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 352:194:@33922.4]
  wire  x523_x272_D20; // @[package.scala 96:25:@33907.4 package.scala 96:25:@33908.4]
  wire  _T_1376; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 352:283:@33923.4]
  wire  _T_1377; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 352:291:@33924.4]
  wire [31:0] x278_rdrow_number; // @[Math.scala 195:22:@33943.4 Math.scala 196:14:@33944.4]
  wire [31:0] _T_1394; // @[Math.scala 406:49:@33950.4]
  wire [31:0] _T_1396; // @[Math.scala 406:56:@33952.4]
  wire [31:0] _T_1397; // @[Math.scala 406:56:@33953.4]
  wire [31:0] x483_number; // @[implicits.scala 133:21:@33954.4]
  wire  x280; // @[package.scala 96:25:@33968.4 package.scala 96:25:@33969.4]
  wire  x524_x255_D1; // @[package.scala 96:25:@33977.4 package.scala 96:25:@33978.4]
  wire  x281; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 364:24:@33981.4]
  wire [31:0] _T_1423; // @[Math.scala 406:49:@33990.4]
  wire [31:0] _T_1425; // @[Math.scala 406:56:@33992.4]
  wire [31:0] _T_1426; // @[Math.scala 406:56:@33993.4]
  wire [31:0] _T_1430; // @[package.scala 96:25:@34001.4]
  wire  _T_1434; // @[FixedPoint.scala 50:25:@34008.4]
  wire [1:0] _T_1438; // @[Bitwise.scala 72:12:@34010.4]
  wire [29:0] _T_1439; // @[FixedPoint.scala 18:52:@34011.4]
  wire  _T_1445; // @[Math.scala 451:55:@34013.4]
  wire [1:0] _T_1446; // @[FixedPoint.scala 18:52:@34014.4]
  wire  _T_1452; // @[Math.scala 451:110:@34016.4]
  wire  _T_1453; // @[Math.scala 451:94:@34017.4]
  wire [31:0] _T_1457; // @[package.scala 96:25:@34025.4 package.scala 96:25:@34026.4]
  wire [31:0] x284_1_number; // @[Math.scala 454:20:@34027.4]
  wire [40:0] _GEN_2; // @[Math.scala 461:32:@34032.4]
  wire [40:0] _T_1462; // @[Math.scala 461:32:@34032.4]
  wire [38:0] _GEN_3; // @[Math.scala 461:32:@34037.4]
  wire [38:0] _T_1465; // @[Math.scala 461:32:@34037.4]
  wire  _T_1498; // @[package.scala 96:25:@34114.4 package.scala 96:25:@34115.4]
  wire  _T_1500; // @[implicits.scala 55:10:@34116.4]
  wire  _T_1501; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 399:194:@34117.4]
  wire  x529_x282_D20; // @[package.scala 96:25:@34102.4 package.scala 96:25:@34103.4]
  wire  _T_1502; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 399:283:@34118.4]
  wire  _T_1503; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 399:326:@34119.4]
  wire  x289; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 403:59:@34130.4]
  wire  _T_1532; // @[package.scala 96:25:@34174.4 package.scala 96:25:@34175.4]
  wire  _T_1534; // @[implicits.scala 55:10:@34176.4]
  wire  _T_1535; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 418:194:@34177.4]
  wire  x531_x290_D20; // @[package.scala 96:25:@34162.4 package.scala 96:25:@34163.4]
  wire  _T_1536; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 418:283:@34178.4]
  wire  _T_1537; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 418:291:@34179.4]
  wire  x294; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 422:59:@34190.4]
  wire  _T_1561; // @[package.scala 96:25:@34223.4 package.scala 96:25:@34224.4]
  wire  _T_1563; // @[implicits.scala 55:10:@34225.4]
  wire  _T_1564; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 433:194:@34226.4]
  wire  x532_x295_D20; // @[package.scala 96:25:@34211.4 package.scala 96:25:@34212.4]
  wire  _T_1565; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 433:283:@34227.4]
  wire  _T_1566; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 433:291:@34228.4]
  wire [31:0] x299_rdrow_number; // @[Math.scala 195:22:@34247.4 Math.scala 196:14:@34248.4]
  wire [31:0] _T_1583; // @[Math.scala 406:49:@34254.4]
  wire [31:0] _T_1585; // @[Math.scala 406:56:@34256.4]
  wire [31:0] _T_1586; // @[Math.scala 406:56:@34257.4]
  wire [31:0] x488_number; // @[implicits.scala 133:21:@34258.4]
  wire  x301; // @[package.scala 96:25:@34272.4 package.scala 96:25:@34273.4]
  wire  x302; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 443:24:@34276.4]
  wire [31:0] _T_1609; // @[Math.scala 406:49:@34285.4]
  wire [31:0] _T_1611; // @[Math.scala 406:56:@34287.4]
  wire [31:0] _T_1612; // @[Math.scala 406:56:@34288.4]
  wire [31:0] _T_1616; // @[package.scala 96:25:@34296.4]
  wire  _T_1620; // @[FixedPoint.scala 50:25:@34303.4]
  wire [1:0] _T_1624; // @[Bitwise.scala 72:12:@34305.4]
  wire [29:0] _T_1625; // @[FixedPoint.scala 18:52:@34306.4]
  wire  _T_1631; // @[Math.scala 451:55:@34308.4]
  wire [1:0] _T_1632; // @[FixedPoint.scala 18:52:@34309.4]
  wire  _T_1638; // @[Math.scala 451:110:@34311.4]
  wire  _T_1639; // @[Math.scala 451:94:@34312.4]
  wire [31:0] _T_1643; // @[package.scala 96:25:@34320.4 package.scala 96:25:@34321.4]
  wire [31:0] x305_1_number; // @[Math.scala 454:20:@34322.4]
  wire [40:0] _GEN_4; // @[Math.scala 461:32:@34327.4]
  wire [40:0] _T_1648; // @[Math.scala 461:32:@34327.4]
  wire [38:0] _GEN_5; // @[Math.scala 461:32:@34332.4]
  wire [38:0] _T_1651; // @[Math.scala 461:32:@34332.4]
  wire  _T_1681; // @[package.scala 96:25:@34400.4 package.scala 96:25:@34401.4]
  wire  _T_1683; // @[implicits.scala 55:10:@34402.4]
  wire  _T_1684; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 470:194:@34403.4]
  wire  x536_x303_D20; // @[package.scala 96:25:@34388.4 package.scala 96:25:@34389.4]
  wire  _T_1685; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 470:283:@34404.4]
  wire  _T_1686; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 470:291:@34405.4]
  wire  x310; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 474:24:@34416.4]
  wire  _T_1713; // @[package.scala 96:25:@34458.4 package.scala 96:25:@34459.4]
  wire  _T_1715; // @[implicits.scala 55:10:@34460.4]
  wire  _T_1716; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 487:194:@34461.4]
  wire  x538_x311_D20; // @[package.scala 96:25:@34446.4 package.scala 96:25:@34447.4]
  wire  _T_1717; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 487:283:@34462.4]
  wire  _T_1718; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 487:291:@34463.4]
  wire  x315; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 491:24:@34474.4]
  wire  _T_1742; // @[package.scala 96:25:@34507.4 package.scala 96:25:@34508.4]
  wire  _T_1744; // @[implicits.scala 55:10:@34509.4]
  wire  _T_1745; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 502:194:@34510.4]
  wire  x539_x316_D20; // @[package.scala 96:25:@34495.4 package.scala 96:25:@34496.4]
  wire  _T_1746; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 502:283:@34511.4]
  wire  _T_1747; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 502:291:@34512.4]
  wire [31:0] x267_rd_0_number; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 271:29:@33516.4 sm_x359_inr_Foreach_SAMPLER_BOX.scala 275:338:@33537.4]
  wire [32:0] _GEN_6; // @[Math.scala 461:32:@34524.4]
  wire [32:0] _T_1752; // @[Math.scala 461:32:@34524.4]
  wire [31:0] x287_rd_0_number; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 395:29:@34105.4 sm_x359_inr_Foreach_SAMPLER_BOX.scala 399:443:@34126.4]
  wire [32:0] _GEN_7; // @[Math.scala 461:32:@34529.4]
  wire [32:0] _T_1755; // @[Math.scala 461:32:@34529.4]
  wire [31:0] x292_rd_0_number; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 414:29:@34165.4 sm_x359_inr_Foreach_SAMPLER_BOX.scala 418:408:@34186.4]
  wire [33:0] _GEN_8; // @[Math.scala 461:32:@34534.4]
  wire [33:0] _T_1758; // @[Math.scala 461:32:@34534.4]
  wire [31:0] x297_rd_0_number; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 429:29:@34214.4 sm_x359_inr_Foreach_SAMPLER_BOX.scala 433:408:@34235.4]
  wire [32:0] _GEN_9; // @[Math.scala 461:32:@34539.4]
  wire [32:0] _T_1761; // @[Math.scala 461:32:@34539.4]
  wire [31:0] x313_rd_0_number; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 483:29:@34449.4 sm_x359_inr_Foreach_SAMPLER_BOX.scala 487:408:@34470.4]
  wire [32:0] _GEN_10; // @[Math.scala 461:32:@34546.4]
  wire [32:0] _T_1766; // @[Math.scala 461:32:@34546.4]
  wire  _T_1830; // @[package.scala 96:25:@34730.4 package.scala 96:25:@34731.4]
  wire  _T_1832; // @[implicits.scala 55:10:@34732.4]
  wire  _T_1833; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 564:167:@34733.4]
  wire  _T_1835; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 564:256:@34735.4]
  wire  _T_1836; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 564:275:@34736.4]
  wire  x543_b237_D58; // @[package.scala 96:25:@34692.4 package.scala 96:25:@34693.4]
  wire  _T_1837; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 564:301:@34737.4]
  wire  x541_b238_D58; // @[package.scala 96:25:@34674.4 package.scala 96:25:@34675.4]
  wire  _T_1868; // @[package.scala 96:25:@34808.4 package.scala 96:25:@34809.4]
  wire  _T_1870; // @[implicits.scala 55:10:@34810.4]
  wire  _T_1871; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 582:195:@34811.4]
  wire  x547_x257_D35; // @[package.scala 96:25:@34751.4 package.scala 96:25:@34752.4]
  wire  _T_1872; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 582:284:@34812.4]
  wire  x550_b237_D59; // @[package.scala 96:25:@34778.4 package.scala 96:25:@34779.4]
  wire  _T_1873; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 582:292:@34813.4]
  wire  x548_b238_D59; // @[package.scala 96:25:@34760.4 package.scala 96:25:@34761.4]
  wire  _T_1896; // @[package.scala 96:25:@34859.4 package.scala 96:25:@34860.4]
  wire  _T_1898; // @[implicits.scala 55:10:@34861.4]
  wire  _T_1899; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 595:195:@34862.4]
  wire  x555_x263_D34; // @[package.scala 96:25:@34847.4 package.scala 96:25:@34848.4]
  wire  _T_1900; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 595:284:@34863.4]
  wire  _T_1901; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 595:292:@34864.4]
  wire  _T_1924; // @[package.scala 96:25:@34910.4 package.scala 96:25:@34911.4]
  wire  _T_1926; // @[implicits.scala 55:10:@34912.4]
  wire  _T_1927; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 608:195:@34913.4]
  wire  x558_x282_D34; // @[package.scala 96:25:@34898.4 package.scala 96:25:@34899.4]
  wire  _T_1928; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 608:284:@34914.4]
  wire  _T_1929; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 608:292:@34915.4]
  wire  _T_1949; // @[package.scala 96:25:@34952.4 package.scala 96:25:@34953.4]
  wire  _T_1951; // @[implicits.scala 55:10:@34954.4]
  wire  _T_1952; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 619:195:@34955.4]
  wire  x560_x290_D34; // @[package.scala 96:25:@34940.4 package.scala 96:25:@34941.4]
  wire  _T_1953; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 619:284:@34956.4]
  wire  _T_1954; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 619:292:@34957.4]
  wire [31:0] x341_rd_0_number; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 591:29:@34850.4 sm_x359_inr_Foreach_SAMPLER_BOX.scala 595:339:@34871.4]
  wire [32:0] _GEN_11; // @[Math.scala 461:32:@34969.4]
  wire [31:0] x343_rd_0_number; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 604:29:@34901.4 sm_x359_inr_Foreach_SAMPLER_BOX.scala 608:339:@34922.4]
  wire [33:0] _GEN_12; // @[Math.scala 461:32:@34981.4]
  wire  _T_2016; // @[package.scala 96:25:@35108.4 package.scala 96:25:@35109.4]
  wire  _T_2018; // @[implicits.scala 55:10:@35110.4]
  wire  x563_b237_D73; // @[package.scala 96:25:@35090.4 package.scala 96:25:@35091.4]
  wire  _T_2019; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 659:117:@35111.4]
  wire  x564_b238_D73; // @[package.scala 96:25:@35099.4 package.scala 96:25:@35100.4]
  wire  _T_2020; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 659:123:@35112.4]
  wire [31:0] x251_sum_number; // @[Math.scala 154:22:@32927.4 Math.scala 155:14:@32928.4]
  wire [31:0] x504_x435_D13_number; // @[package.scala 96:25:@32945.4 package.scala 96:25:@32946.4]
  wire [31:0] x506_x413_D21_number; // @[package.scala 96:25:@32963.4 package.scala 96:25:@32964.4]
  wire [31:0] x512_x435_D37_number; // @[package.scala 96:25:@33076.4 package.scala 96:25:@33077.4]
  wire [31:0] x514_x413_D45_number; // @[package.scala 96:25:@33094.4 package.scala 96:25:@33095.4]
  wire [31:0] x515_x251_sum_D24_number; // @[package.scala 96:25:@33103.4 package.scala 96:25:@33104.4]
  wire [31:0] x266_sum_number; // @[Math.scala 154:22:@33495.4 Math.scala 155:14:@33496.4]
  wire [31:0] x519_x460_D13_number; // @[package.scala 96:25:@33504.4 package.scala 96:25:@33505.4]
  wire [31:0] x275_sum_number; // @[Math.scala 154:22:@33889.4 Math.scala 155:14:@33890.4]
  wire [31:0] x522_x482_D13_number; // @[package.scala 96:25:@33898.4 package.scala 96:25:@33899.4]
  wire [31:0] x527_x484_D20_number; // @[package.scala 96:25:@34084.4 package.scala 96:25:@34085.4]
  wire [31:0] x528_x286_sum_D1_number; // @[package.scala 96:25:@34093.4 package.scala 96:25:@34094.4]
  wire [31:0] x291_sum_number; // @[Math.scala 154:22:@34153.4 Math.scala 155:14:@34154.4]
  wire [31:0] x296_sum_number; // @[Math.scala 154:22:@34202.4 Math.scala 155:14:@34203.4]
  wire [31:0] x534_x307_sum_D1_number; // @[package.scala 96:25:@34370.4 package.scala 96:25:@34371.4]
  wire [31:0] x535_x489_D20_number; // @[package.scala 96:25:@34379.4 package.scala 96:25:@34380.4]
  wire [31:0] x312_sum_number; // @[Math.scala 154:22:@34437.4 Math.scala 155:14:@34438.4]
  wire [31:0] x317_sum_number; // @[Math.scala 154:22:@34486.4 Math.scala 155:14:@34487.4]
  wire [31:0] x542_x435_D50_number; // @[package.scala 96:25:@34683.4 package.scala 96:25:@34684.4]
  wire [31:0] x544_x413_D58_number; // @[package.scala 96:25:@34701.4 package.scala 96:25:@34702.4]
  wire [31:0] x546_x251_sum_D37_number; // @[package.scala 96:25:@34719.4 package.scala 96:25:@34720.4]
  wire [31:0] x549_x435_D51_number; // @[package.scala 96:25:@34769.4 package.scala 96:25:@34770.4]
  wire [31:0] x551_x413_D59_number; // @[package.scala 96:25:@34787.4 package.scala 96:25:@34788.4]
  wire [31:0] x552_x251_sum_D38_number; // @[package.scala 96:25:@34796.4 package.scala 96:25:@34797.4]
  wire [31:0] x553_x460_D27_number; // @[package.scala 96:25:@34829.4 package.scala 96:25:@34830.4]
  wire [31:0] x554_x266_sum_D14_number; // @[package.scala 96:25:@34838.4 package.scala 96:25:@34839.4]
  wire [31:0] x556_x484_D34_number; // @[package.scala 96:25:@34880.4 package.scala 96:25:@34881.4]
  wire [31:0] x557_x286_sum_D15_number; // @[package.scala 96:25:@34889.4 package.scala 96:25:@34890.4]
  wire [31:0] x559_x291_sum_D14_number; // @[package.scala 96:25:@34931.4 package.scala 96:25:@34932.4]
  wire [32:0] _T_1961; // @[package.scala 96:25:@34975.4 package.scala 96:25:@34976.4]
  wire [33:0] _T_1966; // @[package.scala 96:25:@34987.4 package.scala 96:25:@34988.4]
  _ _ ( // @[Math.scala 720:24:@32384.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@32396.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@32419.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x241_lb_0 x241_lb_0 ( // @[m_x241_lb_0.scala 35:17:@32429.4]
    .clock(x241_lb_0_clock),
    .reset(x241_lb_0_reset),
    .io_rPort_8_banks_1(x241_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x241_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x241_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x241_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x241_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x241_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x241_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x241_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x241_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x241_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x241_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x241_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x241_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x241_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x241_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x241_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x241_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x241_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x241_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x241_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x241_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x241_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x241_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x241_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x241_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x241_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x241_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x241_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x241_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x241_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x241_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x241_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x241_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x241_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x241_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x241_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x241_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x241_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x241_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x241_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x241_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x241_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x241_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x241_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x241_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x241_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x241_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x241_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x241_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x241_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x241_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x241_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x241_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x241_lb_0_io_rPort_0_output_0),
    .io_wPort_0_banks_1(x241_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x241_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x241_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x241_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x241_lb_0_io_wPort_0_en_0)
  );
  x242_lb2_0 x242_lb2_0 ( // @[m_x242_lb2_0.scala 30:17:@32496.4]
    .clock(x242_lb2_0_clock),
    .reset(x242_lb2_0_reset),
    .io_rPort_3_banks_1(x242_lb2_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x242_lb2_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x242_lb2_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x242_lb2_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x242_lb2_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x242_lb2_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x242_lb2_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x242_lb2_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x242_lb2_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x242_lb2_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x242_lb2_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x242_lb2_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x242_lb2_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x242_lb2_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x242_lb2_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x242_lb2_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x242_lb2_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x242_lb2_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x242_lb2_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x242_lb2_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x242_lb2_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x242_lb2_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x242_lb2_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x242_lb2_0_io_rPort_0_output_0),
    .io_wPort_0_banks_1(x242_lb2_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x242_lb2_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x242_lb2_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x242_lb2_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x242_lb2_0_io_wPort_0_en_0)
  );
  x223_sum x416_sum_1 ( // @[Math.scala 150:24:@32591.4]
    .clock(x416_sum_1_clock),
    .reset(x416_sum_1_reset),
    .io_a(x416_sum_1_io_a),
    .io_b(x416_sum_1_io_b),
    .io_flow(x416_sum_1_io_flow),
    .io_result(x416_sum_1_io_result)
  );
  x223_sum x419_sum_1 ( // @[Math.scala 150:24:@32629.4]
    .clock(x419_sum_1_clock),
    .reset(x419_sum_1_reset),
    .io_a(x419_sum_1_io_a),
    .io_b(x419_sum_1_io_b),
    .io_flow(x419_sum_1_io_flow),
    .io_result(x419_sum_1_io_result)
  );
  x223_sum x422_sum_1 ( // @[Math.scala 150:24:@32667.4]
    .clock(x422_sum_1_clock),
    .reset(x422_sum_1_reset),
    .io_a(x422_sum_1_io_a),
    .io_b(x422_sum_1_io_b),
    .io_flow(x422_sum_1_io_flow),
    .io_result(x422_sum_1_io_result)
  );
  x223_sum x425_sum_1 ( // @[Math.scala 150:24:@32705.4]
    .clock(x425_sum_1_clock),
    .reset(x425_sum_1_reset),
    .io_a(x425_sum_1_io_a),
    .io_b(x425_sum_1_io_b),
    .io_flow(x425_sum_1_io_flow),
    .io_result(x425_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_1 ( // @[package.scala 93:22:@32728.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_2 ( // @[package.scala 93:22:@32746.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x223_sum x428_sum_1 ( // @[Math.scala 150:24:@32759.4]
    .clock(x428_sum_1_clock),
    .reset(x428_sum_1_reset),
    .io_a(x428_sum_1_io_a),
    .io_b(x428_sum_1_io_b),
    .io_flow(x428_sum_1_io_flow),
    .io_result(x428_sum_1_io_result)
  );
  x223_sum x431_sum_1 ( // @[Math.scala 150:24:@32797.4]
    .clock(x431_sum_1_clock),
    .reset(x431_sum_1_reset),
    .io_a(x431_sum_1_io_a),
    .io_b(x431_sum_1_io_b),
    .io_flow(x431_sum_1_io_flow),
    .io_result(x431_sum_1_io_result)
  );
  x410_sub x434_sub_1 ( // @[Math.scala 191:24:@32823.4]
    .clock(x434_sub_1_clock),
    .reset(x434_sub_1_reset),
    .io_a(x434_sub_1_io_a),
    .io_b(x434_sub_1_io_b),
    .io_flow(x434_sub_1_io_flow),
    .io_result(x434_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@32833.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@32842.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_5 ( // @[package.scala 93:22:@32851.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  x223_sum x438_sum_1 ( // @[Math.scala 150:24:@32890.4]
    .clock(x438_sum_1_clock),
    .reset(x438_sum_1_reset),
    .io_a(x438_sum_1_io_a),
    .io_b(x438_sum_1_io_b),
    .io_flow(x438_sum_1_io_flow),
    .io_result(x438_sum_1_io_result)
  );
  x250_div x250_div_1 ( // @[Math.scala 327:24:@32902.4]
    .clock(x250_div_1_clock),
    .io_a(x250_div_1_io_a),
    .io_flow(x250_div_1_io_flow),
    .io_result(x250_div_1_io_result)
  );
  RetimeWrapper_243 RetimeWrapper_6 ( // @[package.scala 93:22:@32912.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x223_sum x251_sum_1 ( // @[Math.scala 150:24:@32921.4]
    .clock(x251_sum_1_clock),
    .reset(x251_sum_1_reset),
    .io_a(x251_sum_1_io_a),
    .io_b(x251_sum_1_io_b),
    .io_flow(x251_sum_1_io_flow),
    .io_result(x251_sum_1_io_result)
  );
  RetimeWrapper_245 RetimeWrapper_7 ( // @[package.scala 93:22:@32931.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_8 ( // @[package.scala 93:22:@32940.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_245 RetimeWrapper_9 ( // @[package.scala 93:22:@32949.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_10 ( // @[package.scala 93:22:@32958.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_249 RetimeWrapper_11 ( // @[package.scala 93:22:@32967.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_245 RetimeWrapper_12 ( // @[package.scala 93:22:@32978.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_251 RetimeWrapper_13 ( // @[package.scala 93:22:@32999.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@33015.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_251 RetimeWrapper_15 ( // @[package.scala 93:22:@33024.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 ( // @[package.scala 93:22:@33038.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_245 RetimeWrapper_17 ( // @[package.scala 93:22:@33053.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_256 RetimeWrapper_18 ( // @[package.scala 93:22:@33062.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_257 RetimeWrapper_19 ( // @[package.scala 93:22:@33071.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_256 RetimeWrapper_20 ( // @[package.scala 93:22:@33080.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_259 RetimeWrapper_21 ( // @[package.scala 93:22:@33089.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_260 RetimeWrapper_22 ( // @[package.scala 93:22:@33098.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_256 RetimeWrapper_23 ( // @[package.scala 93:22:@33110.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  x410_sub x260_rdcol_1 ( // @[Math.scala 191:24:@33133.4]
    .clock(x260_rdcol_1_clock),
    .reset(x260_rdcol_1_reset),
    .io_a(x260_rdcol_1_io_a),
    .io_b(x260_rdcol_1_io_b),
    .io_flow(x260_rdcol_1_io_flow),
    .io_result(x260_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_24 ( // @[package.scala 93:22:@33148.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@33157.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  x223_sum x441_sum_1 ( // @[Math.scala 150:24:@33200.4]
    .clock(x441_sum_1_clock),
    .reset(x441_sum_1_reset),
    .io_a(x441_sum_1_io_a),
    .io_b(x441_sum_1_io_b),
    .io_flow(x441_sum_1_io_flow),
    .io_result(x441_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_26 ( // @[package.scala 93:22:@33223.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_27 ( // @[package.scala 93:22:@33241.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x223_sum x444_sum_1 ( // @[Math.scala 150:24:@33254.4]
    .clock(x444_sum_1_clock),
    .reset(x444_sum_1_reset),
    .io_a(x444_sum_1_io_a),
    .io_b(x444_sum_1_io_b),
    .io_flow(x444_sum_1_io_flow),
    .io_result(x444_sum_1_io_result)
  );
  x223_sum x447_sum_1 ( // @[Math.scala 150:24:@33292.4]
    .clock(x447_sum_1_clock),
    .reset(x447_sum_1_reset),
    .io_a(x447_sum_1_io_a),
    .io_b(x447_sum_1_io_b),
    .io_flow(x447_sum_1_io_flow),
    .io_result(x447_sum_1_io_result)
  );
  x223_sum x450_sum_1 ( // @[Math.scala 150:24:@33330.4]
    .clock(x450_sum_1_clock),
    .reset(x450_sum_1_reset),
    .io_a(x450_sum_1_io_a),
    .io_b(x450_sum_1_io_b),
    .io_flow(x450_sum_1_io_flow),
    .io_result(x450_sum_1_io_result)
  );
  x223_sum x453_sum_1 ( // @[Math.scala 150:24:@33368.4]
    .clock(x453_sum_1_clock),
    .reset(x453_sum_1_reset),
    .io_a(x453_sum_1_io_a),
    .io_b(x453_sum_1_io_b),
    .io_flow(x453_sum_1_io_flow),
    .io_result(x453_sum_1_io_result)
  );
  x223_sum x456_sum_1 ( // @[Math.scala 150:24:@33406.4]
    .clock(x456_sum_1_clock),
    .reset(x456_sum_1_reset),
    .io_a(x456_sum_1_io_a),
    .io_b(x456_sum_1_io_b),
    .io_flow(x456_sum_1_io_flow),
    .io_result(x456_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_28 ( // @[package.scala 93:22:@33421.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper RetimeWrapper_29 ( // @[package.scala 93:22:@33435.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  x410_sub x459_sub_1 ( // @[Math.scala 191:24:@33446.4]
    .clock(x459_sub_1_clock),
    .reset(x459_sub_1_reset),
    .io_a(x459_sub_1_io_a),
    .io_b(x459_sub_1_io_b),
    .io_flow(x459_sub_1_io_flow),
    .io_result(x459_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_30 ( // @[package.scala 93:22:@33456.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  x250_div x265_div_1 ( // @[Math.scala 327:24:@33470.4]
    .clock(x265_div_1_clock),
    .io_a(x265_div_1_io_a),
    .io_flow(x265_div_1_io_flow),
    .io_result(x265_div_1_io_result)
  );
  RetimeWrapper_277 RetimeWrapper_31 ( // @[package.scala 93:22:@33480.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  x223_sum x266_sum_1 ( // @[Math.scala 150:24:@33489.4]
    .clock(x266_sum_1_clock),
    .reset(x266_sum_1_reset),
    .io_a(x266_sum_1_io_a),
    .io_b(x266_sum_1_io_b),
    .io_flow(x266_sum_1_io_flow),
    .io_result(x266_sum_1_io_result)
  );
  RetimeWrapper_246 RetimeWrapper_32 ( // @[package.scala 93:22:@33499.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_280 RetimeWrapper_33 ( // @[package.scala 93:22:@33508.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_256 RetimeWrapper_34 ( // @[package.scala 93:22:@33520.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  x410_sub x269_rdcol_1 ( // @[Math.scala 191:24:@33543.4]
    .clock(x269_rdcol_1_clock),
    .reset(x269_rdcol_1_reset),
    .io_a(x269_rdcol_1_io_a),
    .io_b(x269_rdcol_1_io_b),
    .io_flow(x269_rdcol_1_io_flow),
    .io_result(x269_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_35 ( // @[package.scala 93:22:@33560.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  x223_sum x463_sum_1 ( // @[Math.scala 150:24:@33603.4]
    .clock(x463_sum_1_clock),
    .reset(x463_sum_1_reset),
    .io_a(x463_sum_1_io_a),
    .io_b(x463_sum_1_io_b),
    .io_flow(x463_sum_1_io_flow),
    .io_result(x463_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_36 ( // @[package.scala 93:22:@33626.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_37 ( // @[package.scala 93:22:@33644.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  x223_sum x466_sum_1 ( // @[Math.scala 150:24:@33657.4]
    .clock(x466_sum_1_clock),
    .reset(x466_sum_1_reset),
    .io_a(x466_sum_1_io_a),
    .io_b(x466_sum_1_io_b),
    .io_flow(x466_sum_1_io_flow),
    .io_result(x466_sum_1_io_result)
  );
  x223_sum x469_sum_1 ( // @[Math.scala 150:24:@33695.4]
    .clock(x469_sum_1_clock),
    .reset(x469_sum_1_reset),
    .io_a(x469_sum_1_io_a),
    .io_b(x469_sum_1_io_b),
    .io_flow(x469_sum_1_io_flow),
    .io_result(x469_sum_1_io_result)
  );
  x223_sum x472_sum_1 ( // @[Math.scala 150:24:@33733.4]
    .clock(x472_sum_1_clock),
    .reset(x472_sum_1_reset),
    .io_a(x472_sum_1_io_a),
    .io_b(x472_sum_1_io_b),
    .io_flow(x472_sum_1_io_flow),
    .io_result(x472_sum_1_io_result)
  );
  x223_sum x475_sum_1 ( // @[Math.scala 150:24:@33771.4]
    .clock(x475_sum_1_clock),
    .reset(x475_sum_1_reset),
    .io_a(x475_sum_1_io_a),
    .io_b(x475_sum_1_io_b),
    .io_flow(x475_sum_1_io_flow),
    .io_result(x475_sum_1_io_result)
  );
  x223_sum x478_sum_1 ( // @[Math.scala 150:24:@33809.4]
    .clock(x478_sum_1_clock),
    .reset(x478_sum_1_reset),
    .io_a(x478_sum_1_io_a),
    .io_b(x478_sum_1_io_b),
    .io_flow(x478_sum_1_io_flow),
    .io_result(x478_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_38 ( // @[package.scala 93:22:@33824.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper RetimeWrapper_39 ( // @[package.scala 93:22:@33838.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  x410_sub x481_sub_1 ( // @[Math.scala 191:24:@33849.4]
    .clock(x481_sub_1_clock),
    .reset(x481_sub_1_reset),
    .io_a(x481_sub_1_io_a),
    .io_b(x481_sub_1_io_b),
    .io_flow(x481_sub_1_io_flow),
    .io_result(x481_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_40 ( // @[package.scala 93:22:@33859.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  x250_div x274_div_1 ( // @[Math.scala 327:24:@33873.4]
    .clock(x274_div_1_clock),
    .io_a(x274_div_1_io_a),
    .io_flow(x274_div_1_io_flow),
    .io_result(x274_div_1_io_result)
  );
  x223_sum x275_sum_1 ( // @[Math.scala 150:24:@33883.4]
    .clock(x275_sum_1_clock),
    .reset(x275_sum_1_reset),
    .io_a(x275_sum_1_io_a),
    .io_b(x275_sum_1_io_b),
    .io_flow(x275_sum_1_io_flow),
    .io_result(x275_sum_1_io_result)
  );
  RetimeWrapper_246 RetimeWrapper_41 ( // @[package.scala 93:22:@33893.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_280 RetimeWrapper_42 ( // @[package.scala 93:22:@33902.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_256 RetimeWrapper_43 ( // @[package.scala 93:22:@33914.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  x410_sub x278_rdrow_1 ( // @[Math.scala 191:24:@33937.4]
    .clock(x278_rdrow_1_clock),
    .reset(x278_rdrow_1_reset),
    .io_a(x278_rdrow_1_io_a),
    .io_b(x278_rdrow_1_io_b),
    .io_flow(x278_rdrow_1_io_flow),
    .io_result(x278_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_44 ( // @[package.scala 93:22:@33963.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper RetimeWrapper_45 ( // @[package.scala 93:22:@33972.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_46 ( // @[package.scala 93:22:@33994.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_47 ( // @[package.scala 93:22:@34020.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  x223_sum x487_sum_1 ( // @[Math.scala 150:24:@34041.4]
    .clock(x487_sum_1_clock),
    .reset(x487_sum_1_reset),
    .io_a(x487_sum_1_io_a),
    .io_b(x487_sum_1_io_b),
    .io_flow(x487_sum_1_io_flow),
    .io_result(x487_sum_1_io_result)
  );
  RetimeWrapper_251 RetimeWrapper_48 ( // @[package.scala 93:22:@34051.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_307 RetimeWrapper_49 ( // @[package.scala 93:22:@34060.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  x223_sum x286_sum_1 ( // @[Math.scala 150:24:@34069.4]
    .clock(x286_sum_1_clock),
    .reset(x286_sum_1_reset),
    .io_a(x286_sum_1_io_a),
    .io_b(x286_sum_1_io_b),
    .io_flow(x286_sum_1_io_flow),
    .io_result(x286_sum_1_io_result)
  );
  RetimeWrapper_249 RetimeWrapper_50 ( // @[package.scala 93:22:@34079.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_51 ( // @[package.scala 93:22:@34088.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_280 RetimeWrapper_52 ( // @[package.scala 93:22:@34097.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_256 RetimeWrapper_53 ( // @[package.scala 93:22:@34109.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_313 RetimeWrapper_54 ( // @[package.scala 93:22:@34136.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  x223_sum x291_sum_1 ( // @[Math.scala 150:24:@34147.4]
    .clock(x291_sum_1_clock),
    .reset(x291_sum_1_reset),
    .io_a(x291_sum_1_io_a),
    .io_b(x291_sum_1_io_b),
    .io_flow(x291_sum_1_io_flow),
    .io_result(x291_sum_1_io_result)
  );
  RetimeWrapper_280 RetimeWrapper_55 ( // @[package.scala 93:22:@34157.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_256 RetimeWrapper_56 ( // @[package.scala 93:22:@34169.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  x223_sum x296_sum_1 ( // @[Math.scala 150:24:@34196.4]
    .clock(x296_sum_1_clock),
    .reset(x296_sum_1_reset),
    .io_a(x296_sum_1_io_a),
    .io_b(x296_sum_1_io_b),
    .io_flow(x296_sum_1_io_flow),
    .io_result(x296_sum_1_io_result)
  );
  RetimeWrapper_280 RetimeWrapper_57 ( // @[package.scala 93:22:@34206.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_256 RetimeWrapper_58 ( // @[package.scala 93:22:@34218.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  x410_sub x299_rdrow_1 ( // @[Math.scala 191:24:@34241.4]
    .clock(x299_rdrow_1_clock),
    .reset(x299_rdrow_1_reset),
    .io_a(x299_rdrow_1_io_a),
    .io_b(x299_rdrow_1_io_b),
    .io_flow(x299_rdrow_1_io_flow),
    .io_result(x299_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_59 ( // @[package.scala 93:22:@34267.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_60 ( // @[package.scala 93:22:@34289.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_61 ( // @[package.scala 93:22:@34315.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x223_sum x492_sum_1 ( // @[Math.scala 150:24:@34336.4]
    .clock(x492_sum_1_clock),
    .reset(x492_sum_1_reset),
    .io_a(x492_sum_1_io_a),
    .io_b(x492_sum_1_io_b),
    .io_flow(x492_sum_1_io_flow),
    .io_result(x492_sum_1_io_result)
  );
  RetimeWrapper_307 RetimeWrapper_62 ( // @[package.scala 93:22:@34346.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  x223_sum x307_sum_1 ( // @[Math.scala 150:24:@34355.4]
    .clock(x307_sum_1_clock),
    .reset(x307_sum_1_reset),
    .io_a(x307_sum_1_io_a),
    .io_b(x307_sum_1_io_b),
    .io_flow(x307_sum_1_io_flow),
    .io_result(x307_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_63 ( // @[package.scala 93:22:@34365.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_249 RetimeWrapper_64 ( // @[package.scala 93:22:@34374.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_280 RetimeWrapper_65 ( // @[package.scala 93:22:@34383.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_256 RetimeWrapper_66 ( // @[package.scala 93:22:@34395.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_313 RetimeWrapper_67 ( // @[package.scala 93:22:@34422.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  x223_sum x312_sum_1 ( // @[Math.scala 150:24:@34431.4]
    .clock(x312_sum_1_clock),
    .reset(x312_sum_1_reset),
    .io_a(x312_sum_1_io_a),
    .io_b(x312_sum_1_io_b),
    .io_flow(x312_sum_1_io_flow),
    .io_result(x312_sum_1_io_result)
  );
  RetimeWrapper_280 RetimeWrapper_68 ( // @[package.scala 93:22:@34441.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_256 RetimeWrapper_69 ( // @[package.scala 93:22:@34453.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  x223_sum x317_sum_1 ( // @[Math.scala 150:24:@34480.4]
    .clock(x317_sum_1_clock),
    .reset(x317_sum_1_reset),
    .io_a(x317_sum_1_io_a),
    .io_b(x317_sum_1_io_b),
    .io_flow(x317_sum_1_io_flow),
    .io_result(x317_sum_1_io_result)
  );
  RetimeWrapper_280 RetimeWrapper_70 ( // @[package.scala 93:22:@34490.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_256 RetimeWrapper_71 ( // @[package.scala 93:22:@34502.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  x325_x7 x325_x7_1 ( // @[Math.scala 150:24:@34550.4]
    .clock(x325_x7_1_clock),
    .reset(x325_x7_1_reset),
    .io_a(x325_x7_1_io_a),
    .io_b(x325_x7_1_io_b),
    .io_flow(x325_x7_1_io_flow),
    .io_result(x325_x7_1_io_result)
  );
  x325_x7 x326_x8_1 ( // @[Math.scala 150:24:@34560.4]
    .clock(x326_x8_1_clock),
    .reset(x326_x8_1_reset),
    .io_a(x326_x8_1_io_a),
    .io_b(x326_x8_1_io_b),
    .io_flow(x326_x8_1_io_flow),
    .io_result(x326_x8_1_io_result)
  );
  x325_x7 x327_x7_1 ( // @[Math.scala 150:24:@34570.4]
    .clock(x327_x7_1_clock),
    .reset(x327_x7_1_reset),
    .io_a(x327_x7_1_io_a),
    .io_b(x327_x7_1_io_b),
    .io_flow(x327_x7_1_io_flow),
    .io_result(x327_x7_1_io_result)
  );
  x325_x7 x328_x8_1 ( // @[Math.scala 150:24:@34580.4]
    .clock(x328_x8_1_clock),
    .reset(x328_x8_1_reset),
    .io_a(x328_x8_1_io_a),
    .io_b(x328_x8_1_io_b),
    .io_flow(x328_x8_1_io_flow),
    .io_result(x328_x8_1_io_result)
  );
  x325_x7 x329_x7_1 ( // @[Math.scala 150:24:@34590.4]
    .clock(x329_x7_1_clock),
    .reset(x329_x7_1_reset),
    .io_a(x329_x7_1_io_a),
    .io_b(x329_x7_1_io_b),
    .io_flow(x329_x7_1_io_flow),
    .io_result(x329_x7_1_io_result)
  );
  x325_x7 x330_x8_1 ( // @[Math.scala 150:24:@34600.4]
    .clock(x330_x8_1_clock),
    .reset(x330_x8_1_reset),
    .io_a(x330_x8_1_io_a),
    .io_b(x330_x8_1_io_b),
    .io_flow(x330_x8_1_io_flow),
    .io_result(x330_x8_1_io_result)
  );
  x325_x7 x331_x7_1 ( // @[Math.scala 150:24:@34610.4]
    .clock(x331_x7_1_clock),
    .reset(x331_x7_1_reset),
    .io_a(x331_x7_1_io_a),
    .io_b(x331_x7_1_io_b),
    .io_flow(x331_x7_1_io_flow),
    .io_result(x331_x7_1_io_result)
  );
  RetimeWrapper_345 RetimeWrapper_72 ( // @[package.scala 93:22:@34620.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  x325_x7 x332_sum_1 ( // @[Math.scala 150:24:@34629.4]
    .clock(x332_sum_1_clock),
    .reset(x332_sum_1_reset),
    .io_a(x332_sum_1_io_a),
    .io_b(x332_sum_1_io_b),
    .io_flow(x332_sum_1_io_flow),
    .io_result(x332_sum_1_io_result)
  );
  x333 x333_1 ( // @[Math.scala 720:24:@34639.4]
    .io_b(x333_1_io_b),
    .io_result(x333_1_io_result)
  );
  x334_mul x334_mul_1 ( // @[Math.scala 262:24:@34650.4]
    .clock(x334_mul_1_clock),
    .io_a(x334_mul_1_io_a),
    .io_b(x334_mul_1_io_b),
    .io_flow(x334_mul_1_io_flow),
    .io_result(x334_mul_1_io_result)
  );
  x335 x335_1 ( // @[Math.scala 720:24:@34660.4]
    .io_b(x335_1_io_b),
    .io_result(x335_1_io_result)
  );
  RetimeWrapper_347 RetimeWrapper_73 ( // @[package.scala 93:22:@34669.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_348 RetimeWrapper_74 ( // @[package.scala 93:22:@34678.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_347 RetimeWrapper_75 ( // @[package.scala 93:22:@34687.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_350 RetimeWrapper_76 ( // @[package.scala 93:22:@34696.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_77 ( // @[package.scala 93:22:@34705.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_257 RetimeWrapper_78 ( // @[package.scala 93:22:@34714.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_347 RetimeWrapper_79 ( // @[package.scala 93:22:@34725.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_354 RetimeWrapper_80 ( // @[package.scala 93:22:@34746.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_355 RetimeWrapper_81 ( // @[package.scala 93:22:@34755.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_356 RetimeWrapper_82 ( // @[package.scala 93:22:@34764.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_355 RetimeWrapper_83 ( // @[package.scala 93:22:@34773.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_358 RetimeWrapper_84 ( // @[package.scala 93:22:@34782.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_359 RetimeWrapper_85 ( // @[package.scala 93:22:@34791.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_355 RetimeWrapper_86 ( // @[package.scala 93:22:@34803.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_361 RetimeWrapper_87 ( // @[package.scala 93:22:@34824.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_362 RetimeWrapper_88 ( // @[package.scala 93:22:@34833.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_363 RetimeWrapper_89 ( // @[package.scala 93:22:@34842.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_355 RetimeWrapper_90 ( // @[package.scala 93:22:@34854.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_365 RetimeWrapper_91 ( // @[package.scala 93:22:@34875.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_366 RetimeWrapper_92 ( // @[package.scala 93:22:@34884.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_363 RetimeWrapper_93 ( // @[package.scala 93:22:@34893.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_355 RetimeWrapper_94 ( // @[package.scala 93:22:@34905.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_362 RetimeWrapper_95 ( // @[package.scala 93:22:@34926.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_363 RetimeWrapper_96 ( // @[package.scala 93:22:@34935.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_355 RetimeWrapper_97 ( // @[package.scala 93:22:@34947.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_372 RetimeWrapper_98 ( // @[package.scala 93:22:@34970.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_373 RetimeWrapper_99 ( // @[package.scala 93:22:@34982.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_100 ( // @[package.scala 93:22:@34992.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  x325_x7 x349_x9_1 ( // @[Math.scala 150:24:@35001.4]
    .clock(x349_x9_1_clock),
    .reset(x349_x9_1_reset),
    .io_a(x349_x9_1_io_a),
    .io_b(x349_x9_1_io_b),
    .io_flow(x349_x9_1_io_flow),
    .io_result(x349_x9_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_101 ( // @[package.scala 93:22:@35011.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  x325_x7 x350_x10_1 ( // @[Math.scala 150:24:@35022.4]
    .clock(x350_x10_1_clock),
    .reset(x350_x10_1_reset),
    .io_a(x350_x10_1_io_a),
    .io_b(x350_x10_1_io_b),
    .io_flow(x350_x10_1_io_flow),
    .io_result(x350_x10_1_io_result)
  );
  x325_x7 x351_sum_1 ( // @[Math.scala 150:24:@35032.4]
    .clock(x351_sum_1_clock),
    .reset(x351_sum_1_reset),
    .io_a(x351_sum_1_io_a),
    .io_b(x351_sum_1_io_b),
    .io_flow(x351_sum_1_io_flow),
    .io_result(x351_sum_1_io_result)
  );
  x333 x352_1 ( // @[Math.scala 720:24:@35042.4]
    .io_b(x352_1_io_b),
    .io_result(x352_1_io_result)
  );
  x334_mul x353_mul_1 ( // @[Math.scala 262:24:@35053.4]
    .clock(x353_mul_1_clock),
    .io_a(x353_mul_1_io_a),
    .io_b(x353_mul_1_io_b),
    .io_flow(x353_mul_1_io_flow),
    .io_result(x353_mul_1_io_result)
  );
  x335 x354_1 ( // @[Math.scala 720:24:@35063.4]
    .io_b(x354_1_io_b),
    .io_result(x354_1_io_result)
  );
  RetimeWrapper_345 RetimeWrapper_102 ( // @[package.scala 93:22:@35076.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_380 RetimeWrapper_103 ( // @[package.scala 93:22:@35085.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_380 RetimeWrapper_104 ( // @[package.scala 93:22:@35094.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_380 RetimeWrapper_105 ( // @[package.scala 93:22:@35103.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  assign b237 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 62:18:@32404.4]
  assign b238 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 63:18:@32405.4]
  assign _T_205 = b237 & b238; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 67:30:@32407.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 67:37:@32408.4]
  assign _T_210 = io_in_x209_TID == 8'h0; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 69:76:@32413.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 69:62:@32414.4]
  assign _T_213 = io_in_x209_TDEST == 8'h0; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 69:101:@32415.4]
  assign b235_number = __io_result; // @[Math.scala 723:22:@32389.4 Math.scala 724:14:@32390.4]
  assign _T_242 = $signed(b235_number); // @[Math.scala 406:49:@32542.4]
  assign _T_244 = $signed(_T_242) & $signed(32'sh3); // @[Math.scala 406:56:@32544.4]
  assign _T_245 = $signed(_T_244); // @[Math.scala 406:56:@32545.4]
  assign x412_number = $unsigned(_T_245); // @[implicits.scala 133:21:@32546.4]
  assign _T_255 = $signed(x412_number); // @[Math.scala 406:49:@32555.4]
  assign _T_257 = $signed(_T_255) & $signed(32'sh3); // @[Math.scala 406:56:@32557.4]
  assign _T_258 = $signed(_T_257); // @[Math.scala 406:56:@32558.4]
  assign b236_number = __1_io_result; // @[Math.scala 723:22:@32401.4 Math.scala 724:14:@32402.4]
  assign _T_262 = b236_number[31]; // @[FixedPoint.scala 50:25:@32564.4]
  assign _T_266 = _T_262 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@32566.4]
  assign _T_267 = b236_number[31:16]; // @[FixedPoint.scala 18:52:@32567.4]
  assign _T_273 = _T_267 == 16'hffff; // @[Math.scala 451:55:@32569.4]
  assign _T_274 = b236_number[15:0]; // @[FixedPoint.scala 18:52:@32570.4]
  assign _T_280 = _T_274 != 16'h0; // @[Math.scala 451:110:@32572.4]
  assign _T_281 = _T_273 & _T_280; // @[Math.scala 451:94:@32573.4]
  assign _T_283 = {_T_266,_T_267}; // @[Cat.scala 30:58:@32575.4]
  assign _T_293 = $signed(b236_number); // @[Math.scala 406:49:@32583.4]
  assign _T_295 = $signed(_T_293) & $signed(32'shffff); // @[Math.scala 406:56:@32585.4]
  assign _T_296 = $signed(_T_295); // @[Math.scala 406:56:@32586.4]
  assign x416_sum_number = x416_sum_1_io_result; // @[Math.scala 154:22:@32597.4 Math.scala 155:14:@32598.4]
  assign _T_303 = x416_sum_number[31]; // @[FixedPoint.scala 50:25:@32602.4]
  assign _T_307 = _T_303 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@32604.4]
  assign _T_308 = x416_sum_number[31:8]; // @[FixedPoint.scala 18:52:@32605.4]
  assign _T_314 = _T_308 == 24'hffffff; // @[Math.scala 451:55:@32607.4]
  assign _T_315 = x416_sum_number[7:0]; // @[FixedPoint.scala 18:52:@32608.4]
  assign _T_321 = _T_315 != 8'h0; // @[Math.scala 451:110:@32610.4]
  assign _T_322 = _T_314 & _T_321; // @[Math.scala 451:94:@32611.4]
  assign _T_324 = {_T_307,_T_308}; // @[Cat.scala 30:58:@32613.4]
  assign _T_334 = $signed(x416_sum_number); // @[Math.scala 406:49:@32621.4]
  assign _T_336 = $signed(_T_334) & $signed(32'shff); // @[Math.scala 406:56:@32623.4]
  assign _T_337 = $signed(_T_336); // @[Math.scala 406:56:@32624.4]
  assign x419_sum_number = x419_sum_1_io_result; // @[Math.scala 154:22:@32635.4 Math.scala 155:14:@32636.4]
  assign _T_344 = x419_sum_number[31]; // @[FixedPoint.scala 50:25:@32640.4]
  assign _T_348 = _T_344 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@32642.4]
  assign _T_349 = x419_sum_number[31:4]; // @[FixedPoint.scala 18:52:@32643.4]
  assign _T_355 = _T_349 == 28'hfffffff; // @[Math.scala 451:55:@32645.4]
  assign _T_356 = x419_sum_number[3:0]; // @[FixedPoint.scala 18:52:@32646.4]
  assign _T_362 = _T_356 != 4'h0; // @[Math.scala 451:110:@32648.4]
  assign _T_363 = _T_355 & _T_362; // @[Math.scala 451:94:@32649.4]
  assign _T_365 = {_T_348,_T_349}; // @[Cat.scala 30:58:@32651.4]
  assign _T_375 = $signed(x419_sum_number); // @[Math.scala 406:49:@32659.4]
  assign _T_377 = $signed(_T_375) & $signed(32'shf); // @[Math.scala 406:56:@32661.4]
  assign _T_378 = $signed(_T_377); // @[Math.scala 406:56:@32662.4]
  assign x422_sum_number = x422_sum_1_io_result; // @[Math.scala 154:22:@32673.4 Math.scala 155:14:@32674.4]
  assign _T_385 = x422_sum_number[31]; // @[FixedPoint.scala 50:25:@32678.4]
  assign _T_389 = _T_385 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@32680.4]
  assign _T_390 = x422_sum_number[31:2]; // @[FixedPoint.scala 18:52:@32681.4]
  assign _T_396 = _T_390 == 30'h3fffffff; // @[Math.scala 451:55:@32683.4]
  assign _T_397 = x422_sum_number[1:0]; // @[FixedPoint.scala 18:52:@32684.4]
  assign _T_403 = _T_397 != 2'h0; // @[Math.scala 451:110:@32686.4]
  assign _T_404 = _T_396 & _T_403; // @[Math.scala 451:94:@32687.4]
  assign _T_406 = {_T_389,_T_390}; // @[Cat.scala 30:58:@32689.4]
  assign _T_416 = $signed(x422_sum_number); // @[Math.scala 406:49:@32697.4]
  assign _T_418 = $signed(_T_416) & $signed(32'sh3); // @[Math.scala 406:56:@32699.4]
  assign _T_419 = $signed(_T_418); // @[Math.scala 406:56:@32700.4]
  assign x425_sum_number = x425_sum_1_io_result; // @[Math.scala 154:22:@32711.4 Math.scala 155:14:@32712.4]
  assign _T_426 = x425_sum_number[31]; // @[FixedPoint.scala 50:25:@32716.4]
  assign _T_430 = _T_426 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@32718.4]
  assign _T_431 = x425_sum_number[31:2]; // @[FixedPoint.scala 18:52:@32719.4]
  assign _T_437 = _T_431 == 30'h3fffffff; // @[Math.scala 451:55:@32721.4]
  assign _T_438 = x425_sum_number[1:0]; // @[FixedPoint.scala 18:52:@32722.4]
  assign _T_444 = _T_438 != 2'h0; // @[Math.scala 451:110:@32724.4]
  assign _T_445 = _T_437 & _T_444; // @[Math.scala 451:94:@32725.4]
  assign _T_449 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@32733.4 package.scala 96:25:@32734.4]
  assign _T_459 = $signed(x425_sum_number); // @[Math.scala 406:49:@32742.4]
  assign _T_461 = $signed(_T_459) & $signed(32'sh3); // @[Math.scala 406:56:@32744.4]
  assign _T_462 = $signed(_T_461); // @[Math.scala 406:56:@32745.4]
  assign _T_466 = $signed(RetimeWrapper_2_io_out); // @[package.scala 96:25:@32753.4]
  assign x428_sum_number = x428_sum_1_io_result; // @[Math.scala 154:22:@32765.4 Math.scala 155:14:@32766.4]
  assign _T_473 = x428_sum_number[31]; // @[FixedPoint.scala 50:25:@32770.4]
  assign _T_477 = _T_473 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@32772.4]
  assign _T_478 = x428_sum_number[31:2]; // @[FixedPoint.scala 18:52:@32773.4]
  assign _T_484 = _T_478 == 30'h3fffffff; // @[Math.scala 451:55:@32775.4]
  assign _T_485 = x428_sum_number[1:0]; // @[FixedPoint.scala 18:52:@32776.4]
  assign _T_491 = _T_485 != 2'h0; // @[Math.scala 451:110:@32778.4]
  assign _T_492 = _T_484 & _T_491; // @[Math.scala 451:94:@32779.4]
  assign _T_494 = {_T_477,_T_478}; // @[Cat.scala 30:58:@32781.4]
  assign _T_504 = $signed(x428_sum_number); // @[Math.scala 406:49:@32789.4]
  assign _T_506 = $signed(_T_504) & $signed(32'sh3); // @[Math.scala 406:56:@32791.4]
  assign _T_507 = $signed(_T_506); // @[Math.scala 406:56:@32792.4]
  assign x431_sum_number = x431_sum_1_io_result; // @[Math.scala 154:22:@32803.4 Math.scala 155:14:@32804.4]
  assign _T_517 = $signed(x431_sum_number); // @[Math.scala 476:37:@32809.4]
  assign x499_x432_D1 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@32838.4 package.scala 96:25:@32839.4]
  assign x501_x431_sum_D1_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@32856.4 package.scala 96:25:@32857.4]
  assign x434_sub_number = x434_sub_1_io_result; // @[Math.scala 195:22:@32829.4 Math.scala 196:14:@32830.4]
  assign _T_548 = x412_number[31]; // @[FixedPoint.scala 50:25:@32864.4]
  assign _T_552 = _T_548 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@32866.4]
  assign _T_553 = x412_number[31:2]; // @[FixedPoint.scala 18:52:@32867.4]
  assign _T_559 = _T_553 == 30'h3fffffff; // @[Math.scala 451:55:@32869.4]
  assign _T_560 = x412_number[1:0]; // @[FixedPoint.scala 18:52:@32870.4]
  assign _T_566 = _T_560 != 2'h0; // @[Math.scala 451:110:@32872.4]
  assign _T_567 = _T_559 & _T_566; // @[Math.scala 451:94:@32873.4]
  assign _T_569 = {_T_552,_T_553}; // @[Cat.scala 30:58:@32875.4]
  assign x248_1_number = _T_567 ? 32'h0 : _T_569; // @[Math.scala 454:20:@32876.4]
  assign _GEN_0 = {{9'd0}, x248_1_number}; // @[Math.scala 461:32:@32881.4]
  assign _T_574 = _GEN_0 << 9; // @[Math.scala 461:32:@32881.4]
  assign _GEN_1 = {{7'd0}, x248_1_number}; // @[Math.scala 461:32:@32886.4]
  assign _T_577 = _GEN_1 << 7; // @[Math.scala 461:32:@32886.4]
  assign _T_610 = ~ io_sigsIn_break; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 164:101:@32975.4]
  assign _T_614 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@32983.4 package.scala 96:25:@32984.4]
  assign _T_616 = io_rr ? _T_614 : 1'h0; // @[implicits.scala 55:10:@32985.4]
  assign _T_617 = _T_610 & _T_616; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 164:118:@32986.4]
  assign _T_619 = _T_617 & _T_610; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 164:207:@32988.4]
  assign _T_620 = _T_619 & io_sigsIn_backpressure; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 164:226:@32989.4]
  assign x505_b237_D21 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@32954.4 package.scala 96:25:@32955.4]
  assign _T_621 = _T_620 & x505_b237_D21; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 164:252:@32990.4]
  assign x503_b238_D21 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@32936.4 package.scala 96:25:@32937.4]
  assign x508_b235_D23_number = RetimeWrapper_13_io_out; // @[package.scala 96:25:@33004.4 package.scala 96:25:@33005.4]
  assign _T_633 = $signed(x508_b235_D23_number); // @[Math.scala 476:37:@33012.4]
  assign x509_b236_D23_number = RetimeWrapper_15_io_out; // @[package.scala 96:25:@33029.4 package.scala 96:25:@33030.4]
  assign _T_646 = $signed(x509_b236_D23_number); // @[Math.scala 476:37:@33035.4]
  assign x254 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@33020.4 package.scala 96:25:@33021.4]
  assign x255 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@33043.4 package.scala 96:25:@33044.4]
  assign x256 = x254 | x255; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 183:24:@33047.4]
  assign _T_684 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@33115.4 package.scala 96:25:@33116.4]
  assign _T_686 = io_rr ? _T_684 : 1'h0; // @[implicits.scala 55:10:@33117.4]
  assign _T_687 = _T_610 & _T_686; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 202:194:@33118.4]
  assign x510_x257_D21 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@33058.4 package.scala 96:25:@33059.4]
  assign _T_688 = _T_687 & x510_x257_D21; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 202:283:@33119.4]
  assign x513_b237_D45 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@33085.4 package.scala 96:25:@33086.4]
  assign _T_689 = _T_688 & x513_b237_D45; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 202:291:@33120.4]
  assign x511_b238_D45 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@33067.4 package.scala 96:25:@33068.4]
  assign x260_rdcol_number = x260_rdcol_1_io_result; // @[Math.scala 195:22:@33139.4 Math.scala 196:14:@33140.4]
  assign _T_704 = $signed(x260_rdcol_number); // @[Math.scala 476:37:@33145.4]
  assign x516_x254_D1 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@33162.4 package.scala 96:25:@33163.4]
  assign x261 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@33153.4 package.scala 96:25:@33154.4]
  assign x262 = x516_x254_D1 | x261; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 212:24:@33166.4]
  assign _T_718 = x260_rdcol_number[31]; // @[FixedPoint.scala 50:25:@33173.4]
  assign _T_722 = _T_718 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@33175.4]
  assign _T_723 = x260_rdcol_number[31:16]; // @[FixedPoint.scala 18:52:@33176.4]
  assign _T_729 = _T_723 == 16'hffff; // @[Math.scala 451:55:@33178.4]
  assign _T_730 = x260_rdcol_number[15:0]; // @[FixedPoint.scala 18:52:@33179.4]
  assign _T_736 = _T_730 != 16'h0; // @[Math.scala 451:110:@33181.4]
  assign _T_737 = _T_729 & _T_736; // @[Math.scala 451:94:@33182.4]
  assign _T_739 = {_T_722,_T_723}; // @[Cat.scala 30:58:@33184.4]
  assign _T_751 = $signed(_T_704) & $signed(32'shffff); // @[Math.scala 406:56:@33194.4]
  assign _T_752 = $signed(_T_751); // @[Math.scala 406:56:@33195.4]
  assign x441_sum_number = x441_sum_1_io_result; // @[Math.scala 154:22:@33206.4 Math.scala 155:14:@33207.4]
  assign _T_759 = x441_sum_number[31]; // @[FixedPoint.scala 50:25:@33211.4]
  assign _T_763 = _T_759 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@33213.4]
  assign _T_764 = x441_sum_number[31:8]; // @[FixedPoint.scala 18:52:@33214.4]
  assign _T_770 = _T_764 == 24'hffffff; // @[Math.scala 451:55:@33216.4]
  assign _T_771 = x441_sum_number[7:0]; // @[FixedPoint.scala 18:52:@33217.4]
  assign _T_777 = _T_771 != 8'h0; // @[Math.scala 451:110:@33219.4]
  assign _T_778 = _T_770 & _T_777; // @[Math.scala 451:94:@33220.4]
  assign _T_782 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@33228.4 package.scala 96:25:@33229.4]
  assign _T_792 = $signed(x441_sum_number); // @[Math.scala 406:49:@33237.4]
  assign _T_794 = $signed(_T_792) & $signed(32'shff); // @[Math.scala 406:56:@33239.4]
  assign _T_795 = $signed(_T_794); // @[Math.scala 406:56:@33240.4]
  assign _T_799 = $signed(RetimeWrapper_27_io_out); // @[package.scala 96:25:@33248.4]
  assign x444_sum_number = x444_sum_1_io_result; // @[Math.scala 154:22:@33260.4 Math.scala 155:14:@33261.4]
  assign _T_806 = x444_sum_number[31]; // @[FixedPoint.scala 50:25:@33265.4]
  assign _T_810 = _T_806 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@33267.4]
  assign _T_811 = x444_sum_number[31:4]; // @[FixedPoint.scala 18:52:@33268.4]
  assign _T_817 = _T_811 == 28'hfffffff; // @[Math.scala 451:55:@33270.4]
  assign _T_818 = x444_sum_number[3:0]; // @[FixedPoint.scala 18:52:@33271.4]
  assign _T_824 = _T_818 != 4'h0; // @[Math.scala 451:110:@33273.4]
  assign _T_825 = _T_817 & _T_824; // @[Math.scala 451:94:@33274.4]
  assign _T_827 = {_T_810,_T_811}; // @[Cat.scala 30:58:@33276.4]
  assign _T_837 = $signed(x444_sum_number); // @[Math.scala 406:49:@33284.4]
  assign _T_839 = $signed(_T_837) & $signed(32'shf); // @[Math.scala 406:56:@33286.4]
  assign _T_840 = $signed(_T_839); // @[Math.scala 406:56:@33287.4]
  assign x447_sum_number = x447_sum_1_io_result; // @[Math.scala 154:22:@33298.4 Math.scala 155:14:@33299.4]
  assign _T_847 = x447_sum_number[31]; // @[FixedPoint.scala 50:25:@33303.4]
  assign _T_851 = _T_847 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33305.4]
  assign _T_852 = x447_sum_number[31:2]; // @[FixedPoint.scala 18:52:@33306.4]
  assign _T_858 = _T_852 == 30'h3fffffff; // @[Math.scala 451:55:@33308.4]
  assign _T_859 = x447_sum_number[1:0]; // @[FixedPoint.scala 18:52:@33309.4]
  assign _T_865 = _T_859 != 2'h0; // @[Math.scala 451:110:@33311.4]
  assign _T_866 = _T_858 & _T_865; // @[Math.scala 451:94:@33312.4]
  assign _T_868 = {_T_851,_T_852}; // @[Cat.scala 30:58:@33314.4]
  assign _T_878 = $signed(x447_sum_number); // @[Math.scala 406:49:@33322.4]
  assign _T_880 = $signed(_T_878) & $signed(32'sh3); // @[Math.scala 406:56:@33324.4]
  assign _T_881 = $signed(_T_880); // @[Math.scala 406:56:@33325.4]
  assign x450_sum_number = x450_sum_1_io_result; // @[Math.scala 154:22:@33336.4 Math.scala 155:14:@33337.4]
  assign _T_888 = x450_sum_number[31]; // @[FixedPoint.scala 50:25:@33341.4]
  assign _T_892 = _T_888 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33343.4]
  assign _T_893 = x450_sum_number[31:2]; // @[FixedPoint.scala 18:52:@33344.4]
  assign _T_899 = _T_893 == 30'h3fffffff; // @[Math.scala 451:55:@33346.4]
  assign _T_900 = x450_sum_number[1:0]; // @[FixedPoint.scala 18:52:@33347.4]
  assign _T_906 = _T_900 != 2'h0; // @[Math.scala 451:110:@33349.4]
  assign _T_907 = _T_899 & _T_906; // @[Math.scala 451:94:@33350.4]
  assign _T_909 = {_T_892,_T_893}; // @[Cat.scala 30:58:@33352.4]
  assign _T_919 = $signed(x450_sum_number); // @[Math.scala 406:49:@33360.4]
  assign _T_921 = $signed(_T_919) & $signed(32'sh3); // @[Math.scala 406:56:@33362.4]
  assign _T_922 = $signed(_T_921); // @[Math.scala 406:56:@33363.4]
  assign x453_sum_number = x453_sum_1_io_result; // @[Math.scala 154:22:@33374.4 Math.scala 155:14:@33375.4]
  assign _T_929 = x453_sum_number[31]; // @[FixedPoint.scala 50:25:@33379.4]
  assign _T_933 = _T_929 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33381.4]
  assign _T_934 = x453_sum_number[31:2]; // @[FixedPoint.scala 18:52:@33382.4]
  assign _T_940 = _T_934 == 30'h3fffffff; // @[Math.scala 451:55:@33384.4]
  assign _T_941 = x453_sum_number[1:0]; // @[FixedPoint.scala 18:52:@33385.4]
  assign _T_947 = _T_941 != 2'h0; // @[Math.scala 451:110:@33387.4]
  assign _T_948 = _T_940 & _T_947; // @[Math.scala 451:94:@33388.4]
  assign _T_950 = {_T_933,_T_934}; // @[Cat.scala 30:58:@33390.4]
  assign _T_960 = $signed(x453_sum_number); // @[Math.scala 406:49:@33398.4]
  assign _T_962 = $signed(_T_960) & $signed(32'sh3); // @[Math.scala 406:56:@33400.4]
  assign _T_963 = $signed(_T_962); // @[Math.scala 406:56:@33401.4]
  assign x456_sum_number = x456_sum_1_io_result; // @[Math.scala 154:22:@33412.4 Math.scala 155:14:@33413.4]
  assign _T_973 = $signed(x456_sum_number); // @[Math.scala 476:37:@33418.4]
  assign x457 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@33426.4 package.scala 96:25:@33427.4]
  assign x517_x456_sum_D1_number = RetimeWrapper_30_io_out; // @[package.scala 96:25:@33461.4 package.scala 96:25:@33462.4]
  assign x459_sub_number = x459_sub_1_io_result; // @[Math.scala 195:22:@33452.4 Math.scala 196:14:@33453.4]
  assign _T_1030 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@33525.4 package.scala 96:25:@33526.4]
  assign _T_1032 = io_rr ? _T_1030 : 1'h0; // @[implicits.scala 55:10:@33527.4]
  assign _T_1033 = _T_610 & _T_1032; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 275:194:@33528.4]
  assign x520_x263_D20 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@33513.4 package.scala 96:25:@33514.4]
  assign _T_1034 = _T_1033 & x520_x263_D20; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 275:283:@33529.4]
  assign _T_1035 = _T_1034 & x513_b237_D45; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 275:291:@33530.4]
  assign x269_rdcol_number = x269_rdcol_1_io_result; // @[Math.scala 195:22:@33549.4 Math.scala 196:14:@33550.4]
  assign _T_1052 = $signed(x269_rdcol_number); // @[Math.scala 476:37:@33557.4]
  assign x270 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@33565.4 package.scala 96:25:@33566.4]
  assign x271 = x516_x254_D1 | x270; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 291:59:@33569.4]
  assign _T_1063 = x269_rdcol_number[31]; // @[FixedPoint.scala 50:25:@33576.4]
  assign _T_1067 = _T_1063 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@33578.4]
  assign _T_1068 = x269_rdcol_number[31:16]; // @[FixedPoint.scala 18:52:@33579.4]
  assign _T_1074 = _T_1068 == 16'hffff; // @[Math.scala 451:55:@33581.4]
  assign _T_1075 = x269_rdcol_number[15:0]; // @[FixedPoint.scala 18:52:@33582.4]
  assign _T_1081 = _T_1075 != 16'h0; // @[Math.scala 451:110:@33584.4]
  assign _T_1082 = _T_1074 & _T_1081; // @[Math.scala 451:94:@33585.4]
  assign _T_1084 = {_T_1067,_T_1068}; // @[Cat.scala 30:58:@33587.4]
  assign _T_1096 = $signed(_T_1052) & $signed(32'shffff); // @[Math.scala 406:56:@33597.4]
  assign _T_1097 = $signed(_T_1096); // @[Math.scala 406:56:@33598.4]
  assign x463_sum_number = x463_sum_1_io_result; // @[Math.scala 154:22:@33609.4 Math.scala 155:14:@33610.4]
  assign _T_1104 = x463_sum_number[31]; // @[FixedPoint.scala 50:25:@33614.4]
  assign _T_1108 = _T_1104 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@33616.4]
  assign _T_1109 = x463_sum_number[31:8]; // @[FixedPoint.scala 18:52:@33617.4]
  assign _T_1115 = _T_1109 == 24'hffffff; // @[Math.scala 451:55:@33619.4]
  assign _T_1116 = x463_sum_number[7:0]; // @[FixedPoint.scala 18:52:@33620.4]
  assign _T_1122 = _T_1116 != 8'h0; // @[Math.scala 451:110:@33622.4]
  assign _T_1123 = _T_1115 & _T_1122; // @[Math.scala 451:94:@33623.4]
  assign _T_1127 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@33631.4 package.scala 96:25:@33632.4]
  assign _T_1137 = $signed(x463_sum_number); // @[Math.scala 406:49:@33640.4]
  assign _T_1139 = $signed(_T_1137) & $signed(32'shff); // @[Math.scala 406:56:@33642.4]
  assign _T_1140 = $signed(_T_1139); // @[Math.scala 406:56:@33643.4]
  assign _T_1144 = $signed(RetimeWrapper_37_io_out); // @[package.scala 96:25:@33651.4]
  assign x466_sum_number = x466_sum_1_io_result; // @[Math.scala 154:22:@33663.4 Math.scala 155:14:@33664.4]
  assign _T_1151 = x466_sum_number[31]; // @[FixedPoint.scala 50:25:@33668.4]
  assign _T_1155 = _T_1151 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@33670.4]
  assign _T_1156 = x466_sum_number[31:4]; // @[FixedPoint.scala 18:52:@33671.4]
  assign _T_1162 = _T_1156 == 28'hfffffff; // @[Math.scala 451:55:@33673.4]
  assign _T_1163 = x466_sum_number[3:0]; // @[FixedPoint.scala 18:52:@33674.4]
  assign _T_1169 = _T_1163 != 4'h0; // @[Math.scala 451:110:@33676.4]
  assign _T_1170 = _T_1162 & _T_1169; // @[Math.scala 451:94:@33677.4]
  assign _T_1172 = {_T_1155,_T_1156}; // @[Cat.scala 30:58:@33679.4]
  assign _T_1182 = $signed(x466_sum_number); // @[Math.scala 406:49:@33687.4]
  assign _T_1184 = $signed(_T_1182) & $signed(32'shf); // @[Math.scala 406:56:@33689.4]
  assign _T_1185 = $signed(_T_1184); // @[Math.scala 406:56:@33690.4]
  assign x469_sum_number = x469_sum_1_io_result; // @[Math.scala 154:22:@33701.4 Math.scala 155:14:@33702.4]
  assign _T_1192 = x469_sum_number[31]; // @[FixedPoint.scala 50:25:@33706.4]
  assign _T_1196 = _T_1192 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33708.4]
  assign _T_1197 = x469_sum_number[31:2]; // @[FixedPoint.scala 18:52:@33709.4]
  assign _T_1203 = _T_1197 == 30'h3fffffff; // @[Math.scala 451:55:@33711.4]
  assign _T_1204 = x469_sum_number[1:0]; // @[FixedPoint.scala 18:52:@33712.4]
  assign _T_1210 = _T_1204 != 2'h0; // @[Math.scala 451:110:@33714.4]
  assign _T_1211 = _T_1203 & _T_1210; // @[Math.scala 451:94:@33715.4]
  assign _T_1213 = {_T_1196,_T_1197}; // @[Cat.scala 30:58:@33717.4]
  assign _T_1223 = $signed(x469_sum_number); // @[Math.scala 406:49:@33725.4]
  assign _T_1225 = $signed(_T_1223) & $signed(32'sh3); // @[Math.scala 406:56:@33727.4]
  assign _T_1226 = $signed(_T_1225); // @[Math.scala 406:56:@33728.4]
  assign x472_sum_number = x472_sum_1_io_result; // @[Math.scala 154:22:@33739.4 Math.scala 155:14:@33740.4]
  assign _T_1233 = x472_sum_number[31]; // @[FixedPoint.scala 50:25:@33744.4]
  assign _T_1237 = _T_1233 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33746.4]
  assign _T_1238 = x472_sum_number[31:2]; // @[FixedPoint.scala 18:52:@33747.4]
  assign _T_1244 = _T_1238 == 30'h3fffffff; // @[Math.scala 451:55:@33749.4]
  assign _T_1245 = x472_sum_number[1:0]; // @[FixedPoint.scala 18:52:@33750.4]
  assign _T_1251 = _T_1245 != 2'h0; // @[Math.scala 451:110:@33752.4]
  assign _T_1252 = _T_1244 & _T_1251; // @[Math.scala 451:94:@33753.4]
  assign _T_1254 = {_T_1237,_T_1238}; // @[Cat.scala 30:58:@33755.4]
  assign _T_1264 = $signed(x472_sum_number); // @[Math.scala 406:49:@33763.4]
  assign _T_1266 = $signed(_T_1264) & $signed(32'sh3); // @[Math.scala 406:56:@33765.4]
  assign _T_1267 = $signed(_T_1266); // @[Math.scala 406:56:@33766.4]
  assign x475_sum_number = x475_sum_1_io_result; // @[Math.scala 154:22:@33777.4 Math.scala 155:14:@33778.4]
  assign _T_1274 = x475_sum_number[31]; // @[FixedPoint.scala 50:25:@33782.4]
  assign _T_1278 = _T_1274 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33784.4]
  assign _T_1279 = x475_sum_number[31:2]; // @[FixedPoint.scala 18:52:@33785.4]
  assign _T_1285 = _T_1279 == 30'h3fffffff; // @[Math.scala 451:55:@33787.4]
  assign _T_1286 = x475_sum_number[1:0]; // @[FixedPoint.scala 18:52:@33788.4]
  assign _T_1292 = _T_1286 != 2'h0; // @[Math.scala 451:110:@33790.4]
  assign _T_1293 = _T_1285 & _T_1292; // @[Math.scala 451:94:@33791.4]
  assign _T_1295 = {_T_1278,_T_1279}; // @[Cat.scala 30:58:@33793.4]
  assign _T_1305 = $signed(x475_sum_number); // @[Math.scala 406:49:@33801.4]
  assign _T_1307 = $signed(_T_1305) & $signed(32'sh3); // @[Math.scala 406:56:@33803.4]
  assign _T_1308 = $signed(_T_1307); // @[Math.scala 406:56:@33804.4]
  assign x478_sum_number = x478_sum_1_io_result; // @[Math.scala 154:22:@33815.4 Math.scala 155:14:@33816.4]
  assign _T_1318 = $signed(x478_sum_number); // @[Math.scala 476:37:@33821.4]
  assign x479 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@33829.4 package.scala 96:25:@33830.4]
  assign x521_x478_sum_D1_number = RetimeWrapper_40_io_out; // @[package.scala 96:25:@33864.4 package.scala 96:25:@33865.4]
  assign x481_sub_number = x481_sub_1_io_result; // @[Math.scala 195:22:@33855.4 Math.scala 196:14:@33856.4]
  assign _T_1372 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@33919.4 package.scala 96:25:@33920.4]
  assign _T_1374 = io_rr ? _T_1372 : 1'h0; // @[implicits.scala 55:10:@33921.4]
  assign _T_1375 = _T_610 & _T_1374; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 352:194:@33922.4]
  assign x523_x272_D20 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@33907.4 package.scala 96:25:@33908.4]
  assign _T_1376 = _T_1375 & x523_x272_D20; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 352:283:@33923.4]
  assign _T_1377 = _T_1376 & x513_b237_D45; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 352:291:@33924.4]
  assign x278_rdrow_number = x278_rdrow_1_io_result; // @[Math.scala 195:22:@33943.4 Math.scala 196:14:@33944.4]
  assign _T_1394 = $signed(x278_rdrow_number); // @[Math.scala 406:49:@33950.4]
  assign _T_1396 = $signed(_T_1394) & $signed(32'sh3); // @[Math.scala 406:56:@33952.4]
  assign _T_1397 = $signed(_T_1396); // @[Math.scala 406:56:@33953.4]
  assign x483_number = $unsigned(_T_1397); // @[implicits.scala 133:21:@33954.4]
  assign x280 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@33968.4 package.scala 96:25:@33969.4]
  assign x524_x255_D1 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@33977.4 package.scala 96:25:@33978.4]
  assign x281 = x280 | x524_x255_D1; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 364:24:@33981.4]
  assign _T_1423 = $signed(x483_number); // @[Math.scala 406:49:@33990.4]
  assign _T_1425 = $signed(_T_1423) & $signed(32'sh3); // @[Math.scala 406:56:@33992.4]
  assign _T_1426 = $signed(_T_1425); // @[Math.scala 406:56:@33993.4]
  assign _T_1430 = $signed(RetimeWrapper_46_io_out); // @[package.scala 96:25:@34001.4]
  assign _T_1434 = x483_number[31]; // @[FixedPoint.scala 50:25:@34008.4]
  assign _T_1438 = _T_1434 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34010.4]
  assign _T_1439 = x483_number[31:2]; // @[FixedPoint.scala 18:52:@34011.4]
  assign _T_1445 = _T_1439 == 30'h3fffffff; // @[Math.scala 451:55:@34013.4]
  assign _T_1446 = x483_number[1:0]; // @[FixedPoint.scala 18:52:@34014.4]
  assign _T_1452 = _T_1446 != 2'h0; // @[Math.scala 451:110:@34016.4]
  assign _T_1453 = _T_1445 & _T_1452; // @[Math.scala 451:94:@34017.4]
  assign _T_1457 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@34025.4 package.scala 96:25:@34026.4]
  assign x284_1_number = _T_1453 ? 32'h0 : _T_1457; // @[Math.scala 454:20:@34027.4]
  assign _GEN_2 = {{9'd0}, x284_1_number}; // @[Math.scala 461:32:@34032.4]
  assign _T_1462 = _GEN_2 << 9; // @[Math.scala 461:32:@34032.4]
  assign _GEN_3 = {{7'd0}, x284_1_number}; // @[Math.scala 461:32:@34037.4]
  assign _T_1465 = _GEN_3 << 7; // @[Math.scala 461:32:@34037.4]
  assign _T_1498 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@34114.4 package.scala 96:25:@34115.4]
  assign _T_1500 = io_rr ? _T_1498 : 1'h0; // @[implicits.scala 55:10:@34116.4]
  assign _T_1501 = _T_610 & _T_1500; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 399:194:@34117.4]
  assign x529_x282_D20 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@34102.4 package.scala 96:25:@34103.4]
  assign _T_1502 = _T_1501 & x529_x282_D20; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 399:283:@34118.4]
  assign _T_1503 = _T_1502 & x513_b237_D45; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 399:326:@34119.4]
  assign x289 = x280 | x261; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 403:59:@34130.4]
  assign _T_1532 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@34174.4 package.scala 96:25:@34175.4]
  assign _T_1534 = io_rr ? _T_1532 : 1'h0; // @[implicits.scala 55:10:@34176.4]
  assign _T_1535 = _T_610 & _T_1534; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 418:194:@34177.4]
  assign x531_x290_D20 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@34162.4 package.scala 96:25:@34163.4]
  assign _T_1536 = _T_1535 & x531_x290_D20; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 418:283:@34178.4]
  assign _T_1537 = _T_1536 & x513_b237_D45; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 418:291:@34179.4]
  assign x294 = x280 | x270; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 422:59:@34190.4]
  assign _T_1561 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@34223.4 package.scala 96:25:@34224.4]
  assign _T_1563 = io_rr ? _T_1561 : 1'h0; // @[implicits.scala 55:10:@34225.4]
  assign _T_1564 = _T_610 & _T_1563; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 433:194:@34226.4]
  assign x532_x295_D20 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@34211.4 package.scala 96:25:@34212.4]
  assign _T_1565 = _T_1564 & x532_x295_D20; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 433:283:@34227.4]
  assign _T_1566 = _T_1565 & x513_b237_D45; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 433:291:@34228.4]
  assign x299_rdrow_number = x299_rdrow_1_io_result; // @[Math.scala 195:22:@34247.4 Math.scala 196:14:@34248.4]
  assign _T_1583 = $signed(x299_rdrow_number); // @[Math.scala 406:49:@34254.4]
  assign _T_1585 = $signed(_T_1583) & $signed(32'sh3); // @[Math.scala 406:56:@34256.4]
  assign _T_1586 = $signed(_T_1585); // @[Math.scala 406:56:@34257.4]
  assign x488_number = $unsigned(_T_1586); // @[implicits.scala 133:21:@34258.4]
  assign x301 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@34272.4 package.scala 96:25:@34273.4]
  assign x302 = x301 | x524_x255_D1; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 443:24:@34276.4]
  assign _T_1609 = $signed(x488_number); // @[Math.scala 406:49:@34285.4]
  assign _T_1611 = $signed(_T_1609) & $signed(32'sh3); // @[Math.scala 406:56:@34287.4]
  assign _T_1612 = $signed(_T_1611); // @[Math.scala 406:56:@34288.4]
  assign _T_1616 = $signed(RetimeWrapper_60_io_out); // @[package.scala 96:25:@34296.4]
  assign _T_1620 = x488_number[31]; // @[FixedPoint.scala 50:25:@34303.4]
  assign _T_1624 = _T_1620 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34305.4]
  assign _T_1625 = x488_number[31:2]; // @[FixedPoint.scala 18:52:@34306.4]
  assign _T_1631 = _T_1625 == 30'h3fffffff; // @[Math.scala 451:55:@34308.4]
  assign _T_1632 = x488_number[1:0]; // @[FixedPoint.scala 18:52:@34309.4]
  assign _T_1638 = _T_1632 != 2'h0; // @[Math.scala 451:110:@34311.4]
  assign _T_1639 = _T_1631 & _T_1638; // @[Math.scala 451:94:@34312.4]
  assign _T_1643 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@34320.4 package.scala 96:25:@34321.4]
  assign x305_1_number = _T_1639 ? 32'h0 : _T_1643; // @[Math.scala 454:20:@34322.4]
  assign _GEN_4 = {{9'd0}, x305_1_number}; // @[Math.scala 461:32:@34327.4]
  assign _T_1648 = _GEN_4 << 9; // @[Math.scala 461:32:@34327.4]
  assign _GEN_5 = {{7'd0}, x305_1_number}; // @[Math.scala 461:32:@34332.4]
  assign _T_1651 = _GEN_5 << 7; // @[Math.scala 461:32:@34332.4]
  assign _T_1681 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@34400.4 package.scala 96:25:@34401.4]
  assign _T_1683 = io_rr ? _T_1681 : 1'h0; // @[implicits.scala 55:10:@34402.4]
  assign _T_1684 = _T_610 & _T_1683; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 470:194:@34403.4]
  assign x536_x303_D20 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@34388.4 package.scala 96:25:@34389.4]
  assign _T_1685 = _T_1684 & x536_x303_D20; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 470:283:@34404.4]
  assign _T_1686 = _T_1685 & x513_b237_D45; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 470:291:@34405.4]
  assign x310 = x301 | x261; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 474:24:@34416.4]
  assign _T_1713 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@34458.4 package.scala 96:25:@34459.4]
  assign _T_1715 = io_rr ? _T_1713 : 1'h0; // @[implicits.scala 55:10:@34460.4]
  assign _T_1716 = _T_610 & _T_1715; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 487:194:@34461.4]
  assign x538_x311_D20 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@34446.4 package.scala 96:25:@34447.4]
  assign _T_1717 = _T_1716 & x538_x311_D20; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 487:283:@34462.4]
  assign _T_1718 = _T_1717 & x513_b237_D45; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 487:291:@34463.4]
  assign x315 = x301 | x270; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 491:24:@34474.4]
  assign _T_1742 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@34507.4 package.scala 96:25:@34508.4]
  assign _T_1744 = io_rr ? _T_1742 : 1'h0; // @[implicits.scala 55:10:@34509.4]
  assign _T_1745 = _T_610 & _T_1744; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 502:194:@34510.4]
  assign x539_x316_D20 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@34495.4 package.scala 96:25:@34496.4]
  assign _T_1746 = _T_1745 & x539_x316_D20; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 502:283:@34511.4]
  assign _T_1747 = _T_1746 & x513_b237_D45; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 502:291:@34512.4]
  assign x267_rd_0_number = x241_lb_0_io_rPort_6_output_0; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 271:29:@33516.4 sm_x359_inr_Foreach_SAMPLER_BOX.scala 275:338:@33537.4]
  assign _GEN_6 = {{1'd0}, x267_rd_0_number}; // @[Math.scala 461:32:@34524.4]
  assign _T_1752 = _GEN_6 << 1; // @[Math.scala 461:32:@34524.4]
  assign x287_rd_0_number = x241_lb_0_io_rPort_8_output_0; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 395:29:@34105.4 sm_x359_inr_Foreach_SAMPLER_BOX.scala 399:443:@34126.4]
  assign _GEN_7 = {{1'd0}, x287_rd_0_number}; // @[Math.scala 461:32:@34529.4]
  assign _T_1755 = _GEN_7 << 1; // @[Math.scala 461:32:@34529.4]
  assign x292_rd_0_number = x241_lb_0_io_rPort_2_output_0; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 414:29:@34165.4 sm_x359_inr_Foreach_SAMPLER_BOX.scala 418:408:@34186.4]
  assign _GEN_8 = {{2'd0}, x292_rd_0_number}; // @[Math.scala 461:32:@34534.4]
  assign _T_1758 = _GEN_8 << 2; // @[Math.scala 461:32:@34534.4]
  assign x297_rd_0_number = x241_lb_0_io_rPort_3_output_0; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 429:29:@34214.4 sm_x359_inr_Foreach_SAMPLER_BOX.scala 433:408:@34235.4]
  assign _GEN_9 = {{1'd0}, x297_rd_0_number}; // @[Math.scala 461:32:@34539.4]
  assign _T_1761 = _GEN_9 << 1; // @[Math.scala 461:32:@34539.4]
  assign x313_rd_0_number = x241_lb_0_io_rPort_4_output_0; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 483:29:@34449.4 sm_x359_inr_Foreach_SAMPLER_BOX.scala 487:408:@34470.4]
  assign _GEN_10 = {{1'd0}, x313_rd_0_number}; // @[Math.scala 461:32:@34546.4]
  assign _T_1766 = _GEN_10 << 1; // @[Math.scala 461:32:@34546.4]
  assign _T_1830 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@34730.4 package.scala 96:25:@34731.4]
  assign _T_1832 = io_rr ? _T_1830 : 1'h0; // @[implicits.scala 55:10:@34732.4]
  assign _T_1833 = _T_610 & _T_1832; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 564:167:@34733.4]
  assign _T_1835 = _T_1833 & _T_610; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 564:256:@34735.4]
  assign _T_1836 = _T_1835 & io_sigsIn_backpressure; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 564:275:@34736.4]
  assign x543_b237_D58 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@34692.4 package.scala 96:25:@34693.4]
  assign _T_1837 = _T_1836 & x543_b237_D58; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 564:301:@34737.4]
  assign x541_b238_D58 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@34674.4 package.scala 96:25:@34675.4]
  assign _T_1868 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@34808.4 package.scala 96:25:@34809.4]
  assign _T_1870 = io_rr ? _T_1868 : 1'h0; // @[implicits.scala 55:10:@34810.4]
  assign _T_1871 = _T_610 & _T_1870; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 582:195:@34811.4]
  assign x547_x257_D35 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@34751.4 package.scala 96:25:@34752.4]
  assign _T_1872 = _T_1871 & x547_x257_D35; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 582:284:@34812.4]
  assign x550_b237_D59 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@34778.4 package.scala 96:25:@34779.4]
  assign _T_1873 = _T_1872 & x550_b237_D59; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 582:292:@34813.4]
  assign x548_b238_D59 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@34760.4 package.scala 96:25:@34761.4]
  assign _T_1896 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@34859.4 package.scala 96:25:@34860.4]
  assign _T_1898 = io_rr ? _T_1896 : 1'h0; // @[implicits.scala 55:10:@34861.4]
  assign _T_1899 = _T_610 & _T_1898; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 595:195:@34862.4]
  assign x555_x263_D34 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@34847.4 package.scala 96:25:@34848.4]
  assign _T_1900 = _T_1899 & x555_x263_D34; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 595:284:@34863.4]
  assign _T_1901 = _T_1900 & x550_b237_D59; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 595:292:@34864.4]
  assign _T_1924 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@34910.4 package.scala 96:25:@34911.4]
  assign _T_1926 = io_rr ? _T_1924 : 1'h0; // @[implicits.scala 55:10:@34912.4]
  assign _T_1927 = _T_610 & _T_1926; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 608:195:@34913.4]
  assign x558_x282_D34 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@34898.4 package.scala 96:25:@34899.4]
  assign _T_1928 = _T_1927 & x558_x282_D34; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 608:284:@34914.4]
  assign _T_1929 = _T_1928 & x550_b237_D59; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 608:292:@34915.4]
  assign _T_1949 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@34952.4 package.scala 96:25:@34953.4]
  assign _T_1951 = io_rr ? _T_1949 : 1'h0; // @[implicits.scala 55:10:@34954.4]
  assign _T_1952 = _T_610 & _T_1951; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 619:195:@34955.4]
  assign x560_x290_D34 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@34940.4 package.scala 96:25:@34941.4]
  assign _T_1953 = _T_1952 & x560_x290_D34; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 619:284:@34956.4]
  assign _T_1954 = _T_1953 & x550_b237_D59; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 619:292:@34957.4]
  assign x341_rd_0_number = x242_lb2_0_io_rPort_1_output_0; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 591:29:@34850.4 sm_x359_inr_Foreach_SAMPLER_BOX.scala 595:339:@34871.4]
  assign _GEN_11 = {{1'd0}, x341_rd_0_number}; // @[Math.scala 461:32:@34969.4]
  assign x343_rd_0_number = x242_lb2_0_io_rPort_2_output_0; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 604:29:@34901.4 sm_x359_inr_Foreach_SAMPLER_BOX.scala 608:339:@34922.4]
  assign _GEN_12 = {{2'd0}, x343_rd_0_number}; // @[Math.scala 461:32:@34981.4]
  assign _T_2016 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@35108.4 package.scala 96:25:@35109.4]
  assign _T_2018 = io_rr ? _T_2016 : 1'h0; // @[implicits.scala 55:10:@35110.4]
  assign x563_b237_D73 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@35090.4 package.scala 96:25:@35091.4]
  assign _T_2019 = _T_2018 & x563_b237_D73; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 659:117:@35111.4]
  assign x564_b238_D73 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@35099.4 package.scala 96:25:@35100.4]
  assign _T_2020 = _T_2019 & x564_b238_D73; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 659:123:@35112.4]
  assign x251_sum_number = x251_sum_1_io_result; // @[Math.scala 154:22:@32927.4 Math.scala 155:14:@32928.4]
  assign x504_x435_D13_number = RetimeWrapper_8_io_out; // @[package.scala 96:25:@32945.4 package.scala 96:25:@32946.4]
  assign x506_x413_D21_number = RetimeWrapper_10_io_out; // @[package.scala 96:25:@32963.4 package.scala 96:25:@32964.4]
  assign x512_x435_D37_number = RetimeWrapper_19_io_out; // @[package.scala 96:25:@33076.4 package.scala 96:25:@33077.4]
  assign x514_x413_D45_number = RetimeWrapper_21_io_out; // @[package.scala 96:25:@33094.4 package.scala 96:25:@33095.4]
  assign x515_x251_sum_D24_number = RetimeWrapper_22_io_out; // @[package.scala 96:25:@33103.4 package.scala 96:25:@33104.4]
  assign x266_sum_number = x266_sum_1_io_result; // @[Math.scala 154:22:@33495.4 Math.scala 155:14:@33496.4]
  assign x519_x460_D13_number = RetimeWrapper_32_io_out; // @[package.scala 96:25:@33504.4 package.scala 96:25:@33505.4]
  assign x275_sum_number = x275_sum_1_io_result; // @[Math.scala 154:22:@33889.4 Math.scala 155:14:@33890.4]
  assign x522_x482_D13_number = RetimeWrapper_41_io_out; // @[package.scala 96:25:@33898.4 package.scala 96:25:@33899.4]
  assign x527_x484_D20_number = RetimeWrapper_50_io_out; // @[package.scala 96:25:@34084.4 package.scala 96:25:@34085.4]
  assign x528_x286_sum_D1_number = RetimeWrapper_51_io_out; // @[package.scala 96:25:@34093.4 package.scala 96:25:@34094.4]
  assign x291_sum_number = x291_sum_1_io_result; // @[Math.scala 154:22:@34153.4 Math.scala 155:14:@34154.4]
  assign x296_sum_number = x296_sum_1_io_result; // @[Math.scala 154:22:@34202.4 Math.scala 155:14:@34203.4]
  assign x534_x307_sum_D1_number = RetimeWrapper_63_io_out; // @[package.scala 96:25:@34370.4 package.scala 96:25:@34371.4]
  assign x535_x489_D20_number = RetimeWrapper_64_io_out; // @[package.scala 96:25:@34379.4 package.scala 96:25:@34380.4]
  assign x312_sum_number = x312_sum_1_io_result; // @[Math.scala 154:22:@34437.4 Math.scala 155:14:@34438.4]
  assign x317_sum_number = x317_sum_1_io_result; // @[Math.scala 154:22:@34486.4 Math.scala 155:14:@34487.4]
  assign x542_x435_D50_number = RetimeWrapper_74_io_out; // @[package.scala 96:25:@34683.4 package.scala 96:25:@34684.4]
  assign x544_x413_D58_number = RetimeWrapper_76_io_out; // @[package.scala 96:25:@34701.4 package.scala 96:25:@34702.4]
  assign x546_x251_sum_D37_number = RetimeWrapper_78_io_out; // @[package.scala 96:25:@34719.4 package.scala 96:25:@34720.4]
  assign x549_x435_D51_number = RetimeWrapper_82_io_out; // @[package.scala 96:25:@34769.4 package.scala 96:25:@34770.4]
  assign x551_x413_D59_number = RetimeWrapper_84_io_out; // @[package.scala 96:25:@34787.4 package.scala 96:25:@34788.4]
  assign x552_x251_sum_D38_number = RetimeWrapper_85_io_out; // @[package.scala 96:25:@34796.4 package.scala 96:25:@34797.4]
  assign x553_x460_D27_number = RetimeWrapper_87_io_out; // @[package.scala 96:25:@34829.4 package.scala 96:25:@34830.4]
  assign x554_x266_sum_D14_number = RetimeWrapper_88_io_out; // @[package.scala 96:25:@34838.4 package.scala 96:25:@34839.4]
  assign x556_x484_D34_number = RetimeWrapper_91_io_out; // @[package.scala 96:25:@34880.4 package.scala 96:25:@34881.4]
  assign x557_x286_sum_D15_number = RetimeWrapper_92_io_out; // @[package.scala 96:25:@34889.4 package.scala 96:25:@34890.4]
  assign x559_x291_sum_D14_number = RetimeWrapper_95_io_out; // @[package.scala 96:25:@34931.4 package.scala 96:25:@34932.4]
  assign _T_1961 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@34975.4 package.scala 96:25:@34976.4]
  assign _T_1966 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@34987.4 package.scala 96:25:@34988.4]
  assign io_in_x209_TREADY = _T_211 & _T_213; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 67:22:@32409.4 sm_x359_inr_Foreach_SAMPLER_BOX.scala 69:22:@32417.4]
  assign io_in_x210_TVALID = _T_2020 & io_sigsIn_backpressure; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 659:22:@35114.4]
  assign io_in_x210_TDATA = {{224'd0}, RetimeWrapper_102_io_out}; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 660:24:@35115.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@32387.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@32399.4]
  assign RetimeWrapper_clock = clock; // @[:@32420.4]
  assign RetimeWrapper_reset = reset; // @[:@32421.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32423.4]
  assign RetimeWrapper_io_in = io_in_x209_TDATA[31:0]; // @[package.scala 94:16:@32422.4]
  assign x241_lb_0_clock = clock; // @[:@32430.4]
  assign x241_lb_0_reset = reset; // @[:@32431.4]
  assign x241_lb_0_io_rPort_8_banks_1 = x512_x435_D37_number[1:0]; // @[MemInterfaceType.scala 106:58:@34122.4]
  assign x241_lb_0_io_rPort_8_banks_0 = x527_x484_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@34121.4]
  assign x241_lb_0_io_rPort_8_ofs_0 = x528_x286_sum_D1_number[9:0]; // @[MemInterfaceType.scala 107:54:@34123.4]
  assign x241_lb_0_io_rPort_8_en_0 = _T_1503 & x511_b238_D45; // @[MemInterfaceType.scala 110:79:@34125.4]
  assign x241_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34124.4]
  assign x241_lb_0_io_rPort_7_banks_1 = x512_x435_D37_number[1:0]; // @[MemInterfaceType.scala 106:58:@33123.4]
  assign x241_lb_0_io_rPort_7_banks_0 = x514_x413_D45_number[2:0]; // @[MemInterfaceType.scala 106:58:@33122.4]
  assign x241_lb_0_io_rPort_7_ofs_0 = x515_x251_sum_D24_number[9:0]; // @[MemInterfaceType.scala 107:54:@33124.4]
  assign x241_lb_0_io_rPort_7_en_0 = _T_689 & x511_b238_D45; // @[MemInterfaceType.scala 110:79:@33126.4]
  assign x241_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33125.4]
  assign x241_lb_0_io_rPort_6_banks_1 = x519_x460_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@33533.4]
  assign x241_lb_0_io_rPort_6_banks_0 = x514_x413_D45_number[2:0]; // @[MemInterfaceType.scala 106:58:@33532.4]
  assign x241_lb_0_io_rPort_6_ofs_0 = x266_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@33534.4]
  assign x241_lb_0_io_rPort_6_en_0 = _T_1035 & x511_b238_D45; // @[MemInterfaceType.scala 110:79:@33536.4]
  assign x241_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33535.4]
  assign x241_lb_0_io_rPort_5_banks_1 = x522_x482_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@34515.4]
  assign x241_lb_0_io_rPort_5_banks_0 = x535_x489_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@34514.4]
  assign x241_lb_0_io_rPort_5_ofs_0 = x317_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@34516.4]
  assign x241_lb_0_io_rPort_5_en_0 = _T_1747 & x511_b238_D45; // @[MemInterfaceType.scala 110:79:@34518.4]
  assign x241_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34517.4]
  assign x241_lb_0_io_rPort_4_banks_1 = x519_x460_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@34466.4]
  assign x241_lb_0_io_rPort_4_banks_0 = x535_x489_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@34465.4]
  assign x241_lb_0_io_rPort_4_ofs_0 = x312_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@34467.4]
  assign x241_lb_0_io_rPort_4_en_0 = _T_1718 & x511_b238_D45; // @[MemInterfaceType.scala 110:79:@34469.4]
  assign x241_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34468.4]
  assign x241_lb_0_io_rPort_3_banks_1 = x522_x482_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@34231.4]
  assign x241_lb_0_io_rPort_3_banks_0 = x527_x484_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@34230.4]
  assign x241_lb_0_io_rPort_3_ofs_0 = x296_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@34232.4]
  assign x241_lb_0_io_rPort_3_en_0 = _T_1566 & x511_b238_D45; // @[MemInterfaceType.scala 110:79:@34234.4]
  assign x241_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34233.4]
  assign x241_lb_0_io_rPort_2_banks_1 = x519_x460_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@34182.4]
  assign x241_lb_0_io_rPort_2_banks_0 = x527_x484_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@34181.4]
  assign x241_lb_0_io_rPort_2_ofs_0 = x291_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@34183.4]
  assign x241_lb_0_io_rPort_2_en_0 = _T_1537 & x511_b238_D45; // @[MemInterfaceType.scala 110:79:@34185.4]
  assign x241_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34184.4]
  assign x241_lb_0_io_rPort_1_banks_1 = x512_x435_D37_number[1:0]; // @[MemInterfaceType.scala 106:58:@34408.4]
  assign x241_lb_0_io_rPort_1_banks_0 = x535_x489_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@34407.4]
  assign x241_lb_0_io_rPort_1_ofs_0 = x534_x307_sum_D1_number[9:0]; // @[MemInterfaceType.scala 107:54:@34409.4]
  assign x241_lb_0_io_rPort_1_en_0 = _T_1686 & x511_b238_D45; // @[MemInterfaceType.scala 110:79:@34411.4]
  assign x241_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34410.4]
  assign x241_lb_0_io_rPort_0_banks_1 = x522_x482_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@33927.4]
  assign x241_lb_0_io_rPort_0_banks_0 = x514_x413_D45_number[2:0]; // @[MemInterfaceType.scala 106:58:@33926.4]
  assign x241_lb_0_io_rPort_0_ofs_0 = x275_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@33928.4]
  assign x241_lb_0_io_rPort_0_en_0 = _T_1377 & x511_b238_D45; // @[MemInterfaceType.scala 110:79:@33930.4]
  assign x241_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33929.4]
  assign x241_lb_0_io_wPort_0_banks_1 = x504_x435_D13_number[1:0]; // @[MemInterfaceType.scala 88:58:@32993.4]
  assign x241_lb_0_io_wPort_0_banks_0 = x506_x413_D21_number[2:0]; // @[MemInterfaceType.scala 88:58:@32992.4]
  assign x241_lb_0_io_wPort_0_ofs_0 = x251_sum_number[9:0]; // @[MemInterfaceType.scala 89:54:@32994.4]
  assign x241_lb_0_io_wPort_0_data_0 = RetimeWrapper_11_io_out; // @[MemInterfaceType.scala 90:56:@32995.4]
  assign x241_lb_0_io_wPort_0_en_0 = _T_621 & x503_b238_D21; // @[MemInterfaceType.scala 93:57:@32997.4]
  assign x242_lb2_0_clock = clock; // @[:@32497.4]
  assign x242_lb2_0_reset = reset; // @[:@32498.4]
  assign x242_lb2_0_io_rPort_3_banks_1 = x553_x460_D27_number[1:0]; // @[MemInterfaceType.scala 106:58:@34960.4]
  assign x242_lb2_0_io_rPort_3_banks_0 = x556_x484_D34_number[2:0]; // @[MemInterfaceType.scala 106:58:@34959.4]
  assign x242_lb2_0_io_rPort_3_ofs_0 = x559_x291_sum_D14_number[9:0]; // @[MemInterfaceType.scala 107:54:@34961.4]
  assign x242_lb2_0_io_rPort_3_en_0 = _T_1954 & x548_b238_D59; // @[MemInterfaceType.scala 110:79:@34963.4]
  assign x242_lb2_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34962.4]
  assign x242_lb2_0_io_rPort_2_banks_1 = x549_x435_D51_number[1:0]; // @[MemInterfaceType.scala 106:58:@34918.4]
  assign x242_lb2_0_io_rPort_2_banks_0 = x556_x484_D34_number[2:0]; // @[MemInterfaceType.scala 106:58:@34917.4]
  assign x242_lb2_0_io_rPort_2_ofs_0 = x557_x286_sum_D15_number[9:0]; // @[MemInterfaceType.scala 107:54:@34919.4]
  assign x242_lb2_0_io_rPort_2_en_0 = _T_1929 & x548_b238_D59; // @[MemInterfaceType.scala 110:79:@34921.4]
  assign x242_lb2_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34920.4]
  assign x242_lb2_0_io_rPort_1_banks_1 = x553_x460_D27_number[1:0]; // @[MemInterfaceType.scala 106:58:@34867.4]
  assign x242_lb2_0_io_rPort_1_banks_0 = x551_x413_D59_number[2:0]; // @[MemInterfaceType.scala 106:58:@34866.4]
  assign x242_lb2_0_io_rPort_1_ofs_0 = x554_x266_sum_D14_number[9:0]; // @[MemInterfaceType.scala 107:54:@34868.4]
  assign x242_lb2_0_io_rPort_1_en_0 = _T_1901 & x548_b238_D59; // @[MemInterfaceType.scala 110:79:@34870.4]
  assign x242_lb2_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34869.4]
  assign x242_lb2_0_io_rPort_0_banks_1 = x549_x435_D51_number[1:0]; // @[MemInterfaceType.scala 106:58:@34816.4]
  assign x242_lb2_0_io_rPort_0_banks_0 = x551_x413_D59_number[2:0]; // @[MemInterfaceType.scala 106:58:@34815.4]
  assign x242_lb2_0_io_rPort_0_ofs_0 = x552_x251_sum_D38_number[9:0]; // @[MemInterfaceType.scala 107:54:@34817.4]
  assign x242_lb2_0_io_rPort_0_en_0 = _T_1873 & x548_b238_D59; // @[MemInterfaceType.scala 110:79:@34819.4]
  assign x242_lb2_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34818.4]
  assign x242_lb2_0_io_wPort_0_banks_1 = x542_x435_D50_number[1:0]; // @[MemInterfaceType.scala 88:58:@34740.4]
  assign x242_lb2_0_io_wPort_0_banks_0 = x544_x413_D58_number[2:0]; // @[MemInterfaceType.scala 88:58:@34739.4]
  assign x242_lb2_0_io_wPort_0_ofs_0 = x546_x251_sum_D37_number[9:0]; // @[MemInterfaceType.scala 89:54:@34741.4]
  assign x242_lb2_0_io_wPort_0_data_0 = RetimeWrapper_77_io_out; // @[MemInterfaceType.scala 90:56:@34742.4]
  assign x242_lb2_0_io_wPort_0_en_0 = _T_1837 & x541_b238_D58; // @[MemInterfaceType.scala 93:57:@34744.4]
  assign x416_sum_1_clock = clock; // @[:@32592.4]
  assign x416_sum_1_reset = reset; // @[:@32593.4]
  assign x416_sum_1_io_a = _T_281 ? 32'h0 : _T_283; // @[Math.scala 151:17:@32594.4]
  assign x416_sum_1_io_b = $unsigned(_T_296); // @[Math.scala 152:17:@32595.4]
  assign x416_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@32596.4]
  assign x419_sum_1_clock = clock; // @[:@32630.4]
  assign x419_sum_1_reset = reset; // @[:@32631.4]
  assign x419_sum_1_io_a = _T_322 ? 32'h0 : _T_324; // @[Math.scala 151:17:@32632.4]
  assign x419_sum_1_io_b = $unsigned(_T_337); // @[Math.scala 152:17:@32633.4]
  assign x419_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@32634.4]
  assign x422_sum_1_clock = clock; // @[:@32668.4]
  assign x422_sum_1_reset = reset; // @[:@32669.4]
  assign x422_sum_1_io_a = _T_363 ? 32'h0 : _T_365; // @[Math.scala 151:17:@32670.4]
  assign x422_sum_1_io_b = $unsigned(_T_378); // @[Math.scala 152:17:@32671.4]
  assign x422_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@32672.4]
  assign x425_sum_1_clock = clock; // @[:@32706.4]
  assign x425_sum_1_reset = reset; // @[:@32707.4]
  assign x425_sum_1_io_a = _T_404 ? 32'h0 : _T_406; // @[Math.scala 151:17:@32708.4]
  assign x425_sum_1_io_b = $unsigned(_T_419); // @[Math.scala 152:17:@32709.4]
  assign x425_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@32710.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32729.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32730.4]
  assign RetimeWrapper_1_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@32732.4]
  assign RetimeWrapper_1_io_in = {_T_430,_T_431}; // @[package.scala 94:16:@32731.4]
  assign RetimeWrapper_2_clock = clock; // @[:@32747.4]
  assign RetimeWrapper_2_reset = reset; // @[:@32748.4]
  assign RetimeWrapper_2_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@32751.4]
  assign RetimeWrapper_2_io_in = $unsigned(_T_462); // @[package.scala 94:16:@32750.4]
  assign x428_sum_1_clock = clock; // @[:@32760.4]
  assign x428_sum_1_reset = reset; // @[:@32761.4]
  assign x428_sum_1_io_a = _T_445 ? 32'h0 : _T_449; // @[Math.scala 151:17:@32762.4]
  assign x428_sum_1_io_b = $unsigned(_T_466); // @[Math.scala 152:17:@32763.4]
  assign x428_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@32764.4]
  assign x431_sum_1_clock = clock; // @[:@32798.4]
  assign x431_sum_1_reset = reset; // @[:@32799.4]
  assign x431_sum_1_io_a = _T_492 ? 32'h0 : _T_494; // @[Math.scala 151:17:@32800.4]
  assign x431_sum_1_io_b = $unsigned(_T_507); // @[Math.scala 152:17:@32801.4]
  assign x431_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@32802.4]
  assign x434_sub_1_clock = clock; // @[:@32824.4]
  assign x434_sub_1_reset = reset; // @[:@32825.4]
  assign x434_sub_1_io_a = x431_sum_1_io_result; // @[Math.scala 192:17:@32826.4]
  assign x434_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@32827.4]
  assign x434_sub_1_io_flow = io_in_x210_TREADY; // @[Math.scala 194:20:@32828.4]
  assign RetimeWrapper_3_clock = clock; // @[:@32834.4]
  assign RetimeWrapper_3_reset = reset; // @[:@32835.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32837.4]
  assign RetimeWrapper_3_io_in = $signed(_T_517) < $signed(32'sh3); // @[package.scala 94:16:@32836.4]
  assign RetimeWrapper_4_clock = clock; // @[:@32843.4]
  assign RetimeWrapper_4_reset = reset; // @[:@32844.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32846.4]
  assign RetimeWrapper_4_io_in = $signed(_T_517) < $signed(32'sh6); // @[package.scala 94:16:@32845.4]
  assign RetimeWrapper_5_clock = clock; // @[:@32852.4]
  assign RetimeWrapper_5_reset = reset; // @[:@32853.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32855.4]
  assign RetimeWrapper_5_io_in = x431_sum_1_io_result; // @[package.scala 94:16:@32854.4]
  assign x438_sum_1_clock = clock; // @[:@32891.4]
  assign x438_sum_1_reset = reset; // @[:@32892.4]
  assign x438_sum_1_io_a = _T_574[31:0]; // @[Math.scala 151:17:@32893.4]
  assign x438_sum_1_io_b = _T_577[31:0]; // @[Math.scala 152:17:@32894.4]
  assign x438_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@32895.4]
  assign x250_div_1_clock = clock; // @[:@32903.4]
  assign x250_div_1_io_a = __1_io_result; // @[Math.scala 328:17:@32905.4]
  assign x250_div_1_io_flow = io_in_x210_TREADY; // @[Math.scala 330:20:@32907.4]
  assign RetimeWrapper_6_clock = clock; // @[:@32913.4]
  assign RetimeWrapper_6_reset = reset; // @[:@32914.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32916.4]
  assign RetimeWrapper_6_io_in = x438_sum_1_io_result; // @[package.scala 94:16:@32915.4]
  assign x251_sum_1_clock = clock; // @[:@32922.4]
  assign x251_sum_1_reset = reset; // @[:@32923.4]
  assign x251_sum_1_io_a = RetimeWrapper_6_io_out; // @[Math.scala 151:17:@32924.4]
  assign x251_sum_1_io_b = x250_div_1_io_result; // @[Math.scala 152:17:@32925.4]
  assign x251_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@32926.4]
  assign RetimeWrapper_7_clock = clock; // @[:@32932.4]
  assign RetimeWrapper_7_reset = reset; // @[:@32933.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32935.4]
  assign RetimeWrapper_7_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@32934.4]
  assign RetimeWrapper_8_clock = clock; // @[:@32941.4]
  assign RetimeWrapper_8_reset = reset; // @[:@32942.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32944.4]
  assign RetimeWrapper_8_io_in = x499_x432_D1 ? x501_x431_sum_D1_number : x434_sub_number; // @[package.scala 94:16:@32943.4]
  assign RetimeWrapper_9_clock = clock; // @[:@32950.4]
  assign RetimeWrapper_9_reset = reset; // @[:@32951.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32953.4]
  assign RetimeWrapper_9_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@32952.4]
  assign RetimeWrapper_10_clock = clock; // @[:@32959.4]
  assign RetimeWrapper_10_reset = reset; // @[:@32960.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32962.4]
  assign RetimeWrapper_10_io_in = $unsigned(_T_258); // @[package.scala 94:16:@32961.4]
  assign RetimeWrapper_11_clock = clock; // @[:@32968.4]
  assign RetimeWrapper_11_reset = reset; // @[:@32969.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32971.4]
  assign RetimeWrapper_11_io_in = RetimeWrapper_io_out; // @[package.scala 94:16:@32970.4]
  assign RetimeWrapper_12_clock = clock; // @[:@32979.4]
  assign RetimeWrapper_12_reset = reset; // @[:@32980.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32982.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32981.4]
  assign RetimeWrapper_13_clock = clock; // @[:@33000.4]
  assign RetimeWrapper_13_reset = reset; // @[:@33001.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33003.4]
  assign RetimeWrapper_13_io_in = __io_result; // @[package.scala 94:16:@33002.4]
  assign RetimeWrapper_14_clock = clock; // @[:@33016.4]
  assign RetimeWrapper_14_reset = reset; // @[:@33017.4]
  assign RetimeWrapper_14_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@33019.4]
  assign RetimeWrapper_14_io_in = $signed(_T_633) < $signed(32'sh0); // @[package.scala 94:16:@33018.4]
  assign RetimeWrapper_15_clock = clock; // @[:@33025.4]
  assign RetimeWrapper_15_reset = reset; // @[:@33026.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33028.4]
  assign RetimeWrapper_15_io_in = __1_io_result; // @[package.scala 94:16:@33027.4]
  assign RetimeWrapper_16_clock = clock; // @[:@33039.4]
  assign RetimeWrapper_16_reset = reset; // @[:@33040.4]
  assign RetimeWrapper_16_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@33042.4]
  assign RetimeWrapper_16_io_in = $signed(_T_646) < $signed(32'sh0); // @[package.scala 94:16:@33041.4]
  assign RetimeWrapper_17_clock = clock; // @[:@33054.4]
  assign RetimeWrapper_17_reset = reset; // @[:@33055.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33057.4]
  assign RetimeWrapper_17_io_in = ~ x256; // @[package.scala 94:16:@33056.4]
  assign RetimeWrapper_18_clock = clock; // @[:@33063.4]
  assign RetimeWrapper_18_reset = reset; // @[:@33064.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33066.4]
  assign RetimeWrapper_18_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@33065.4]
  assign RetimeWrapper_19_clock = clock; // @[:@33072.4]
  assign RetimeWrapper_19_reset = reset; // @[:@33073.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33075.4]
  assign RetimeWrapper_19_io_in = x499_x432_D1 ? x501_x431_sum_D1_number : x434_sub_number; // @[package.scala 94:16:@33074.4]
  assign RetimeWrapper_20_clock = clock; // @[:@33081.4]
  assign RetimeWrapper_20_reset = reset; // @[:@33082.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33084.4]
  assign RetimeWrapper_20_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@33083.4]
  assign RetimeWrapper_21_clock = clock; // @[:@33090.4]
  assign RetimeWrapper_21_reset = reset; // @[:@33091.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33093.4]
  assign RetimeWrapper_21_io_in = $unsigned(_T_258); // @[package.scala 94:16:@33092.4]
  assign RetimeWrapper_22_clock = clock; // @[:@33099.4]
  assign RetimeWrapper_22_reset = reset; // @[:@33100.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33102.4]
  assign RetimeWrapper_22_io_in = x251_sum_1_io_result; // @[package.scala 94:16:@33101.4]
  assign RetimeWrapper_23_clock = clock; // @[:@33111.4]
  assign RetimeWrapper_23_reset = reset; // @[:@33112.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33114.4]
  assign RetimeWrapper_23_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33113.4]
  assign x260_rdcol_1_clock = clock; // @[:@33134.4]
  assign x260_rdcol_1_reset = reset; // @[:@33135.4]
  assign x260_rdcol_1_io_a = RetimeWrapper_15_io_out; // @[Math.scala 192:17:@33136.4]
  assign x260_rdcol_1_io_b = 32'h1; // @[Math.scala 193:17:@33137.4]
  assign x260_rdcol_1_io_flow = io_in_x210_TREADY; // @[Math.scala 194:20:@33138.4]
  assign RetimeWrapper_24_clock = clock; // @[:@33149.4]
  assign RetimeWrapper_24_reset = reset; // @[:@33150.4]
  assign RetimeWrapper_24_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@33152.4]
  assign RetimeWrapper_24_io_in = $signed(_T_704) < $signed(32'sh0); // @[package.scala 94:16:@33151.4]
  assign RetimeWrapper_25_clock = clock; // @[:@33158.4]
  assign RetimeWrapper_25_reset = reset; // @[:@33159.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33161.4]
  assign RetimeWrapper_25_io_in = RetimeWrapper_14_io_out; // @[package.scala 94:16:@33160.4]
  assign x441_sum_1_clock = clock; // @[:@33201.4]
  assign x441_sum_1_reset = reset; // @[:@33202.4]
  assign x441_sum_1_io_a = _T_737 ? 32'h0 : _T_739; // @[Math.scala 151:17:@33203.4]
  assign x441_sum_1_io_b = $unsigned(_T_752); // @[Math.scala 152:17:@33204.4]
  assign x441_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@33205.4]
  assign RetimeWrapper_26_clock = clock; // @[:@33224.4]
  assign RetimeWrapper_26_reset = reset; // @[:@33225.4]
  assign RetimeWrapper_26_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@33227.4]
  assign RetimeWrapper_26_io_in = {_T_763,_T_764}; // @[package.scala 94:16:@33226.4]
  assign RetimeWrapper_27_clock = clock; // @[:@33242.4]
  assign RetimeWrapper_27_reset = reset; // @[:@33243.4]
  assign RetimeWrapper_27_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@33246.4]
  assign RetimeWrapper_27_io_in = $unsigned(_T_795); // @[package.scala 94:16:@33245.4]
  assign x444_sum_1_clock = clock; // @[:@33255.4]
  assign x444_sum_1_reset = reset; // @[:@33256.4]
  assign x444_sum_1_io_a = _T_778 ? 32'h0 : _T_782; // @[Math.scala 151:17:@33257.4]
  assign x444_sum_1_io_b = $unsigned(_T_799); // @[Math.scala 152:17:@33258.4]
  assign x444_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@33259.4]
  assign x447_sum_1_clock = clock; // @[:@33293.4]
  assign x447_sum_1_reset = reset; // @[:@33294.4]
  assign x447_sum_1_io_a = _T_825 ? 32'h0 : _T_827; // @[Math.scala 151:17:@33295.4]
  assign x447_sum_1_io_b = $unsigned(_T_840); // @[Math.scala 152:17:@33296.4]
  assign x447_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@33297.4]
  assign x450_sum_1_clock = clock; // @[:@33331.4]
  assign x450_sum_1_reset = reset; // @[:@33332.4]
  assign x450_sum_1_io_a = _T_866 ? 32'h0 : _T_868; // @[Math.scala 151:17:@33333.4]
  assign x450_sum_1_io_b = $unsigned(_T_881); // @[Math.scala 152:17:@33334.4]
  assign x450_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@33335.4]
  assign x453_sum_1_clock = clock; // @[:@33369.4]
  assign x453_sum_1_reset = reset; // @[:@33370.4]
  assign x453_sum_1_io_a = _T_907 ? 32'h0 : _T_909; // @[Math.scala 151:17:@33371.4]
  assign x453_sum_1_io_b = $unsigned(_T_922); // @[Math.scala 152:17:@33372.4]
  assign x453_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@33373.4]
  assign x456_sum_1_clock = clock; // @[:@33407.4]
  assign x456_sum_1_reset = reset; // @[:@33408.4]
  assign x456_sum_1_io_a = _T_948 ? 32'h0 : _T_950; // @[Math.scala 151:17:@33409.4]
  assign x456_sum_1_io_b = $unsigned(_T_963); // @[Math.scala 152:17:@33410.4]
  assign x456_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@33411.4]
  assign RetimeWrapper_28_clock = clock; // @[:@33422.4]
  assign RetimeWrapper_28_reset = reset; // @[:@33423.4]
  assign RetimeWrapper_28_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@33425.4]
  assign RetimeWrapper_28_io_in = $signed(_T_973) < $signed(32'sh3); // @[package.scala 94:16:@33424.4]
  assign RetimeWrapper_29_clock = clock; // @[:@33436.4]
  assign RetimeWrapper_29_reset = reset; // @[:@33437.4]
  assign RetimeWrapper_29_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@33439.4]
  assign RetimeWrapper_29_io_in = $signed(_T_973) < $signed(32'sh6); // @[package.scala 94:16:@33438.4]
  assign x459_sub_1_clock = clock; // @[:@33447.4]
  assign x459_sub_1_reset = reset; // @[:@33448.4]
  assign x459_sub_1_io_a = x456_sum_1_io_result; // @[Math.scala 192:17:@33449.4]
  assign x459_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@33450.4]
  assign x459_sub_1_io_flow = io_in_x210_TREADY; // @[Math.scala 194:20:@33451.4]
  assign RetimeWrapper_30_clock = clock; // @[:@33457.4]
  assign RetimeWrapper_30_reset = reset; // @[:@33458.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33460.4]
  assign RetimeWrapper_30_io_in = x456_sum_1_io_result; // @[package.scala 94:16:@33459.4]
  assign x265_div_1_clock = clock; // @[:@33471.4]
  assign x265_div_1_io_a = x260_rdcol_1_io_result; // @[Math.scala 328:17:@33473.4]
  assign x265_div_1_io_flow = io_in_x210_TREADY; // @[Math.scala 330:20:@33475.4]
  assign RetimeWrapper_31_clock = clock; // @[:@33481.4]
  assign RetimeWrapper_31_reset = reset; // @[:@33482.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33484.4]
  assign RetimeWrapper_31_io_in = x438_sum_1_io_result; // @[package.scala 94:16:@33483.4]
  assign x266_sum_1_clock = clock; // @[:@33490.4]
  assign x266_sum_1_reset = reset; // @[:@33491.4]
  assign x266_sum_1_io_a = RetimeWrapper_31_io_out; // @[Math.scala 151:17:@33492.4]
  assign x266_sum_1_io_b = x265_div_1_io_result; // @[Math.scala 152:17:@33493.4]
  assign x266_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@33494.4]
  assign RetimeWrapper_32_clock = clock; // @[:@33500.4]
  assign RetimeWrapper_32_reset = reset; // @[:@33501.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33503.4]
  assign RetimeWrapper_32_io_in = x457 ? x517_x456_sum_D1_number : x459_sub_number; // @[package.scala 94:16:@33502.4]
  assign RetimeWrapper_33_clock = clock; // @[:@33509.4]
  assign RetimeWrapper_33_reset = reset; // @[:@33510.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33512.4]
  assign RetimeWrapper_33_io_in = ~ x262; // @[package.scala 94:16:@33511.4]
  assign RetimeWrapper_34_clock = clock; // @[:@33521.4]
  assign RetimeWrapper_34_reset = reset; // @[:@33522.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33524.4]
  assign RetimeWrapper_34_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33523.4]
  assign x269_rdcol_1_clock = clock; // @[:@33544.4]
  assign x269_rdcol_1_reset = reset; // @[:@33545.4]
  assign x269_rdcol_1_io_a = RetimeWrapper_15_io_out; // @[Math.scala 192:17:@33546.4]
  assign x269_rdcol_1_io_b = 32'h2; // @[Math.scala 193:17:@33547.4]
  assign x269_rdcol_1_io_flow = io_in_x210_TREADY; // @[Math.scala 194:20:@33548.4]
  assign RetimeWrapper_35_clock = clock; // @[:@33561.4]
  assign RetimeWrapper_35_reset = reset; // @[:@33562.4]
  assign RetimeWrapper_35_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@33564.4]
  assign RetimeWrapper_35_io_in = $signed(_T_1052) < $signed(32'sh0); // @[package.scala 94:16:@33563.4]
  assign x463_sum_1_clock = clock; // @[:@33604.4]
  assign x463_sum_1_reset = reset; // @[:@33605.4]
  assign x463_sum_1_io_a = _T_1082 ? 32'h0 : _T_1084; // @[Math.scala 151:17:@33606.4]
  assign x463_sum_1_io_b = $unsigned(_T_1097); // @[Math.scala 152:17:@33607.4]
  assign x463_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@33608.4]
  assign RetimeWrapper_36_clock = clock; // @[:@33627.4]
  assign RetimeWrapper_36_reset = reset; // @[:@33628.4]
  assign RetimeWrapper_36_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@33630.4]
  assign RetimeWrapper_36_io_in = {_T_1108,_T_1109}; // @[package.scala 94:16:@33629.4]
  assign RetimeWrapper_37_clock = clock; // @[:@33645.4]
  assign RetimeWrapper_37_reset = reset; // @[:@33646.4]
  assign RetimeWrapper_37_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@33649.4]
  assign RetimeWrapper_37_io_in = $unsigned(_T_1140); // @[package.scala 94:16:@33648.4]
  assign x466_sum_1_clock = clock; // @[:@33658.4]
  assign x466_sum_1_reset = reset; // @[:@33659.4]
  assign x466_sum_1_io_a = _T_1123 ? 32'h0 : _T_1127; // @[Math.scala 151:17:@33660.4]
  assign x466_sum_1_io_b = $unsigned(_T_1144); // @[Math.scala 152:17:@33661.4]
  assign x466_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@33662.4]
  assign x469_sum_1_clock = clock; // @[:@33696.4]
  assign x469_sum_1_reset = reset; // @[:@33697.4]
  assign x469_sum_1_io_a = _T_1170 ? 32'h0 : _T_1172; // @[Math.scala 151:17:@33698.4]
  assign x469_sum_1_io_b = $unsigned(_T_1185); // @[Math.scala 152:17:@33699.4]
  assign x469_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@33700.4]
  assign x472_sum_1_clock = clock; // @[:@33734.4]
  assign x472_sum_1_reset = reset; // @[:@33735.4]
  assign x472_sum_1_io_a = _T_1211 ? 32'h0 : _T_1213; // @[Math.scala 151:17:@33736.4]
  assign x472_sum_1_io_b = $unsigned(_T_1226); // @[Math.scala 152:17:@33737.4]
  assign x472_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@33738.4]
  assign x475_sum_1_clock = clock; // @[:@33772.4]
  assign x475_sum_1_reset = reset; // @[:@33773.4]
  assign x475_sum_1_io_a = _T_1252 ? 32'h0 : _T_1254; // @[Math.scala 151:17:@33774.4]
  assign x475_sum_1_io_b = $unsigned(_T_1267); // @[Math.scala 152:17:@33775.4]
  assign x475_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@33776.4]
  assign x478_sum_1_clock = clock; // @[:@33810.4]
  assign x478_sum_1_reset = reset; // @[:@33811.4]
  assign x478_sum_1_io_a = _T_1293 ? 32'h0 : _T_1295; // @[Math.scala 151:17:@33812.4]
  assign x478_sum_1_io_b = $unsigned(_T_1308); // @[Math.scala 152:17:@33813.4]
  assign x478_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@33814.4]
  assign RetimeWrapper_38_clock = clock; // @[:@33825.4]
  assign RetimeWrapper_38_reset = reset; // @[:@33826.4]
  assign RetimeWrapper_38_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@33828.4]
  assign RetimeWrapper_38_io_in = $signed(_T_1318) < $signed(32'sh3); // @[package.scala 94:16:@33827.4]
  assign RetimeWrapper_39_clock = clock; // @[:@33839.4]
  assign RetimeWrapper_39_reset = reset; // @[:@33840.4]
  assign RetimeWrapper_39_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@33842.4]
  assign RetimeWrapper_39_io_in = $signed(_T_1318) < $signed(32'sh6); // @[package.scala 94:16:@33841.4]
  assign x481_sub_1_clock = clock; // @[:@33850.4]
  assign x481_sub_1_reset = reset; // @[:@33851.4]
  assign x481_sub_1_io_a = x478_sum_1_io_result; // @[Math.scala 192:17:@33852.4]
  assign x481_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@33853.4]
  assign x481_sub_1_io_flow = io_in_x210_TREADY; // @[Math.scala 194:20:@33854.4]
  assign RetimeWrapper_40_clock = clock; // @[:@33860.4]
  assign RetimeWrapper_40_reset = reset; // @[:@33861.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33863.4]
  assign RetimeWrapper_40_io_in = x478_sum_1_io_result; // @[package.scala 94:16:@33862.4]
  assign x274_div_1_clock = clock; // @[:@33874.4]
  assign x274_div_1_io_a = x269_rdcol_1_io_result; // @[Math.scala 328:17:@33876.4]
  assign x274_div_1_io_flow = io_in_x210_TREADY; // @[Math.scala 330:20:@33878.4]
  assign x275_sum_1_clock = clock; // @[:@33884.4]
  assign x275_sum_1_reset = reset; // @[:@33885.4]
  assign x275_sum_1_io_a = RetimeWrapper_31_io_out; // @[Math.scala 151:17:@33886.4]
  assign x275_sum_1_io_b = x274_div_1_io_result; // @[Math.scala 152:17:@33887.4]
  assign x275_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@33888.4]
  assign RetimeWrapper_41_clock = clock; // @[:@33894.4]
  assign RetimeWrapper_41_reset = reset; // @[:@33895.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33897.4]
  assign RetimeWrapper_41_io_in = x479 ? x521_x478_sum_D1_number : x481_sub_number; // @[package.scala 94:16:@33896.4]
  assign RetimeWrapper_42_clock = clock; // @[:@33903.4]
  assign RetimeWrapper_42_reset = reset; // @[:@33904.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33906.4]
  assign RetimeWrapper_42_io_in = ~ x271; // @[package.scala 94:16:@33905.4]
  assign RetimeWrapper_43_clock = clock; // @[:@33915.4]
  assign RetimeWrapper_43_reset = reset; // @[:@33916.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33918.4]
  assign RetimeWrapper_43_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33917.4]
  assign x278_rdrow_1_clock = clock; // @[:@33938.4]
  assign x278_rdrow_1_reset = reset; // @[:@33939.4]
  assign x278_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@33940.4]
  assign x278_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@33941.4]
  assign x278_rdrow_1_io_flow = io_in_x210_TREADY; // @[Math.scala 194:20:@33942.4]
  assign RetimeWrapper_44_clock = clock; // @[:@33964.4]
  assign RetimeWrapper_44_reset = reset; // @[:@33965.4]
  assign RetimeWrapper_44_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@33967.4]
  assign RetimeWrapper_44_io_in = $signed(_T_1394) < $signed(32'sh0); // @[package.scala 94:16:@33966.4]
  assign RetimeWrapper_45_clock = clock; // @[:@33973.4]
  assign RetimeWrapper_45_reset = reset; // @[:@33974.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33976.4]
  assign RetimeWrapper_45_io_in = RetimeWrapper_16_io_out; // @[package.scala 94:16:@33975.4]
  assign RetimeWrapper_46_clock = clock; // @[:@33995.4]
  assign RetimeWrapper_46_reset = reset; // @[:@33996.4]
  assign RetimeWrapper_46_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@33999.4]
  assign RetimeWrapper_46_io_in = $unsigned(_T_1426); // @[package.scala 94:16:@33998.4]
  assign RetimeWrapper_47_clock = clock; // @[:@34021.4]
  assign RetimeWrapper_47_reset = reset; // @[:@34022.4]
  assign RetimeWrapper_47_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@34024.4]
  assign RetimeWrapper_47_io_in = {_T_1438,_T_1439}; // @[package.scala 94:16:@34023.4]
  assign x487_sum_1_clock = clock; // @[:@34042.4]
  assign x487_sum_1_reset = reset; // @[:@34043.4]
  assign x487_sum_1_io_a = _T_1462[31:0]; // @[Math.scala 151:17:@34044.4]
  assign x487_sum_1_io_b = _T_1465[31:0]; // @[Math.scala 152:17:@34045.4]
  assign x487_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34046.4]
  assign RetimeWrapper_48_clock = clock; // @[:@34052.4]
  assign RetimeWrapper_48_reset = reset; // @[:@34053.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34055.4]
  assign RetimeWrapper_48_io_in = x250_div_1_io_result; // @[package.scala 94:16:@34054.4]
  assign RetimeWrapper_49_clock = clock; // @[:@34061.4]
  assign RetimeWrapper_49_reset = reset; // @[:@34062.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34064.4]
  assign RetimeWrapper_49_io_in = x487_sum_1_io_result; // @[package.scala 94:16:@34063.4]
  assign x286_sum_1_clock = clock; // @[:@34070.4]
  assign x286_sum_1_reset = reset; // @[:@34071.4]
  assign x286_sum_1_io_a = RetimeWrapper_49_io_out; // @[Math.scala 151:17:@34072.4]
  assign x286_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@34073.4]
  assign x286_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34074.4]
  assign RetimeWrapper_50_clock = clock; // @[:@34080.4]
  assign RetimeWrapper_50_reset = reset; // @[:@34081.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34083.4]
  assign RetimeWrapper_50_io_in = $unsigned(_T_1430); // @[package.scala 94:16:@34082.4]
  assign RetimeWrapper_51_clock = clock; // @[:@34089.4]
  assign RetimeWrapper_51_reset = reset; // @[:@34090.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34092.4]
  assign RetimeWrapper_51_io_in = x286_sum_1_io_result; // @[package.scala 94:16:@34091.4]
  assign RetimeWrapper_52_clock = clock; // @[:@34098.4]
  assign RetimeWrapper_52_reset = reset; // @[:@34099.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34101.4]
  assign RetimeWrapper_52_io_in = ~ x281; // @[package.scala 94:16:@34100.4]
  assign RetimeWrapper_53_clock = clock; // @[:@34110.4]
  assign RetimeWrapper_53_reset = reset; // @[:@34111.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34113.4]
  assign RetimeWrapper_53_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34112.4]
  assign RetimeWrapper_54_clock = clock; // @[:@34137.4]
  assign RetimeWrapper_54_reset = reset; // @[:@34138.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34140.4]
  assign RetimeWrapper_54_io_in = x487_sum_1_io_result; // @[package.scala 94:16:@34139.4]
  assign x291_sum_1_clock = clock; // @[:@34148.4]
  assign x291_sum_1_reset = reset; // @[:@34149.4]
  assign x291_sum_1_io_a = RetimeWrapper_54_io_out; // @[Math.scala 151:17:@34150.4]
  assign x291_sum_1_io_b = x265_div_1_io_result; // @[Math.scala 152:17:@34151.4]
  assign x291_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34152.4]
  assign RetimeWrapper_55_clock = clock; // @[:@34158.4]
  assign RetimeWrapper_55_reset = reset; // @[:@34159.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34161.4]
  assign RetimeWrapper_55_io_in = ~ x289; // @[package.scala 94:16:@34160.4]
  assign RetimeWrapper_56_clock = clock; // @[:@34170.4]
  assign RetimeWrapper_56_reset = reset; // @[:@34171.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34173.4]
  assign RetimeWrapper_56_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34172.4]
  assign x296_sum_1_clock = clock; // @[:@34197.4]
  assign x296_sum_1_reset = reset; // @[:@34198.4]
  assign x296_sum_1_io_a = RetimeWrapper_54_io_out; // @[Math.scala 151:17:@34199.4]
  assign x296_sum_1_io_b = x274_div_1_io_result; // @[Math.scala 152:17:@34200.4]
  assign x296_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34201.4]
  assign RetimeWrapper_57_clock = clock; // @[:@34207.4]
  assign RetimeWrapper_57_reset = reset; // @[:@34208.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34210.4]
  assign RetimeWrapper_57_io_in = ~ x294; // @[package.scala 94:16:@34209.4]
  assign RetimeWrapper_58_clock = clock; // @[:@34219.4]
  assign RetimeWrapper_58_reset = reset; // @[:@34220.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34222.4]
  assign RetimeWrapper_58_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34221.4]
  assign x299_rdrow_1_clock = clock; // @[:@34242.4]
  assign x299_rdrow_1_reset = reset; // @[:@34243.4]
  assign x299_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@34244.4]
  assign x299_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@34245.4]
  assign x299_rdrow_1_io_flow = io_in_x210_TREADY; // @[Math.scala 194:20:@34246.4]
  assign RetimeWrapper_59_clock = clock; // @[:@34268.4]
  assign RetimeWrapper_59_reset = reset; // @[:@34269.4]
  assign RetimeWrapper_59_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@34271.4]
  assign RetimeWrapper_59_io_in = $signed(_T_1583) < $signed(32'sh0); // @[package.scala 94:16:@34270.4]
  assign RetimeWrapper_60_clock = clock; // @[:@34290.4]
  assign RetimeWrapper_60_reset = reset; // @[:@34291.4]
  assign RetimeWrapper_60_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@34294.4]
  assign RetimeWrapper_60_io_in = $unsigned(_T_1612); // @[package.scala 94:16:@34293.4]
  assign RetimeWrapper_61_clock = clock; // @[:@34316.4]
  assign RetimeWrapper_61_reset = reset; // @[:@34317.4]
  assign RetimeWrapper_61_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@34319.4]
  assign RetimeWrapper_61_io_in = {_T_1624,_T_1625}; // @[package.scala 94:16:@34318.4]
  assign x492_sum_1_clock = clock; // @[:@34337.4]
  assign x492_sum_1_reset = reset; // @[:@34338.4]
  assign x492_sum_1_io_a = _T_1648[31:0]; // @[Math.scala 151:17:@34339.4]
  assign x492_sum_1_io_b = _T_1651[31:0]; // @[Math.scala 152:17:@34340.4]
  assign x492_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34341.4]
  assign RetimeWrapper_62_clock = clock; // @[:@34347.4]
  assign RetimeWrapper_62_reset = reset; // @[:@34348.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34350.4]
  assign RetimeWrapper_62_io_in = x492_sum_1_io_result; // @[package.scala 94:16:@34349.4]
  assign x307_sum_1_clock = clock; // @[:@34356.4]
  assign x307_sum_1_reset = reset; // @[:@34357.4]
  assign x307_sum_1_io_a = RetimeWrapper_62_io_out; // @[Math.scala 151:17:@34358.4]
  assign x307_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@34359.4]
  assign x307_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34360.4]
  assign RetimeWrapper_63_clock = clock; // @[:@34366.4]
  assign RetimeWrapper_63_reset = reset; // @[:@34367.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34369.4]
  assign RetimeWrapper_63_io_in = x307_sum_1_io_result; // @[package.scala 94:16:@34368.4]
  assign RetimeWrapper_64_clock = clock; // @[:@34375.4]
  assign RetimeWrapper_64_reset = reset; // @[:@34376.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34378.4]
  assign RetimeWrapper_64_io_in = $unsigned(_T_1616); // @[package.scala 94:16:@34377.4]
  assign RetimeWrapper_65_clock = clock; // @[:@34384.4]
  assign RetimeWrapper_65_reset = reset; // @[:@34385.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34387.4]
  assign RetimeWrapper_65_io_in = ~ x302; // @[package.scala 94:16:@34386.4]
  assign RetimeWrapper_66_clock = clock; // @[:@34396.4]
  assign RetimeWrapper_66_reset = reset; // @[:@34397.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34399.4]
  assign RetimeWrapper_66_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34398.4]
  assign RetimeWrapper_67_clock = clock; // @[:@34423.4]
  assign RetimeWrapper_67_reset = reset; // @[:@34424.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34426.4]
  assign RetimeWrapper_67_io_in = x492_sum_1_io_result; // @[package.scala 94:16:@34425.4]
  assign x312_sum_1_clock = clock; // @[:@34432.4]
  assign x312_sum_1_reset = reset; // @[:@34433.4]
  assign x312_sum_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@34434.4]
  assign x312_sum_1_io_b = x265_div_1_io_result; // @[Math.scala 152:17:@34435.4]
  assign x312_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34436.4]
  assign RetimeWrapper_68_clock = clock; // @[:@34442.4]
  assign RetimeWrapper_68_reset = reset; // @[:@34443.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34445.4]
  assign RetimeWrapper_68_io_in = ~ x310; // @[package.scala 94:16:@34444.4]
  assign RetimeWrapper_69_clock = clock; // @[:@34454.4]
  assign RetimeWrapper_69_reset = reset; // @[:@34455.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34457.4]
  assign RetimeWrapper_69_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34456.4]
  assign x317_sum_1_clock = clock; // @[:@34481.4]
  assign x317_sum_1_reset = reset; // @[:@34482.4]
  assign x317_sum_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@34483.4]
  assign x317_sum_1_io_b = x274_div_1_io_result; // @[Math.scala 152:17:@34484.4]
  assign x317_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34485.4]
  assign RetimeWrapper_70_clock = clock; // @[:@34491.4]
  assign RetimeWrapper_70_reset = reset; // @[:@34492.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34494.4]
  assign RetimeWrapper_70_io_in = ~ x315; // @[package.scala 94:16:@34493.4]
  assign RetimeWrapper_71_clock = clock; // @[:@34503.4]
  assign RetimeWrapper_71_reset = reset; // @[:@34504.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34506.4]
  assign RetimeWrapper_71_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34505.4]
  assign x325_x7_1_clock = clock; // @[:@34551.4]
  assign x325_x7_1_reset = reset; // @[:@34552.4]
  assign x325_x7_1_io_a = x241_lb_0_io_rPort_7_output_0; // @[Math.scala 151:17:@34553.4]
  assign x325_x7_1_io_b = _T_1752[31:0]; // @[Math.scala 152:17:@34554.4]
  assign x325_x7_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34555.4]
  assign x326_x8_1_clock = clock; // @[:@34561.4]
  assign x326_x8_1_reset = reset; // @[:@34562.4]
  assign x326_x8_1_io_a = x241_lb_0_io_rPort_0_output_0; // @[Math.scala 151:17:@34563.4]
  assign x326_x8_1_io_b = _T_1755[31:0]; // @[Math.scala 152:17:@34564.4]
  assign x326_x8_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34565.4]
  assign x327_x7_1_clock = clock; // @[:@34571.4]
  assign x327_x7_1_reset = reset; // @[:@34572.4]
  assign x327_x7_1_io_a = _T_1758[31:0]; // @[Math.scala 151:17:@34573.4]
  assign x327_x7_1_io_b = _T_1761[31:0]; // @[Math.scala 152:17:@34574.4]
  assign x327_x7_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34575.4]
  assign x328_x8_1_clock = clock; // @[:@34581.4]
  assign x328_x8_1_reset = reset; // @[:@34582.4]
  assign x328_x8_1_io_a = x241_lb_0_io_rPort_1_output_0; // @[Math.scala 151:17:@34583.4]
  assign x328_x8_1_io_b = _T_1766[31:0]; // @[Math.scala 152:17:@34584.4]
  assign x328_x8_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34585.4]
  assign x329_x7_1_clock = clock; // @[:@34591.4]
  assign x329_x7_1_reset = reset; // @[:@34592.4]
  assign x329_x7_1_io_a = x325_x7_1_io_result; // @[Math.scala 151:17:@34593.4]
  assign x329_x7_1_io_b = x326_x8_1_io_result; // @[Math.scala 152:17:@34594.4]
  assign x329_x7_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34595.4]
  assign x330_x8_1_clock = clock; // @[:@34601.4]
  assign x330_x8_1_reset = reset; // @[:@34602.4]
  assign x330_x8_1_io_a = x327_x7_1_io_result; // @[Math.scala 151:17:@34603.4]
  assign x330_x8_1_io_b = x328_x8_1_io_result; // @[Math.scala 152:17:@34604.4]
  assign x330_x8_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34605.4]
  assign x331_x7_1_clock = clock; // @[:@34611.4]
  assign x331_x7_1_reset = reset; // @[:@34612.4]
  assign x331_x7_1_io_a = x329_x7_1_io_result; // @[Math.scala 151:17:@34613.4]
  assign x331_x7_1_io_b = x330_x8_1_io_result; // @[Math.scala 152:17:@34614.4]
  assign x331_x7_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34615.4]
  assign RetimeWrapper_72_clock = clock; // @[:@34621.4]
  assign RetimeWrapper_72_reset = reset; // @[:@34622.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34624.4]
  assign RetimeWrapper_72_io_in = x241_lb_0_io_rPort_5_output_0; // @[package.scala 94:16:@34623.4]
  assign x332_sum_1_clock = clock; // @[:@34630.4]
  assign x332_sum_1_reset = reset; // @[:@34631.4]
  assign x332_sum_1_io_a = x331_x7_1_io_result; // @[Math.scala 151:17:@34632.4]
  assign x332_sum_1_io_b = RetimeWrapper_72_io_out; // @[Math.scala 152:17:@34633.4]
  assign x332_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@34634.4]
  assign x333_1_io_b = x332_sum_1_io_result; // @[Math.scala 721:17:@34642.4]
  assign x334_mul_1_clock = clock; // @[:@34651.4]
  assign x334_mul_1_io_a = x333_1_io_result; // @[Math.scala 263:17:@34653.4]
  assign x334_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@34654.4]
  assign x334_mul_1_io_flow = io_in_x210_TREADY; // @[Math.scala 265:20:@34655.4]
  assign x335_1_io_b = x334_mul_1_io_result; // @[Math.scala 721:17:@34663.4]
  assign RetimeWrapper_73_clock = clock; // @[:@34670.4]
  assign RetimeWrapper_73_reset = reset; // @[:@34671.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34673.4]
  assign RetimeWrapper_73_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@34672.4]
  assign RetimeWrapper_74_clock = clock; // @[:@34679.4]
  assign RetimeWrapper_74_reset = reset; // @[:@34680.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34682.4]
  assign RetimeWrapper_74_io_in = x499_x432_D1 ? x501_x431_sum_D1_number : x434_sub_number; // @[package.scala 94:16:@34681.4]
  assign RetimeWrapper_75_clock = clock; // @[:@34688.4]
  assign RetimeWrapper_75_reset = reset; // @[:@34689.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34691.4]
  assign RetimeWrapper_75_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@34690.4]
  assign RetimeWrapper_76_clock = clock; // @[:@34697.4]
  assign RetimeWrapper_76_reset = reset; // @[:@34698.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34700.4]
  assign RetimeWrapper_76_io_in = $unsigned(_T_258); // @[package.scala 94:16:@34699.4]
  assign RetimeWrapper_77_clock = clock; // @[:@34706.4]
  assign RetimeWrapper_77_reset = reset; // @[:@34707.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34709.4]
  assign RetimeWrapper_77_io_in = x335_1_io_result; // @[package.scala 94:16:@34708.4]
  assign RetimeWrapper_78_clock = clock; // @[:@34715.4]
  assign RetimeWrapper_78_reset = reset; // @[:@34716.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34718.4]
  assign RetimeWrapper_78_io_in = x251_sum_1_io_result; // @[package.scala 94:16:@34717.4]
  assign RetimeWrapper_79_clock = clock; // @[:@34726.4]
  assign RetimeWrapper_79_reset = reset; // @[:@34727.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34729.4]
  assign RetimeWrapper_79_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34728.4]
  assign RetimeWrapper_80_clock = clock; // @[:@34747.4]
  assign RetimeWrapper_80_reset = reset; // @[:@34748.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34750.4]
  assign RetimeWrapper_80_io_in = ~ x256; // @[package.scala 94:16:@34749.4]
  assign RetimeWrapper_81_clock = clock; // @[:@34756.4]
  assign RetimeWrapper_81_reset = reset; // @[:@34757.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34759.4]
  assign RetimeWrapper_81_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@34758.4]
  assign RetimeWrapper_82_clock = clock; // @[:@34765.4]
  assign RetimeWrapper_82_reset = reset; // @[:@34766.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34768.4]
  assign RetimeWrapper_82_io_in = x499_x432_D1 ? x501_x431_sum_D1_number : x434_sub_number; // @[package.scala 94:16:@34767.4]
  assign RetimeWrapper_83_clock = clock; // @[:@34774.4]
  assign RetimeWrapper_83_reset = reset; // @[:@34775.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34777.4]
  assign RetimeWrapper_83_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@34776.4]
  assign RetimeWrapper_84_clock = clock; // @[:@34783.4]
  assign RetimeWrapper_84_reset = reset; // @[:@34784.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34786.4]
  assign RetimeWrapper_84_io_in = $unsigned(_T_258); // @[package.scala 94:16:@34785.4]
  assign RetimeWrapper_85_clock = clock; // @[:@34792.4]
  assign RetimeWrapper_85_reset = reset; // @[:@34793.4]
  assign RetimeWrapper_85_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34795.4]
  assign RetimeWrapper_85_io_in = x251_sum_1_io_result; // @[package.scala 94:16:@34794.4]
  assign RetimeWrapper_86_clock = clock; // @[:@34804.4]
  assign RetimeWrapper_86_reset = reset; // @[:@34805.4]
  assign RetimeWrapper_86_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34807.4]
  assign RetimeWrapper_86_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34806.4]
  assign RetimeWrapper_87_clock = clock; // @[:@34825.4]
  assign RetimeWrapper_87_reset = reset; // @[:@34826.4]
  assign RetimeWrapper_87_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34828.4]
  assign RetimeWrapper_87_io_in = x457 ? x517_x456_sum_D1_number : x459_sub_number; // @[package.scala 94:16:@34827.4]
  assign RetimeWrapper_88_clock = clock; // @[:@34834.4]
  assign RetimeWrapper_88_reset = reset; // @[:@34835.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34837.4]
  assign RetimeWrapper_88_io_in = x266_sum_1_io_result; // @[package.scala 94:16:@34836.4]
  assign RetimeWrapper_89_clock = clock; // @[:@34843.4]
  assign RetimeWrapper_89_reset = reset; // @[:@34844.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34846.4]
  assign RetimeWrapper_89_io_in = ~ x262; // @[package.scala 94:16:@34845.4]
  assign RetimeWrapper_90_clock = clock; // @[:@34855.4]
  assign RetimeWrapper_90_reset = reset; // @[:@34856.4]
  assign RetimeWrapper_90_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34858.4]
  assign RetimeWrapper_90_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34857.4]
  assign RetimeWrapper_91_clock = clock; // @[:@34876.4]
  assign RetimeWrapper_91_reset = reset; // @[:@34877.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34879.4]
  assign RetimeWrapper_91_io_in = $unsigned(_T_1430); // @[package.scala 94:16:@34878.4]
  assign RetimeWrapper_92_clock = clock; // @[:@34885.4]
  assign RetimeWrapper_92_reset = reset; // @[:@34886.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34888.4]
  assign RetimeWrapper_92_io_in = x286_sum_1_io_result; // @[package.scala 94:16:@34887.4]
  assign RetimeWrapper_93_clock = clock; // @[:@34894.4]
  assign RetimeWrapper_93_reset = reset; // @[:@34895.4]
  assign RetimeWrapper_93_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34897.4]
  assign RetimeWrapper_93_io_in = ~ x281; // @[package.scala 94:16:@34896.4]
  assign RetimeWrapper_94_clock = clock; // @[:@34906.4]
  assign RetimeWrapper_94_reset = reset; // @[:@34907.4]
  assign RetimeWrapper_94_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34909.4]
  assign RetimeWrapper_94_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34908.4]
  assign RetimeWrapper_95_clock = clock; // @[:@34927.4]
  assign RetimeWrapper_95_reset = reset; // @[:@34928.4]
  assign RetimeWrapper_95_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34930.4]
  assign RetimeWrapper_95_io_in = x291_sum_1_io_result; // @[package.scala 94:16:@34929.4]
  assign RetimeWrapper_96_clock = clock; // @[:@34936.4]
  assign RetimeWrapper_96_reset = reset; // @[:@34937.4]
  assign RetimeWrapper_96_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34939.4]
  assign RetimeWrapper_96_io_in = ~ x289; // @[package.scala 94:16:@34938.4]
  assign RetimeWrapper_97_clock = clock; // @[:@34948.4]
  assign RetimeWrapper_97_reset = reset; // @[:@34949.4]
  assign RetimeWrapper_97_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34951.4]
  assign RetimeWrapper_97_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34950.4]
  assign RetimeWrapper_98_clock = clock; // @[:@34971.4]
  assign RetimeWrapper_98_reset = reset; // @[:@34972.4]
  assign RetimeWrapper_98_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@34974.4]
  assign RetimeWrapper_98_io_in = _GEN_11 << 1; // @[package.scala 94:16:@34973.4]
  assign RetimeWrapper_99_clock = clock; // @[:@34983.4]
  assign RetimeWrapper_99_reset = reset; // @[:@34984.4]
  assign RetimeWrapper_99_io_flow = io_in_x210_TREADY; // @[package.scala 95:18:@34986.4]
  assign RetimeWrapper_99_io_in = _GEN_12 << 2; // @[package.scala 94:16:@34985.4]
  assign RetimeWrapper_100_clock = clock; // @[:@34993.4]
  assign RetimeWrapper_100_reset = reset; // @[:@34994.4]
  assign RetimeWrapper_100_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34996.4]
  assign RetimeWrapper_100_io_in = x242_lb2_0_io_rPort_0_output_0; // @[package.scala 94:16:@34995.4]
  assign x349_x9_1_clock = clock; // @[:@35002.4]
  assign x349_x9_1_reset = reset; // @[:@35003.4]
  assign x349_x9_1_io_a = RetimeWrapper_100_io_out; // @[Math.scala 151:17:@35004.4]
  assign x349_x9_1_io_b = _T_1961[31:0]; // @[Math.scala 152:17:@35005.4]
  assign x349_x9_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@35006.4]
  assign RetimeWrapper_101_clock = clock; // @[:@35012.4]
  assign RetimeWrapper_101_reset = reset; // @[:@35013.4]
  assign RetimeWrapper_101_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35015.4]
  assign RetimeWrapper_101_io_in = x242_lb2_0_io_rPort_3_output_0; // @[package.scala 94:16:@35014.4]
  assign x350_x10_1_clock = clock; // @[:@35023.4]
  assign x350_x10_1_reset = reset; // @[:@35024.4]
  assign x350_x10_1_io_a = _T_1966[31:0]; // @[Math.scala 151:17:@35025.4]
  assign x350_x10_1_io_b = RetimeWrapper_101_io_out; // @[Math.scala 152:17:@35026.4]
  assign x350_x10_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@35027.4]
  assign x351_sum_1_clock = clock; // @[:@35033.4]
  assign x351_sum_1_reset = reset; // @[:@35034.4]
  assign x351_sum_1_io_a = x349_x9_1_io_result; // @[Math.scala 151:17:@35035.4]
  assign x351_sum_1_io_b = x350_x10_1_io_result; // @[Math.scala 152:17:@35036.4]
  assign x351_sum_1_io_flow = io_in_x210_TREADY; // @[Math.scala 153:20:@35037.4]
  assign x352_1_io_b = x351_sum_1_io_result; // @[Math.scala 721:17:@35045.4]
  assign x353_mul_1_clock = clock; // @[:@35054.4]
  assign x353_mul_1_io_a = x352_1_io_result; // @[Math.scala 263:17:@35056.4]
  assign x353_mul_1_io_b = 32'h10; // @[Math.scala 264:17:@35057.4]
  assign x353_mul_1_io_flow = io_in_x210_TREADY; // @[Math.scala 265:20:@35058.4]
  assign x354_1_io_b = x353_mul_1_io_result; // @[Math.scala 721:17:@35066.4]
  assign RetimeWrapper_102_clock = clock; // @[:@35077.4]
  assign RetimeWrapper_102_reset = reset; // @[:@35078.4]
  assign RetimeWrapper_102_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35080.4]
  assign RetimeWrapper_102_io_in = x354_1_io_result; // @[package.scala 94:16:@35079.4]
  assign RetimeWrapper_103_clock = clock; // @[:@35086.4]
  assign RetimeWrapper_103_reset = reset; // @[:@35087.4]
  assign RetimeWrapper_103_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35089.4]
  assign RetimeWrapper_103_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@35088.4]
  assign RetimeWrapper_104_clock = clock; // @[:@35095.4]
  assign RetimeWrapper_104_reset = reset; // @[:@35096.4]
  assign RetimeWrapper_104_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35098.4]
  assign RetimeWrapper_104_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@35097.4]
  assign RetimeWrapper_105_clock = clock; // @[:@35104.4]
  assign RetimeWrapper_105_reset = reset; // @[:@35105.4]
  assign RetimeWrapper_105_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35107.4]
  assign RetimeWrapper_105_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35106.4]
endmodule
module x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1( // @[:@35125.2]
  input          clock, // @[:@35126.4]
  input          reset, // @[:@35127.4]
  input          io_in_x209_TVALID, // @[:@35128.4]
  output         io_in_x209_TREADY, // @[:@35128.4]
  input  [255:0] io_in_x209_TDATA, // @[:@35128.4]
  input  [7:0]   io_in_x209_TID, // @[:@35128.4]
  input  [7:0]   io_in_x209_TDEST, // @[:@35128.4]
  output         io_in_x210_TVALID, // @[:@35128.4]
  input          io_in_x210_TREADY, // @[:@35128.4]
  output [255:0] io_in_x210_TDATA, // @[:@35128.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@35128.4]
  input          io_sigsIn_smChildAcks_0, // @[:@35128.4]
  output         io_sigsOut_smDoneIn_0, // @[:@35128.4]
  input          io_rr // @[:@35128.4]
);
  wire  x234_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@35162.4]
  wire  x234_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@35162.4]
  wire  x234_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@35162.4]
  wire  x234_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@35162.4]
  wire [12:0] x234_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@35162.4]
  wire [12:0] x234_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@35162.4]
  wire  x234_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@35162.4]
  wire  x234_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@35162.4]
  wire  x234_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@35162.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 32:18:@35222.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 32:18:@35222.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 32:18:@35222.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 32:18:@35222.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 32:18:@35222.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 32:18:@35222.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 32:18:@35222.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 32:18:@35222.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 32:18:@35222.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 32:18:@35222.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 32:18:@35222.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 32:18:@35222.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@35250.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@35250.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@35250.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@35250.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@35250.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@35292.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@35292.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@35292.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@35292.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@35292.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@35300.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@35300.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@35300.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@35300.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@35300.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x209_TREADY; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire [255:0] x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x209_TDATA; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire [7:0] x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x209_TID; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire [7:0] x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x209_TDEST; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x210_TVALID; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x210_TREADY; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire [255:0] x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x210_TDATA; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire [31:0] x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire [31:0] x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
  wire  _T_240; // @[package.scala 96:25:@35255.4 package.scala 96:25:@35256.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x360_outr_UnitPipe.scala 69:66:@35261.4]
  wire  _T_253; // @[package.scala 96:25:@35297.4 package.scala 96:25:@35298.4]
  wire  _T_259; // @[package.scala 96:25:@35305.4 package.scala 96:25:@35306.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@35308.4]
  wire  x359_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@35309.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@35317.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@35318.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@35330.4]
  x217_ctrchain x234_ctrchain ( // @[SpatialBlocks.scala 37:22:@35162.4]
    .clock(x234_ctrchain_clock),
    .reset(x234_ctrchain_reset),
    .io_input_reset(x234_ctrchain_io_input_reset),
    .io_input_enable(x234_ctrchain_io_input_enable),
    .io_output_counts_1(x234_ctrchain_io_output_counts_1),
    .io_output_counts_0(x234_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x234_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x234_ctrchain_io_output_oobs_1),
    .io_output_done(x234_ctrchain_io_output_done)
  );
  x359_inr_Foreach_SAMPLER_BOX_sm x359_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 32:18:@35222.4]
    .clock(x359_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x359_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x359_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x359_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x359_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x359_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x359_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x359_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x359_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x359_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x359_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x359_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@35250.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@35292.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@35300.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1 x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 672:24:@35334.4]
    .clock(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x209_TREADY(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x209_TREADY),
    .io_in_x209_TDATA(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x209_TDATA),
    .io_in_x209_TID(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x209_TID),
    .io_in_x209_TDEST(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x209_TDEST),
    .io_in_x210_TVALID(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x210_TVALID),
    .io_in_x210_TREADY(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x210_TREADY),
    .io_in_x210_TDATA(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x210_TDATA),
    .io_sigsIn_backpressure(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@35255.4 package.scala 96:25:@35256.4]
  assign x359_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x209_TVALID | x359_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x360_outr_UnitPipe.scala 69:66:@35261.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@35297.4 package.scala 96:25:@35298.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@35305.4 package.scala 96:25:@35306.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@35308.4]
  assign x359_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@35309.4]
  assign _T_264 = x359_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@35317.4]
  assign _T_265 = ~ x359_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@35318.4]
  assign _T_272 = x359_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@35330.4]
  assign io_in_x209_TREADY = x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x209_TREADY; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 48:23:@35392.4]
  assign io_in_x210_TVALID = x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x210_TVALID; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 49:23:@35402.4]
  assign io_in_x210_TDATA = x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x210_TDATA; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 49:23:@35400.4]
  assign io_sigsOut_smDoneIn_0 = x359_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@35315.4]
  assign x234_ctrchain_clock = clock; // @[:@35163.4]
  assign x234_ctrchain_reset = reset; // @[:@35164.4]
  assign x234_ctrchain_io_input_reset = x359_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@35333.4]
  assign x234_ctrchain_io_input_enable = _T_272 & x359_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@35285.4 SpatialBlocks.scala 159:42:@35332.4]
  assign x359_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@35223.4]
  assign x359_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@35224.4]
  assign x359_inr_Foreach_SAMPLER_BOX_sm_io_enable = x359_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x359_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@35312.4]
  assign x359_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x360_outr_UnitPipe.scala 67:50:@35258.4]
  assign x359_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@35314.4]
  assign x359_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x210_TREADY | x359_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@35286.4]
  assign x359_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x360_outr_UnitPipe.scala 71:48:@35264.4]
  assign RetimeWrapper_clock = clock; // @[:@35251.4]
  assign RetimeWrapper_reset = reset; // @[:@35252.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@35254.4]
  assign RetimeWrapper_io_in = x234_ctrchain_io_output_done; // @[package.scala 94:16:@35253.4]
  assign RetimeWrapper_1_clock = clock; // @[:@35293.4]
  assign RetimeWrapper_1_reset = reset; // @[:@35294.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@35296.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@35295.4]
  assign RetimeWrapper_2_clock = clock; // @[:@35301.4]
  assign RetimeWrapper_2_reset = reset; // @[:@35302.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@35304.4]
  assign RetimeWrapper_2_io_in = x359_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@35303.4]
  assign x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@35335.4]
  assign x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@35336.4]
  assign x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x209_TDATA = io_in_x209_TDATA; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 48:23:@35391.4]
  assign x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x209_TID = io_in_x209_TID; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 48:23:@35387.4]
  assign x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x209_TDEST = io_in_x209_TDEST; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 48:23:@35386.4]
  assign x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x210_TREADY = io_in_x210_TREADY; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 49:23:@35401.4]
  assign x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x210_TREADY | x359_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 677:22:@35419.4]
  assign x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 677:22:@35417.4]
  assign x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x359_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 677:22:@35415.4]
  assign x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x234_ctrchain_io_output_counts_1[12]}},x234_ctrchain_io_output_counts_1}; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 677:22:@35410.4]
  assign x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x234_ctrchain_io_output_counts_0[12]}},x234_ctrchain_io_output_counts_0}; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 677:22:@35409.4]
  assign x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x234_ctrchain_io_output_oobs_0; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 677:22:@35407.4]
  assign x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x234_ctrchain_io_output_oobs_1; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 677:22:@35408.4]
  assign x359_inr_Foreach_SAMPLER_BOX_kernelx359_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x359_inr_Foreach_SAMPLER_BOX.scala 676:18:@35403.4]
endmodule
module x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1( // @[:@35433.2]
  input          clock, // @[:@35434.4]
  input          reset, // @[:@35435.4]
  input          io_in_x209_TVALID, // @[:@35436.4]
  output         io_in_x209_TREADY, // @[:@35436.4]
  input  [255:0] io_in_x209_TDATA, // @[:@35436.4]
  input  [7:0]   io_in_x209_TID, // @[:@35436.4]
  input  [7:0]   io_in_x209_TDEST, // @[:@35436.4]
  output         io_in_x210_TVALID, // @[:@35436.4]
  input          io_in_x210_TREADY, // @[:@35436.4]
  output [255:0] io_in_x210_TDATA, // @[:@35436.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@35436.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@35436.4]
  input          io_sigsIn_smChildAcks_0, // @[:@35436.4]
  input          io_sigsIn_smChildAcks_1, // @[:@35436.4]
  output         io_sigsOut_smDoneIn_0, // @[:@35436.4]
  output         io_sigsOut_smDoneIn_1, // @[:@35436.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@35436.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@35436.4]
  input          io_rr // @[:@35436.4]
);
  wire  x212_fifoinraw_0_clock; // @[m_x212_fifoinraw_0.scala 27:17:@35450.4]
  wire  x212_fifoinraw_0_reset; // @[m_x212_fifoinraw_0.scala 27:17:@35450.4]
  wire  x213_fifoinpacked_0_clock; // @[m_x213_fifoinpacked_0.scala 27:17:@35474.4]
  wire  x213_fifoinpacked_0_reset; // @[m_x213_fifoinpacked_0.scala 27:17:@35474.4]
  wire  x213_fifoinpacked_0_io_wPort_0_en_0; // @[m_x213_fifoinpacked_0.scala 27:17:@35474.4]
  wire  x213_fifoinpacked_0_io_full; // @[m_x213_fifoinpacked_0.scala 27:17:@35474.4]
  wire  x213_fifoinpacked_0_io_active_0_in; // @[m_x213_fifoinpacked_0.scala 27:17:@35474.4]
  wire  x213_fifoinpacked_0_io_active_0_out; // @[m_x213_fifoinpacked_0.scala 27:17:@35474.4]
  wire  x214_fifooutraw_0_clock; // @[m_x214_fifooutraw_0.scala 27:17:@35498.4]
  wire  x214_fifooutraw_0_reset; // @[m_x214_fifooutraw_0.scala 27:17:@35498.4]
  wire  x217_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@35522.4]
  wire  x217_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@35522.4]
  wire  x217_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@35522.4]
  wire  x217_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@35522.4]
  wire [12:0] x217_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@35522.4]
  wire [12:0] x217_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@35522.4]
  wire  x217_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@35522.4]
  wire  x217_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@35522.4]
  wire  x217_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@35522.4]
  wire  x230_inr_Foreach_sm_clock; // @[sm_x230_inr_Foreach.scala 32:18:@35582.4]
  wire  x230_inr_Foreach_sm_reset; // @[sm_x230_inr_Foreach.scala 32:18:@35582.4]
  wire  x230_inr_Foreach_sm_io_enable; // @[sm_x230_inr_Foreach.scala 32:18:@35582.4]
  wire  x230_inr_Foreach_sm_io_done; // @[sm_x230_inr_Foreach.scala 32:18:@35582.4]
  wire  x230_inr_Foreach_sm_io_doneLatch; // @[sm_x230_inr_Foreach.scala 32:18:@35582.4]
  wire  x230_inr_Foreach_sm_io_ctrDone; // @[sm_x230_inr_Foreach.scala 32:18:@35582.4]
  wire  x230_inr_Foreach_sm_io_datapathEn; // @[sm_x230_inr_Foreach.scala 32:18:@35582.4]
  wire  x230_inr_Foreach_sm_io_ctrInc; // @[sm_x230_inr_Foreach.scala 32:18:@35582.4]
  wire  x230_inr_Foreach_sm_io_ctrRst; // @[sm_x230_inr_Foreach.scala 32:18:@35582.4]
  wire  x230_inr_Foreach_sm_io_parentAck; // @[sm_x230_inr_Foreach.scala 32:18:@35582.4]
  wire  x230_inr_Foreach_sm_io_backpressure; // @[sm_x230_inr_Foreach.scala 32:18:@35582.4]
  wire  x230_inr_Foreach_sm_io_break; // @[sm_x230_inr_Foreach.scala 32:18:@35582.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@35610.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@35610.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@35610.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@35610.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@35610.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@35656.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@35656.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@35656.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@35656.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@35656.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@35664.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@35664.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@35664.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@35664.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@35664.4]
  wire  x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_clock; // @[sm_x230_inr_Foreach.scala 92:24:@35699.4]
  wire  x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_reset; // @[sm_x230_inr_Foreach.scala 92:24:@35699.4]
  wire  x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_in_x213_fifoinpacked_0_wPort_0_en_0; // @[sm_x230_inr_Foreach.scala 92:24:@35699.4]
  wire  x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_in_x213_fifoinpacked_0_full; // @[sm_x230_inr_Foreach.scala 92:24:@35699.4]
  wire  x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_in_x213_fifoinpacked_0_active_0_in; // @[sm_x230_inr_Foreach.scala 92:24:@35699.4]
  wire  x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_in_x213_fifoinpacked_0_active_0_out; // @[sm_x230_inr_Foreach.scala 92:24:@35699.4]
  wire  x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x230_inr_Foreach.scala 92:24:@35699.4]
  wire  x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x230_inr_Foreach.scala 92:24:@35699.4]
  wire  x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x230_inr_Foreach.scala 92:24:@35699.4]
  wire [31:0] x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x230_inr_Foreach.scala 92:24:@35699.4]
  wire [31:0] x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x230_inr_Foreach.scala 92:24:@35699.4]
  wire  x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x230_inr_Foreach.scala 92:24:@35699.4]
  wire  x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x230_inr_Foreach.scala 92:24:@35699.4]
  wire  x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_rr; // @[sm_x230_inr_Foreach.scala 92:24:@35699.4]
  wire  x360_outr_UnitPipe_sm_clock; // @[sm_x360_outr_UnitPipe.scala 32:18:@35831.4]
  wire  x360_outr_UnitPipe_sm_reset; // @[sm_x360_outr_UnitPipe.scala 32:18:@35831.4]
  wire  x360_outr_UnitPipe_sm_io_enable; // @[sm_x360_outr_UnitPipe.scala 32:18:@35831.4]
  wire  x360_outr_UnitPipe_sm_io_done; // @[sm_x360_outr_UnitPipe.scala 32:18:@35831.4]
  wire  x360_outr_UnitPipe_sm_io_rst; // @[sm_x360_outr_UnitPipe.scala 32:18:@35831.4]
  wire  x360_outr_UnitPipe_sm_io_ctrDone; // @[sm_x360_outr_UnitPipe.scala 32:18:@35831.4]
  wire  x360_outr_UnitPipe_sm_io_ctrInc; // @[sm_x360_outr_UnitPipe.scala 32:18:@35831.4]
  wire  x360_outr_UnitPipe_sm_io_parentAck; // @[sm_x360_outr_UnitPipe.scala 32:18:@35831.4]
  wire  x360_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x360_outr_UnitPipe.scala 32:18:@35831.4]
  wire  x360_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x360_outr_UnitPipe.scala 32:18:@35831.4]
  wire  x360_outr_UnitPipe_sm_io_childAck_0; // @[sm_x360_outr_UnitPipe.scala 32:18:@35831.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@35888.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@35888.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@35888.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@35888.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@35888.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@35896.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@35896.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@35896.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@35896.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@35896.4]
  wire  x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_clock; // @[sm_x360_outr_UnitPipe.scala 76:24:@35926.4]
  wire  x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_reset; // @[sm_x360_outr_UnitPipe.scala 76:24:@35926.4]
  wire  x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x209_TVALID; // @[sm_x360_outr_UnitPipe.scala 76:24:@35926.4]
  wire  x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x209_TREADY; // @[sm_x360_outr_UnitPipe.scala 76:24:@35926.4]
  wire [255:0] x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x209_TDATA; // @[sm_x360_outr_UnitPipe.scala 76:24:@35926.4]
  wire [7:0] x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x209_TID; // @[sm_x360_outr_UnitPipe.scala 76:24:@35926.4]
  wire [7:0] x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x209_TDEST; // @[sm_x360_outr_UnitPipe.scala 76:24:@35926.4]
  wire  x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x210_TVALID; // @[sm_x360_outr_UnitPipe.scala 76:24:@35926.4]
  wire  x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x210_TREADY; // @[sm_x360_outr_UnitPipe.scala 76:24:@35926.4]
  wire [255:0] x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x210_TDATA; // @[sm_x360_outr_UnitPipe.scala 76:24:@35926.4]
  wire  x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x360_outr_UnitPipe.scala 76:24:@35926.4]
  wire  x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x360_outr_UnitPipe.scala 76:24:@35926.4]
  wire  x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x360_outr_UnitPipe.scala 76:24:@35926.4]
  wire  x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_rr; // @[sm_x360_outr_UnitPipe.scala 76:24:@35926.4]
  wire  _T_254; // @[package.scala 96:25:@35615.4 package.scala 96:25:@35616.4]
  wire  _T_260; // @[implicits.scala 47:10:@35619.4]
  wire  _T_261; // @[sm_x361_outr_UnitPipe.scala 70:41:@35620.4]
  wire  _T_262; // @[sm_x361_outr_UnitPipe.scala 70:78:@35621.4]
  wire  _T_263; // @[sm_x361_outr_UnitPipe.scala 70:76:@35622.4]
  wire  _T_275; // @[package.scala 96:25:@35661.4 package.scala 96:25:@35662.4]
  wire  _T_281; // @[package.scala 96:25:@35669.4 package.scala 96:25:@35670.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@35672.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@35681.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@35682.4]
  wire  _T_354; // @[package.scala 100:49:@35859.4]
  reg  _T_357; // @[package.scala 48:56:@35860.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@35893.4 package.scala 96:25:@35894.4]
  wire  _T_377; // @[package.scala 96:25:@35901.4 package.scala 96:25:@35902.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@35904.4]
  x212_fifoinraw_0 x212_fifoinraw_0 ( // @[m_x212_fifoinraw_0.scala 27:17:@35450.4]
    .clock(x212_fifoinraw_0_clock),
    .reset(x212_fifoinraw_0_reset)
  );
  x213_fifoinpacked_0 x213_fifoinpacked_0 ( // @[m_x213_fifoinpacked_0.scala 27:17:@35474.4]
    .clock(x213_fifoinpacked_0_clock),
    .reset(x213_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x213_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x213_fifoinpacked_0_io_full),
    .io_active_0_in(x213_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x213_fifoinpacked_0_io_active_0_out)
  );
  x212_fifoinraw_0 x214_fifooutraw_0 ( // @[m_x214_fifooutraw_0.scala 27:17:@35498.4]
    .clock(x214_fifooutraw_0_clock),
    .reset(x214_fifooutraw_0_reset)
  );
  x217_ctrchain x217_ctrchain ( // @[SpatialBlocks.scala 37:22:@35522.4]
    .clock(x217_ctrchain_clock),
    .reset(x217_ctrchain_reset),
    .io_input_reset(x217_ctrchain_io_input_reset),
    .io_input_enable(x217_ctrchain_io_input_enable),
    .io_output_counts_1(x217_ctrchain_io_output_counts_1),
    .io_output_counts_0(x217_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x217_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x217_ctrchain_io_output_oobs_1),
    .io_output_done(x217_ctrchain_io_output_done)
  );
  x230_inr_Foreach_sm x230_inr_Foreach_sm ( // @[sm_x230_inr_Foreach.scala 32:18:@35582.4]
    .clock(x230_inr_Foreach_sm_clock),
    .reset(x230_inr_Foreach_sm_reset),
    .io_enable(x230_inr_Foreach_sm_io_enable),
    .io_done(x230_inr_Foreach_sm_io_done),
    .io_doneLatch(x230_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x230_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x230_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x230_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x230_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x230_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x230_inr_Foreach_sm_io_backpressure),
    .io_break(x230_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@35610.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@35656.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@35664.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x230_inr_Foreach_kernelx230_inr_Foreach_concrete1 x230_inr_Foreach_kernelx230_inr_Foreach_concrete1 ( // @[sm_x230_inr_Foreach.scala 92:24:@35699.4]
    .clock(x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_clock),
    .reset(x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_reset),
    .io_in_x213_fifoinpacked_0_wPort_0_en_0(x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_in_x213_fifoinpacked_0_wPort_0_en_0),
    .io_in_x213_fifoinpacked_0_full(x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_in_x213_fifoinpacked_0_full),
    .io_in_x213_fifoinpacked_0_active_0_in(x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_in_x213_fifoinpacked_0_active_0_in),
    .io_in_x213_fifoinpacked_0_active_0_out(x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_in_x213_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x360_outr_UnitPipe_sm ( // @[sm_x360_outr_UnitPipe.scala 32:18:@35831.4]
    .clock(x360_outr_UnitPipe_sm_clock),
    .reset(x360_outr_UnitPipe_sm_reset),
    .io_enable(x360_outr_UnitPipe_sm_io_enable),
    .io_done(x360_outr_UnitPipe_sm_io_done),
    .io_rst(x360_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x360_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x360_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x360_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x360_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x360_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x360_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@35888.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@35896.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1 x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1 ( // @[sm_x360_outr_UnitPipe.scala 76:24:@35926.4]
    .clock(x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_clock),
    .reset(x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_reset),
    .io_in_x209_TVALID(x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x209_TVALID),
    .io_in_x209_TREADY(x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x209_TREADY),
    .io_in_x209_TDATA(x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x209_TDATA),
    .io_in_x209_TID(x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x209_TID),
    .io_in_x209_TDEST(x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x209_TDEST),
    .io_in_x210_TVALID(x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x210_TVALID),
    .io_in_x210_TREADY(x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x210_TREADY),
    .io_in_x210_TDATA(x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x210_TDATA),
    .io_sigsIn_smEnableOuts_0(x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@35615.4 package.scala 96:25:@35616.4]
  assign _T_260 = x213_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@35619.4]
  assign _T_261 = ~ _T_260; // @[sm_x361_outr_UnitPipe.scala 70:41:@35620.4]
  assign _T_262 = ~ x213_fifoinpacked_0_io_active_0_out; // @[sm_x361_outr_UnitPipe.scala 70:78:@35621.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x361_outr_UnitPipe.scala 70:76:@35622.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@35661.4 package.scala 96:25:@35662.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@35669.4 package.scala 96:25:@35670.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@35672.4]
  assign _T_286 = x230_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@35681.4]
  assign _T_287 = ~ x230_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@35682.4]
  assign _T_354 = x360_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@35859.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@35893.4 package.scala 96:25:@35894.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@35901.4 package.scala 96:25:@35902.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@35904.4]
  assign io_in_x209_TREADY = x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x209_TREADY; // @[sm_x360_outr_UnitPipe.scala 48:23:@35982.4]
  assign io_in_x210_TVALID = x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x210_TVALID; // @[sm_x360_outr_UnitPipe.scala 49:23:@35992.4]
  assign io_in_x210_TDATA = x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x210_TDATA; // @[sm_x360_outr_UnitPipe.scala 49:23:@35990.4]
  assign io_sigsOut_smDoneIn_0 = x230_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@35679.4]
  assign io_sigsOut_smDoneIn_1 = x360_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@35911.4]
  assign io_sigsOut_smCtrCopyDone_0 = x230_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@35698.4]
  assign io_sigsOut_smCtrCopyDone_1 = x360_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@35925.4]
  assign x212_fifoinraw_0_clock = clock; // @[:@35451.4]
  assign x212_fifoinraw_0_reset = reset; // @[:@35452.4]
  assign x213_fifoinpacked_0_clock = clock; // @[:@35475.4]
  assign x213_fifoinpacked_0_reset = reset; // @[:@35476.4]
  assign x213_fifoinpacked_0_io_wPort_0_en_0 = x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_in_x213_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@35759.4]
  assign x213_fifoinpacked_0_io_active_0_in = x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_in_x213_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@35758.4]
  assign x214_fifooutraw_0_clock = clock; // @[:@35499.4]
  assign x214_fifooutraw_0_reset = reset; // @[:@35500.4]
  assign x217_ctrchain_clock = clock; // @[:@35523.4]
  assign x217_ctrchain_reset = reset; // @[:@35524.4]
  assign x217_ctrchain_io_input_reset = x230_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@35697.4]
  assign x217_ctrchain_io_input_enable = x230_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@35649.4 SpatialBlocks.scala 159:42:@35696.4]
  assign x230_inr_Foreach_sm_clock = clock; // @[:@35583.4]
  assign x230_inr_Foreach_sm_reset = reset; // @[:@35584.4]
  assign x230_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@35676.4]
  assign x230_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x361_outr_UnitPipe.scala 69:38:@35618.4]
  assign x230_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@35678.4]
  assign x230_inr_Foreach_sm_io_backpressure = _T_263 | x230_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@35650.4]
  assign x230_inr_Foreach_sm_io_break = 1'h0; // @[sm_x361_outr_UnitPipe.scala 73:36:@35628.4]
  assign RetimeWrapper_clock = clock; // @[:@35611.4]
  assign RetimeWrapper_reset = reset; // @[:@35612.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@35614.4]
  assign RetimeWrapper_io_in = x217_ctrchain_io_output_done; // @[package.scala 94:16:@35613.4]
  assign RetimeWrapper_1_clock = clock; // @[:@35657.4]
  assign RetimeWrapper_1_reset = reset; // @[:@35658.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@35660.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@35659.4]
  assign RetimeWrapper_2_clock = clock; // @[:@35665.4]
  assign RetimeWrapper_2_reset = reset; // @[:@35666.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@35668.4]
  assign RetimeWrapper_2_io_in = x230_inr_Foreach_sm_io_done; // @[package.scala 94:16:@35667.4]
  assign x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_clock = clock; // @[:@35700.4]
  assign x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_reset = reset; // @[:@35701.4]
  assign x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_in_x213_fifoinpacked_0_full = x213_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@35753.4]
  assign x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_in_x213_fifoinpacked_0_active_0_out = x213_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@35752.4]
  assign x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x230_inr_Foreach_sm_io_doneLatch; // @[sm_x230_inr_Foreach.scala 97:22:@35782.4]
  assign x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x230_inr_Foreach.scala 97:22:@35780.4]
  assign x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_break = x230_inr_Foreach_sm_io_break; // @[sm_x230_inr_Foreach.scala 97:22:@35778.4]
  assign x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x217_ctrchain_io_output_counts_1[12]}},x217_ctrchain_io_output_counts_1}; // @[sm_x230_inr_Foreach.scala 97:22:@35773.4]
  assign x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x217_ctrchain_io_output_counts_0[12]}},x217_ctrchain_io_output_counts_0}; // @[sm_x230_inr_Foreach.scala 97:22:@35772.4]
  assign x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x217_ctrchain_io_output_oobs_0; // @[sm_x230_inr_Foreach.scala 97:22:@35770.4]
  assign x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x217_ctrchain_io_output_oobs_1; // @[sm_x230_inr_Foreach.scala 97:22:@35771.4]
  assign x230_inr_Foreach_kernelx230_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x230_inr_Foreach.scala 96:18:@35766.4]
  assign x360_outr_UnitPipe_sm_clock = clock; // @[:@35832.4]
  assign x360_outr_UnitPipe_sm_reset = reset; // @[:@35833.4]
  assign x360_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@35908.4]
  assign x360_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@35883.4]
  assign x360_outr_UnitPipe_sm_io_ctrDone = x360_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x361_outr_UnitPipe.scala 78:40:@35863.4]
  assign x360_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@35910.4]
  assign x360_outr_UnitPipe_sm_io_doneIn_0 = x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@35880.4]
  assign RetimeWrapper_3_clock = clock; // @[:@35889.4]
  assign RetimeWrapper_3_reset = reset; // @[:@35890.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@35892.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@35891.4]
  assign RetimeWrapper_4_clock = clock; // @[:@35897.4]
  assign RetimeWrapper_4_reset = reset; // @[:@35898.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@35900.4]
  assign RetimeWrapper_4_io_in = x360_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@35899.4]
  assign x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_clock = clock; // @[:@35927.4]
  assign x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_reset = reset; // @[:@35928.4]
  assign x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x209_TVALID = io_in_x209_TVALID; // @[sm_x360_outr_UnitPipe.scala 48:23:@35983.4]
  assign x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x209_TDATA = io_in_x209_TDATA; // @[sm_x360_outr_UnitPipe.scala 48:23:@35981.4]
  assign x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x209_TID = io_in_x209_TID; // @[sm_x360_outr_UnitPipe.scala 48:23:@35977.4]
  assign x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x209_TDEST = io_in_x209_TDEST; // @[sm_x360_outr_UnitPipe.scala 48:23:@35976.4]
  assign x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_in_x210_TREADY = io_in_x210_TREADY; // @[sm_x360_outr_UnitPipe.scala 49:23:@35991.4]
  assign x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x360_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x360_outr_UnitPipe.scala 81:22:@36001.4]
  assign x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x360_outr_UnitPipe_sm_io_childAck_0; // @[sm_x360_outr_UnitPipe.scala 81:22:@35999.4]
  assign x360_outr_UnitPipe_kernelx360_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x360_outr_UnitPipe.scala 80:18:@35993.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x383_outr_UnitPipe_sm( // @[:@36490.2]
  input   clock, // @[:@36491.4]
  input   reset, // @[:@36492.4]
  input   io_enable, // @[:@36493.4]
  output  io_done, // @[:@36493.4]
  input   io_parentAck, // @[:@36493.4]
  input   io_doneIn_0, // @[:@36493.4]
  input   io_doneIn_1, // @[:@36493.4]
  input   io_doneIn_2, // @[:@36493.4]
  output  io_enableOut_0, // @[:@36493.4]
  output  io_enableOut_1, // @[:@36493.4]
  output  io_enableOut_2, // @[:@36493.4]
  output  io_childAck_0, // @[:@36493.4]
  output  io_childAck_1, // @[:@36493.4]
  output  io_childAck_2, // @[:@36493.4]
  input   io_ctrCopyDone_0, // @[:@36493.4]
  input   io_ctrCopyDone_1, // @[:@36493.4]
  input   io_ctrCopyDone_2 // @[:@36493.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@36496.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@36496.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@36496.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@36496.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@36496.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@36496.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@36499.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@36499.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@36499.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@36499.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@36499.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@36499.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@36502.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@36502.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@36502.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@36502.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@36502.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@36502.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@36505.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@36505.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@36505.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@36505.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@36505.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@36505.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@36508.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@36508.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@36508.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@36508.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@36508.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@36508.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@36511.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@36511.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@36511.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@36511.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@36511.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@36511.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@36552.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@36552.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@36552.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@36552.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@36552.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@36552.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@36555.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@36555.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@36555.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@36555.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@36555.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@36555.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@36558.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@36558.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@36558.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@36558.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@36558.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@36558.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@36609.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@36609.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@36609.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@36609.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@36609.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@36623.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@36623.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@36623.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@36623.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@36623.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@36641.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@36641.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@36641.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@36641.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@36641.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@36678.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@36678.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@36678.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@36678.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@36678.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@36692.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@36692.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@36692.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@36692.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@36692.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@36710.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@36710.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@36710.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@36710.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@36710.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@36747.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@36747.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@36747.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@36747.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@36747.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@36761.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@36761.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@36761.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@36761.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@36761.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@36779.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@36779.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@36779.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@36779.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@36779.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@36836.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@36836.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@36836.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@36836.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@36836.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@36853.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@36853.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@36853.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@36853.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@36853.4]
  wire  _T_77; // @[Controllers.scala 80:47:@36514.4]
  wire  allDone; // @[Controllers.scala 80:47:@36515.4]
  wire  _T_151; // @[Controllers.scala 165:35:@36593.4]
  wire  _T_153; // @[Controllers.scala 165:60:@36594.4]
  wire  _T_154; // @[Controllers.scala 165:58:@36595.4]
  wire  _T_156; // @[Controllers.scala 165:76:@36596.4]
  wire  _T_157; // @[Controllers.scala 165:74:@36597.4]
  wire  _T_161; // @[Controllers.scala 165:109:@36600.4]
  wire  _T_164; // @[Controllers.scala 165:141:@36602.4]
  wire  _T_172; // @[package.scala 96:25:@36614.4 package.scala 96:25:@36615.4]
  wire  _T_176; // @[Controllers.scala 167:54:@36617.4]
  wire  _T_177; // @[Controllers.scala 167:52:@36618.4]
  wire  _T_184; // @[package.scala 96:25:@36628.4 package.scala 96:25:@36629.4]
  wire  _T_202; // @[package.scala 96:25:@36646.4 package.scala 96:25:@36647.4]
  wire  _T_206; // @[Controllers.scala 169:67:@36649.4]
  wire  _T_207; // @[Controllers.scala 169:86:@36650.4]
  wire  _T_219; // @[Controllers.scala 165:35:@36662.4]
  wire  _T_221; // @[Controllers.scala 165:60:@36663.4]
  wire  _T_222; // @[Controllers.scala 165:58:@36664.4]
  wire  _T_224; // @[Controllers.scala 165:76:@36665.4]
  wire  _T_225; // @[Controllers.scala 165:74:@36666.4]
  wire  _T_229; // @[Controllers.scala 165:109:@36669.4]
  wire  _T_232; // @[Controllers.scala 165:141:@36671.4]
  wire  _T_240; // @[package.scala 96:25:@36683.4 package.scala 96:25:@36684.4]
  wire  _T_244; // @[Controllers.scala 167:54:@36686.4]
  wire  _T_245; // @[Controllers.scala 167:52:@36687.4]
  wire  _T_252; // @[package.scala 96:25:@36697.4 package.scala 96:25:@36698.4]
  wire  _T_270; // @[package.scala 96:25:@36715.4 package.scala 96:25:@36716.4]
  wire  _T_274; // @[Controllers.scala 169:67:@36718.4]
  wire  _T_275; // @[Controllers.scala 169:86:@36719.4]
  wire  _T_287; // @[Controllers.scala 165:35:@36731.4]
  wire  _T_289; // @[Controllers.scala 165:60:@36732.4]
  wire  _T_290; // @[Controllers.scala 165:58:@36733.4]
  wire  _T_292; // @[Controllers.scala 165:76:@36734.4]
  wire  _T_293; // @[Controllers.scala 165:74:@36735.4]
  wire  _T_297; // @[Controllers.scala 165:109:@36738.4]
  wire  _T_300; // @[Controllers.scala 165:141:@36740.4]
  wire  _T_308; // @[package.scala 96:25:@36752.4 package.scala 96:25:@36753.4]
  wire  _T_312; // @[Controllers.scala 167:54:@36755.4]
  wire  _T_313; // @[Controllers.scala 167:52:@36756.4]
  wire  _T_320; // @[package.scala 96:25:@36766.4 package.scala 96:25:@36767.4]
  wire  _T_338; // @[package.scala 96:25:@36784.4 package.scala 96:25:@36785.4]
  wire  _T_342; // @[Controllers.scala 169:67:@36787.4]
  wire  _T_343; // @[Controllers.scala 169:86:@36788.4]
  wire  _T_358; // @[Controllers.scala 213:68:@36806.4]
  wire  _T_360; // @[Controllers.scala 213:90:@36808.4]
  wire  _T_362; // @[Controllers.scala 213:132:@36810.4]
  wire  _T_366; // @[Controllers.scala 213:68:@36815.4]
  wire  _T_368; // @[Controllers.scala 213:90:@36817.4]
  wire  _T_374; // @[Controllers.scala 213:68:@36823.4]
  wire  _T_376; // @[Controllers.scala 213:90:@36825.4]
  wire  _T_383; // @[package.scala 100:49:@36831.4]
  reg  _T_386; // @[package.scala 48:56:@36832.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@36834.4]
  reg  _T_400; // @[package.scala 48:56:@36850.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@36496.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@36499.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@36502.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@36505.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@36508.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@36511.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@36552.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@36555.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@36558.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@36609.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@36623.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@36641.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@36678.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@36692.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@36710.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@36747.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@36761.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@36779.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@36836.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@36853.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@36514.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@36515.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@36593.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@36594.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@36595.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@36596.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@36597.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@36600.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@36602.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@36614.4 package.scala 96:25:@36615.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@36617.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@36618.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@36628.4 package.scala 96:25:@36629.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@36646.4 package.scala 96:25:@36647.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@36649.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@36650.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@36662.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@36663.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@36664.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@36665.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@36666.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@36669.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@36671.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@36683.4 package.scala 96:25:@36684.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@36686.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@36687.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@36697.4 package.scala 96:25:@36698.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@36715.4 package.scala 96:25:@36716.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@36718.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@36719.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@36731.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@36732.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@36733.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@36734.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@36735.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@36738.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@36740.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@36752.4 package.scala 96:25:@36753.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@36755.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@36756.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@36766.4 package.scala 96:25:@36767.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@36784.4 package.scala 96:25:@36785.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@36787.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@36788.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@36806.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@36808.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@36810.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@36815.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@36817.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@36823.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@36825.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@36831.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@36834.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@36860.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@36814.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@36822.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@36830.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@36801.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@36803.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@36805.4]
  assign active_0_clock = clock; // @[:@36497.4]
  assign active_0_reset = reset; // @[:@36498.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@36604.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@36608.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@36518.4]
  assign active_1_clock = clock; // @[:@36500.4]
  assign active_1_reset = reset; // @[:@36501.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@36673.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@36677.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@36519.4]
  assign active_2_clock = clock; // @[:@36503.4]
  assign active_2_reset = reset; // @[:@36504.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@36742.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@36746.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@36520.4]
  assign done_0_clock = clock; // @[:@36506.4]
  assign done_0_reset = reset; // @[:@36507.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@36654.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@36532.4 Controllers.scala 170:32:@36661.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@36521.4]
  assign done_1_clock = clock; // @[:@36509.4]
  assign done_1_reset = reset; // @[:@36510.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@36723.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@36541.4 Controllers.scala 170:32:@36730.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@36522.4]
  assign done_2_clock = clock; // @[:@36512.4]
  assign done_2_reset = reset; // @[:@36513.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@36792.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@36550.4 Controllers.scala 170:32:@36799.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@36523.4]
  assign iterDone_0_clock = clock; // @[:@36553.4]
  assign iterDone_0_reset = reset; // @[:@36554.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@36622.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@36572.4 Controllers.scala 168:36:@36638.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@36561.4]
  assign iterDone_1_clock = clock; // @[:@36556.4]
  assign iterDone_1_reset = reset; // @[:@36557.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@36691.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@36581.4 Controllers.scala 168:36:@36707.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@36562.4]
  assign iterDone_2_clock = clock; // @[:@36559.4]
  assign iterDone_2_reset = reset; // @[:@36560.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@36760.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@36590.4 Controllers.scala 168:36:@36776.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@36563.4]
  assign RetimeWrapper_clock = clock; // @[:@36610.4]
  assign RetimeWrapper_reset = reset; // @[:@36611.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@36613.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@36612.4]
  assign RetimeWrapper_1_clock = clock; // @[:@36624.4]
  assign RetimeWrapper_1_reset = reset; // @[:@36625.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@36627.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@36626.4]
  assign RetimeWrapper_2_clock = clock; // @[:@36642.4]
  assign RetimeWrapper_2_reset = reset; // @[:@36643.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@36645.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@36644.4]
  assign RetimeWrapper_3_clock = clock; // @[:@36679.4]
  assign RetimeWrapper_3_reset = reset; // @[:@36680.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@36682.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@36681.4]
  assign RetimeWrapper_4_clock = clock; // @[:@36693.4]
  assign RetimeWrapper_4_reset = reset; // @[:@36694.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@36696.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@36695.4]
  assign RetimeWrapper_5_clock = clock; // @[:@36711.4]
  assign RetimeWrapper_5_reset = reset; // @[:@36712.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@36714.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@36713.4]
  assign RetimeWrapper_6_clock = clock; // @[:@36748.4]
  assign RetimeWrapper_6_reset = reset; // @[:@36749.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@36751.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@36750.4]
  assign RetimeWrapper_7_clock = clock; // @[:@36762.4]
  assign RetimeWrapper_7_reset = reset; // @[:@36763.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@36765.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@36764.4]
  assign RetimeWrapper_8_clock = clock; // @[:@36780.4]
  assign RetimeWrapper_8_reset = reset; // @[:@36781.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@36783.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@36782.4]
  assign RetimeWrapper_9_clock = clock; // @[:@36837.4]
  assign RetimeWrapper_9_reset = reset; // @[:@36838.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@36840.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@36839.4]
  assign RetimeWrapper_10_clock = clock; // @[:@36854.4]
  assign RetimeWrapper_10_reset = reset; // @[:@36855.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@36857.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@36856.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x369_inr_UnitPipe_sm( // @[:@37033.2]
  input   clock, // @[:@37034.4]
  input   reset, // @[:@37035.4]
  input   io_enable, // @[:@37036.4]
  output  io_done, // @[:@37036.4]
  output  io_doneLatch, // @[:@37036.4]
  input   io_ctrDone, // @[:@37036.4]
  output  io_datapathEn, // @[:@37036.4]
  output  io_ctrInc, // @[:@37036.4]
  input   io_parentAck, // @[:@37036.4]
  input   io_backpressure // @[:@37036.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@37038.4]
  wire  active_reset; // @[Controllers.scala 261:22:@37038.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@37038.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@37038.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@37038.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@37038.4]
  wire  done_clock; // @[Controllers.scala 262:20:@37041.4]
  wire  done_reset; // @[Controllers.scala 262:20:@37041.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@37041.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@37041.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@37041.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@37041.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@37095.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@37095.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@37095.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@37095.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@37095.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@37103.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@37103.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@37103.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@37103.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@37103.4]
  wire  _T_80; // @[Controllers.scala 264:48:@37046.4]
  wire  _T_81; // @[Controllers.scala 264:46:@37047.4]
  wire  _T_82; // @[Controllers.scala 264:62:@37048.4]
  wire  _T_83; // @[Controllers.scala 264:60:@37049.4]
  wire  _T_100; // @[package.scala 100:49:@37066.4]
  reg  _T_103; // @[package.scala 48:56:@37067.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@37075.4]
  wire  _T_116; // @[Controllers.scala 283:41:@37083.4]
  wire  _T_117; // @[Controllers.scala 283:59:@37084.4]
  wire  _T_119; // @[Controllers.scala 284:37:@37087.4]
  reg  _T_125; // @[package.scala 48:56:@37091.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@37113.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@37116.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@37118.4]
  wire  _T_152; // @[Controllers.scala 292:61:@37119.4]
  wire  _T_153; // @[Controllers.scala 292:24:@37120.4]
  SRFF active ( // @[Controllers.scala 261:22:@37038.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@37041.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@37095.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@37103.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@37046.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@37047.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@37048.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@37049.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@37066.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@37075.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@37083.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@37084.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@37087.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@37118.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@37119.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@37120.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@37094.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@37122.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@37086.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@37089.4]
  assign active_clock = clock; // @[:@37039.4]
  assign active_reset = reset; // @[:@37040.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@37051.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@37055.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@37056.4]
  assign done_clock = clock; // @[:@37042.4]
  assign done_reset = reset; // @[:@37043.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@37071.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@37064.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@37065.4]
  assign RetimeWrapper_clock = clock; // @[:@37096.4]
  assign RetimeWrapper_reset = reset; // @[:@37097.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@37099.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@37098.4]
  assign RetimeWrapper_1_clock = clock; // @[:@37104.4]
  assign RetimeWrapper_1_reset = reset; // @[:@37105.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@37107.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@37106.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1( // @[:@37197.2]
  output        io_in_x362_valid, // @[:@37200.4]
  output [63:0] io_in_x362_bits_addr, // @[:@37200.4]
  output [31:0] io_in_x362_bits_size, // @[:@37200.4]
  input  [63:0] io_in_x207_outdram_number, // @[:@37200.4]
  input         io_sigsIn_backpressure, // @[:@37200.4]
  input         io_sigsIn_datapathEn, // @[:@37200.4]
  input         io_rr // @[:@37200.4]
);
  wire [96:0] x366_tuple; // @[Cat.scala 30:58:@37214.4]
  wire  _T_135; // @[implicits.scala 55:10:@37217.4]
  assign x366_tuple = {33'h7e9000,io_in_x207_outdram_number}; // @[Cat.scala 30:58:@37214.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@37217.4]
  assign io_in_x362_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x369_inr_UnitPipe.scala 65:18:@37220.4]
  assign io_in_x362_bits_addr = x366_tuple[63:0]; // @[sm_x369_inr_UnitPipe.scala 66:22:@37222.4]
  assign io_in_x362_bits_size = x366_tuple[95:64]; // @[sm_x369_inr_UnitPipe.scala 67:22:@37224.4]
endmodule
module FF_13( // @[:@37226.2]
  input         clock, // @[:@37227.4]
  input         reset, // @[:@37228.4]
  output [22:0] io_rPort_0_output_0, // @[:@37229.4]
  input  [22:0] io_wPort_0_data_0, // @[:@37229.4]
  input         io_wPort_0_reset, // @[:@37229.4]
  input         io_wPort_0_en_0 // @[:@37229.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 321:19:@37244.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 325:32:@37246.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 325:12:@37247.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@37246.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 325:12:@37247.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@37249.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@37264.2]
  input         clock, // @[:@37265.4]
  input         reset, // @[:@37266.4]
  input         io_input_reset, // @[:@37267.4]
  input         io_input_enable, // @[:@37267.4]
  output [22:0] io_output_count_0, // @[:@37267.4]
  output        io_output_oobs_0, // @[:@37267.4]
  output        io_output_done // @[:@37267.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@37280.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@37280.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@37280.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@37280.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@37280.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@37280.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@37296.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@37296.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@37296.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@37296.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@37296.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@37296.4]
  wire  _T_36; // @[Counter.scala 264:45:@37299.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@37324.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@37325.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@37326.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@37327.4]
  wire  _T_57; // @[Counter.scala 293:18:@37329.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@37337.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@37340.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@37341.4]
  wire  _T_75; // @[Counter.scala 322:102:@37345.4]
  wire  _T_77; // @[Counter.scala 322:130:@37346.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@37280.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@37296.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@37299.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@37324.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@37325.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@37326.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@37327.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@37329.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@37337.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@37340.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@37341.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@37345.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@37346.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@37344.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@37348.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@37350.4]
  assign bases_0_clock = clock; // @[:@37281.4]
  assign bases_0_reset = reset; // @[:@37282.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@37343.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@37322.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@37323.4]
  assign SRFF_clock = clock; // @[:@37297.4]
  assign SRFF_reset = reset; // @[:@37298.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@37301.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@37303.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@37304.4]
endmodule
module x371_ctrchain( // @[:@37355.2]
  input         clock, // @[:@37356.4]
  input         reset, // @[:@37357.4]
  input         io_input_reset, // @[:@37358.4]
  input         io_input_enable, // @[:@37358.4]
  output [22:0] io_output_counts_0, // @[:@37358.4]
  output        io_output_oobs_0, // @[:@37358.4]
  output        io_output_done // @[:@37358.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@37360.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@37360.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@37360.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@37360.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@37360.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@37360.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@37360.4]
  reg  wasDone; // @[Counter.scala 542:24:@37369.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@37375.4]
  wire  _T_47; // @[Counter.scala 546:80:@37376.4]
  reg  doneLatch; // @[Counter.scala 550:26:@37381.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@37382.4]
  wire  _T_55; // @[Counter.scala 551:19:@37383.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@37360.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@37375.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@37376.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@37382.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@37383.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@37385.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@37387.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@37378.4]
  assign ctrs_0_clock = clock; // @[:@37361.4]
  assign ctrs_0_reset = reset; // @[:@37362.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@37366.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@37367.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x378_inr_Foreach_sm( // @[:@37575.2]
  input   clock, // @[:@37576.4]
  input   reset, // @[:@37577.4]
  input   io_enable, // @[:@37578.4]
  output  io_done, // @[:@37578.4]
  output  io_doneLatch, // @[:@37578.4]
  input   io_ctrDone, // @[:@37578.4]
  output  io_datapathEn, // @[:@37578.4]
  output  io_ctrInc, // @[:@37578.4]
  output  io_ctrRst, // @[:@37578.4]
  input   io_parentAck, // @[:@37578.4]
  input   io_backpressure, // @[:@37578.4]
  input   io_break // @[:@37578.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@37580.4]
  wire  active_reset; // @[Controllers.scala 261:22:@37580.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@37580.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@37580.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@37580.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@37580.4]
  wire  done_clock; // @[Controllers.scala 262:20:@37583.4]
  wire  done_reset; // @[Controllers.scala 262:20:@37583.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@37583.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@37583.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@37583.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@37583.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@37617.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@37617.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@37617.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@37617.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@37617.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@37639.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@37639.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@37639.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@37639.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@37639.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@37651.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@37651.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@37651.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@37651.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@37651.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@37659.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@37659.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@37659.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@37659.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@37659.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@37675.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@37675.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@37675.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@37675.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@37675.4]
  wire  _T_80; // @[Controllers.scala 264:48:@37588.4]
  wire  _T_81; // @[Controllers.scala 264:46:@37589.4]
  wire  _T_82; // @[Controllers.scala 264:62:@37590.4]
  wire  _T_83; // @[Controllers.scala 264:60:@37591.4]
  wire  _T_100; // @[package.scala 100:49:@37608.4]
  reg  _T_103; // @[package.scala 48:56:@37609.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@37622.4 package.scala 96:25:@37623.4]
  wire  _T_110; // @[package.scala 100:49:@37624.4]
  reg  _T_113; // @[package.scala 48:56:@37625.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@37627.4]
  wire  _T_118; // @[Controllers.scala 283:41:@37632.4]
  wire  _T_119; // @[Controllers.scala 283:59:@37633.4]
  wire  _T_121; // @[Controllers.scala 284:37:@37636.4]
  wire  _T_124; // @[package.scala 96:25:@37644.4 package.scala 96:25:@37645.4]
  wire  _T_126; // @[package.scala 100:49:@37646.4]
  reg  _T_129; // @[package.scala 48:56:@37647.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@37669.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@37671.4]
  reg  _T_153; // @[package.scala 48:56:@37672.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@37680.4 package.scala 96:25:@37681.4]
  wire  _T_158; // @[Controllers.scala 292:61:@37682.4]
  wire  _T_159; // @[Controllers.scala 292:24:@37683.4]
  SRFF active ( // @[Controllers.scala 261:22:@37580.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@37583.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@37617.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@37639.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@37651.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@37659.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@37675.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@37588.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@37589.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@37590.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@37591.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@37608.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@37622.4 package.scala 96:25:@37623.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@37624.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@37627.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@37632.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@37633.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@37636.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@37644.4 package.scala 96:25:@37645.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@37646.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@37671.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@37680.4 package.scala 96:25:@37681.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@37682.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@37683.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@37650.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@37685.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@37635.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@37638.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@37630.4]
  assign active_clock = clock; // @[:@37581.4]
  assign active_reset = reset; // @[:@37582.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@37593.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@37597.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@37598.4]
  assign done_clock = clock; // @[:@37584.4]
  assign done_reset = reset; // @[:@37585.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@37613.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@37606.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@37607.4]
  assign RetimeWrapper_clock = clock; // @[:@37618.4]
  assign RetimeWrapper_reset = reset; // @[:@37619.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@37621.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@37620.4]
  assign RetimeWrapper_1_clock = clock; // @[:@37640.4]
  assign RetimeWrapper_1_reset = reset; // @[:@37641.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@37643.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@37642.4]
  assign RetimeWrapper_2_clock = clock; // @[:@37652.4]
  assign RetimeWrapper_2_reset = reset; // @[:@37653.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@37655.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@37654.4]
  assign RetimeWrapper_3_clock = clock; // @[:@37660.4]
  assign RetimeWrapper_3_reset = reset; // @[:@37661.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@37663.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@37662.4]
  assign RetimeWrapper_4_clock = clock; // @[:@37676.4]
  assign RetimeWrapper_4_reset = reset; // @[:@37677.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@37679.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@37678.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x378_inr_Foreach_kernelx378_inr_Foreach_concrete1( // @[:@37892.2]
  input         clock, // @[:@37893.4]
  input         reset, // @[:@37894.4]
  output [20:0] io_in_x211_outbuf_0_rPort_0_ofs_0, // @[:@37895.4]
  output        io_in_x211_outbuf_0_rPort_0_en_0, // @[:@37895.4]
  output        io_in_x211_outbuf_0_rPort_0_backpressure, // @[:@37895.4]
  input  [31:0] io_in_x211_outbuf_0_rPort_0_output_0, // @[:@37895.4]
  output        io_in_x363_valid, // @[:@37895.4]
  output [31:0] io_in_x363_bits_wdata_0, // @[:@37895.4]
  output        io_in_x363_bits_wstrb, // @[:@37895.4]
  input         io_sigsIn_backpressure, // @[:@37895.4]
  input         io_sigsIn_datapathEn, // @[:@37895.4]
  input         io_sigsIn_break, // @[:@37895.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@37895.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@37895.4]
  input         io_rr // @[:@37895.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@37922.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@37922.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@37951.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@37951.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@37951.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@37951.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@37951.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@37960.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@37960.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@37960.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@37960.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@37960.4]
  wire  b373; // @[sm_x378_inr_Foreach.scala 62:18:@37930.4]
  wire  _T_274; // @[sm_x378_inr_Foreach.scala 67:129:@37934.4]
  wire  _T_278; // @[implicits.scala 55:10:@37937.4]
  wire  _T_279; // @[sm_x378_inr_Foreach.scala 67:146:@37938.4]
  wire [32:0] x376_tuple; // @[Cat.scala 30:58:@37948.4]
  wire  _T_290; // @[package.scala 96:25:@37965.4 package.scala 96:25:@37966.4]
  wire  _T_292; // @[implicits.scala 55:10:@37967.4]
  wire  x565_b373_D2; // @[package.scala 96:25:@37956.4 package.scala 96:25:@37957.4]
  wire  _T_293; // @[sm_x378_inr_Foreach.scala 74:112:@37968.4]
  wire [31:0] b372_number; // @[Math.scala 723:22:@37927.4 Math.scala 724:14:@37928.4]
  _ _ ( // @[Math.scala 720:24:@37922.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@37951.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@37960.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b373 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x378_inr_Foreach.scala 62:18:@37930.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x378_inr_Foreach.scala 67:129:@37934.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@37937.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x378_inr_Foreach.scala 67:146:@37938.4]
  assign x376_tuple = {1'h1,io_in_x211_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@37948.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@37965.4 package.scala 96:25:@37966.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@37967.4]
  assign x565_b373_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@37956.4 package.scala 96:25:@37957.4]
  assign _T_293 = _T_292 & x565_b373_D2; // @[sm_x378_inr_Foreach.scala 74:112:@37968.4]
  assign b372_number = __io_result; // @[Math.scala 723:22:@37927.4 Math.scala 724:14:@37928.4]
  assign io_in_x211_outbuf_0_rPort_0_ofs_0 = b372_number[20:0]; // @[MemInterfaceType.scala 107:54:@37941.4]
  assign io_in_x211_outbuf_0_rPort_0_en_0 = _T_279 & b373; // @[MemInterfaceType.scala 110:79:@37943.4]
  assign io_in_x211_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@37942.4]
  assign io_in_x363_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x378_inr_Foreach.scala 74:18:@37970.4]
  assign io_in_x363_bits_wdata_0 = x376_tuple[31:0]; // @[sm_x378_inr_Foreach.scala 75:26:@37972.4]
  assign io_in_x363_bits_wstrb = x376_tuple[32]; // @[sm_x378_inr_Foreach.scala 76:23:@37974.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@37925.4]
  assign RetimeWrapper_clock = clock; // @[:@37952.4]
  assign RetimeWrapper_reset = reset; // @[:@37953.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37955.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@37954.4]
  assign RetimeWrapper_1_clock = clock; // @[:@37961.4]
  assign RetimeWrapper_1_reset = reset; // @[:@37962.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37964.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@37963.4]
endmodule
module x382_inr_UnitPipe_sm( // @[:@38130.2]
  input   clock, // @[:@38131.4]
  input   reset, // @[:@38132.4]
  input   io_enable, // @[:@38133.4]
  output  io_done, // @[:@38133.4]
  output  io_doneLatch, // @[:@38133.4]
  input   io_ctrDone, // @[:@38133.4]
  output  io_datapathEn, // @[:@38133.4]
  output  io_ctrInc, // @[:@38133.4]
  input   io_parentAck // @[:@38133.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@38135.4]
  wire  active_reset; // @[Controllers.scala 261:22:@38135.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@38135.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@38135.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@38135.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@38135.4]
  wire  done_clock; // @[Controllers.scala 262:20:@38138.4]
  wire  done_reset; // @[Controllers.scala 262:20:@38138.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@38138.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@38138.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@38138.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@38138.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@38172.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@38172.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@38172.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@38172.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@38172.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@38194.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@38194.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@38194.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@38194.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@38194.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@38206.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@38206.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@38206.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@38206.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@38206.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@38214.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@38214.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@38214.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@38214.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@38214.4]
  wire  _T_80; // @[Controllers.scala 264:48:@38143.4]
  wire  _T_81; // @[Controllers.scala 264:46:@38144.4]
  wire  _T_82; // @[Controllers.scala 264:62:@38145.4]
  wire  _T_100; // @[package.scala 100:49:@38163.4]
  reg  _T_103; // @[package.scala 48:56:@38164.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@38187.4]
  wire  _T_124; // @[package.scala 96:25:@38199.4 package.scala 96:25:@38200.4]
  wire  _T_126; // @[package.scala 100:49:@38201.4]
  reg  _T_129; // @[package.scala 48:56:@38202.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@38224.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@38226.4]
  reg  _T_153; // @[package.scala 48:56:@38227.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@38229.4]
  wire  _T_156; // @[Controllers.scala 292:61:@38230.4]
  wire  _T_157; // @[Controllers.scala 292:24:@38231.4]
  SRFF active ( // @[Controllers.scala 261:22:@38135.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@38138.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@38172.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@38194.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@38206.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@38214.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@38143.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@38144.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@38145.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@38163.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@38187.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@38199.4 package.scala 96:25:@38200.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@38201.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@38226.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@38229.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@38230.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@38231.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@38205.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@38233.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@38190.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@38193.4]
  assign active_clock = clock; // @[:@38136.4]
  assign active_reset = reset; // @[:@38137.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@38148.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@38152.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@38153.4]
  assign done_clock = clock; // @[:@38139.4]
  assign done_reset = reset; // @[:@38140.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@38168.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@38161.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@38162.4]
  assign RetimeWrapper_clock = clock; // @[:@38173.4]
  assign RetimeWrapper_reset = reset; // @[:@38174.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@38176.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@38175.4]
  assign RetimeWrapper_1_clock = clock; // @[:@38195.4]
  assign RetimeWrapper_1_reset = reset; // @[:@38196.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@38198.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@38197.4]
  assign RetimeWrapper_2_clock = clock; // @[:@38207.4]
  assign RetimeWrapper_2_reset = reset; // @[:@38208.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@38210.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@38209.4]
  assign RetimeWrapper_3_clock = clock; // @[:@38215.4]
  assign RetimeWrapper_3_reset = reset; // @[:@38216.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@38218.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@38217.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x382_inr_UnitPipe_kernelx382_inr_UnitPipe_concrete1( // @[:@38308.2]
  output  io_in_x364_ready, // @[:@38311.4]
  input   io_sigsIn_datapathEn // @[:@38311.4]
);
  assign io_in_x364_ready = io_sigsIn_datapathEn; // @[sm_x382_inr_UnitPipe.scala 57:18:@38323.4]
endmodule
module x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1( // @[:@38326.2]
  input         clock, // @[:@38327.4]
  input         reset, // @[:@38328.4]
  output [20:0] io_in_x211_outbuf_0_rPort_0_ofs_0, // @[:@38329.4]
  output        io_in_x211_outbuf_0_rPort_0_en_0, // @[:@38329.4]
  output        io_in_x211_outbuf_0_rPort_0_backpressure, // @[:@38329.4]
  input  [31:0] io_in_x211_outbuf_0_rPort_0_output_0, // @[:@38329.4]
  input         io_in_x362_ready, // @[:@38329.4]
  output        io_in_x362_valid, // @[:@38329.4]
  output [63:0] io_in_x362_bits_addr, // @[:@38329.4]
  output [31:0] io_in_x362_bits_size, // @[:@38329.4]
  input         io_in_x363_ready, // @[:@38329.4]
  output        io_in_x363_valid, // @[:@38329.4]
  output [31:0] io_in_x363_bits_wdata_0, // @[:@38329.4]
  output        io_in_x363_bits_wstrb, // @[:@38329.4]
  input  [63:0] io_in_x207_outdram_number, // @[:@38329.4]
  output        io_in_x364_ready, // @[:@38329.4]
  input         io_in_x364_valid, // @[:@38329.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@38329.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@38329.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@38329.4]
  input         io_sigsIn_smChildAcks_0, // @[:@38329.4]
  input         io_sigsIn_smChildAcks_1, // @[:@38329.4]
  input         io_sigsIn_smChildAcks_2, // @[:@38329.4]
  output        io_sigsOut_smDoneIn_0, // @[:@38329.4]
  output        io_sigsOut_smDoneIn_1, // @[:@38329.4]
  output        io_sigsOut_smDoneIn_2, // @[:@38329.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@38329.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@38329.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@38329.4]
  input         io_rr // @[:@38329.4]
);
  wire  x369_inr_UnitPipe_sm_clock; // @[sm_x369_inr_UnitPipe.scala 33:18:@38396.4]
  wire  x369_inr_UnitPipe_sm_reset; // @[sm_x369_inr_UnitPipe.scala 33:18:@38396.4]
  wire  x369_inr_UnitPipe_sm_io_enable; // @[sm_x369_inr_UnitPipe.scala 33:18:@38396.4]
  wire  x369_inr_UnitPipe_sm_io_done; // @[sm_x369_inr_UnitPipe.scala 33:18:@38396.4]
  wire  x369_inr_UnitPipe_sm_io_doneLatch; // @[sm_x369_inr_UnitPipe.scala 33:18:@38396.4]
  wire  x369_inr_UnitPipe_sm_io_ctrDone; // @[sm_x369_inr_UnitPipe.scala 33:18:@38396.4]
  wire  x369_inr_UnitPipe_sm_io_datapathEn; // @[sm_x369_inr_UnitPipe.scala 33:18:@38396.4]
  wire  x369_inr_UnitPipe_sm_io_ctrInc; // @[sm_x369_inr_UnitPipe.scala 33:18:@38396.4]
  wire  x369_inr_UnitPipe_sm_io_parentAck; // @[sm_x369_inr_UnitPipe.scala 33:18:@38396.4]
  wire  x369_inr_UnitPipe_sm_io_backpressure; // @[sm_x369_inr_UnitPipe.scala 33:18:@38396.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@38453.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@38453.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@38453.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@38453.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@38453.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@38461.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@38461.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@38461.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@38461.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@38461.4]
  wire  x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_in_x362_valid; // @[sm_x369_inr_UnitPipe.scala 69:24:@38491.4]
  wire [63:0] x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_in_x362_bits_addr; // @[sm_x369_inr_UnitPipe.scala 69:24:@38491.4]
  wire [31:0] x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_in_x362_bits_size; // @[sm_x369_inr_UnitPipe.scala 69:24:@38491.4]
  wire [63:0] x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_in_x207_outdram_number; // @[sm_x369_inr_UnitPipe.scala 69:24:@38491.4]
  wire  x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x369_inr_UnitPipe.scala 69:24:@38491.4]
  wire  x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x369_inr_UnitPipe.scala 69:24:@38491.4]
  wire  x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_rr; // @[sm_x369_inr_UnitPipe.scala 69:24:@38491.4]
  wire  x371_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@38559.4]
  wire  x371_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@38559.4]
  wire  x371_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@38559.4]
  wire  x371_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@38559.4]
  wire [22:0] x371_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@38559.4]
  wire  x371_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@38559.4]
  wire  x371_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@38559.4]
  wire  x378_inr_Foreach_sm_clock; // @[sm_x378_inr_Foreach.scala 33:18:@38612.4]
  wire  x378_inr_Foreach_sm_reset; // @[sm_x378_inr_Foreach.scala 33:18:@38612.4]
  wire  x378_inr_Foreach_sm_io_enable; // @[sm_x378_inr_Foreach.scala 33:18:@38612.4]
  wire  x378_inr_Foreach_sm_io_done; // @[sm_x378_inr_Foreach.scala 33:18:@38612.4]
  wire  x378_inr_Foreach_sm_io_doneLatch; // @[sm_x378_inr_Foreach.scala 33:18:@38612.4]
  wire  x378_inr_Foreach_sm_io_ctrDone; // @[sm_x378_inr_Foreach.scala 33:18:@38612.4]
  wire  x378_inr_Foreach_sm_io_datapathEn; // @[sm_x378_inr_Foreach.scala 33:18:@38612.4]
  wire  x378_inr_Foreach_sm_io_ctrInc; // @[sm_x378_inr_Foreach.scala 33:18:@38612.4]
  wire  x378_inr_Foreach_sm_io_ctrRst; // @[sm_x378_inr_Foreach.scala 33:18:@38612.4]
  wire  x378_inr_Foreach_sm_io_parentAck; // @[sm_x378_inr_Foreach.scala 33:18:@38612.4]
  wire  x378_inr_Foreach_sm_io_backpressure; // @[sm_x378_inr_Foreach.scala 33:18:@38612.4]
  wire  x378_inr_Foreach_sm_io_break; // @[sm_x378_inr_Foreach.scala 33:18:@38612.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@38640.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@38640.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@38640.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@38640.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@38640.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@38680.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@38680.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@38680.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@38680.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@38680.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@38688.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@38688.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@38688.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@38688.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@38688.4]
  wire  x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_clock; // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
  wire  x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_reset; // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
  wire [20:0] x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x211_outbuf_0_rPort_0_ofs_0; // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
  wire  x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x211_outbuf_0_rPort_0_en_0; // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
  wire  x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x211_outbuf_0_rPort_0_backpressure; // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
  wire [31:0] x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x211_outbuf_0_rPort_0_output_0; // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
  wire  x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x363_valid; // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
  wire [31:0] x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x363_bits_wdata_0; // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
  wire  x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x363_bits_wstrb; // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
  wire  x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
  wire  x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
  wire  x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
  wire [31:0] x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
  wire  x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
  wire  x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_rr; // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
  wire  x382_inr_UnitPipe_sm_clock; // @[sm_x382_inr_UnitPipe.scala 32:18:@38843.4]
  wire  x382_inr_UnitPipe_sm_reset; // @[sm_x382_inr_UnitPipe.scala 32:18:@38843.4]
  wire  x382_inr_UnitPipe_sm_io_enable; // @[sm_x382_inr_UnitPipe.scala 32:18:@38843.4]
  wire  x382_inr_UnitPipe_sm_io_done; // @[sm_x382_inr_UnitPipe.scala 32:18:@38843.4]
  wire  x382_inr_UnitPipe_sm_io_doneLatch; // @[sm_x382_inr_UnitPipe.scala 32:18:@38843.4]
  wire  x382_inr_UnitPipe_sm_io_ctrDone; // @[sm_x382_inr_UnitPipe.scala 32:18:@38843.4]
  wire  x382_inr_UnitPipe_sm_io_datapathEn; // @[sm_x382_inr_UnitPipe.scala 32:18:@38843.4]
  wire  x382_inr_UnitPipe_sm_io_ctrInc; // @[sm_x382_inr_UnitPipe.scala 32:18:@38843.4]
  wire  x382_inr_UnitPipe_sm_io_parentAck; // @[sm_x382_inr_UnitPipe.scala 32:18:@38843.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@38900.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@38900.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@38900.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@38900.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@38900.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@38908.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@38908.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@38908.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@38908.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@38908.4]
  wire  x382_inr_UnitPipe_kernelx382_inr_UnitPipe_concrete1_io_in_x364_ready; // @[sm_x382_inr_UnitPipe.scala 60:24:@38938.4]
  wire  x382_inr_UnitPipe_kernelx382_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x382_inr_UnitPipe.scala 60:24:@38938.4]
  wire  _T_359; // @[package.scala 100:49:@38424.4]
  reg  _T_362; // @[package.scala 48:56:@38425.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@38458.4 package.scala 96:25:@38459.4]
  wire  _T_381; // @[package.scala 96:25:@38466.4 package.scala 96:25:@38467.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@38469.4]
  wire  _T_454; // @[package.scala 96:25:@38645.4 package.scala 96:25:@38646.4]
  wire  _T_468; // @[package.scala 96:25:@38685.4 package.scala 96:25:@38686.4]
  wire  _T_474; // @[package.scala 96:25:@38693.4 package.scala 96:25:@38694.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@38696.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@38705.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@38706.4]
  wire  _T_547; // @[package.scala 100:49:@38871.4]
  reg  _T_550; // @[package.scala 48:56:@38872.4]
  reg [31:0] _RAND_1;
  wire  x382_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x383_outr_UnitPipe.scala 101:55:@38878.4]
  wire  _T_563; // @[package.scala 96:25:@38905.4 package.scala 96:25:@38906.4]
  wire  _T_569; // @[package.scala 96:25:@38913.4 package.scala 96:25:@38914.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@38916.4]
  wire  x382_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@38917.4]
  x369_inr_UnitPipe_sm x369_inr_UnitPipe_sm ( // @[sm_x369_inr_UnitPipe.scala 33:18:@38396.4]
    .clock(x369_inr_UnitPipe_sm_clock),
    .reset(x369_inr_UnitPipe_sm_reset),
    .io_enable(x369_inr_UnitPipe_sm_io_enable),
    .io_done(x369_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x369_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x369_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x369_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x369_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x369_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x369_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@38453.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@38461.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1 x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1 ( // @[sm_x369_inr_UnitPipe.scala 69:24:@38491.4]
    .io_in_x362_valid(x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_in_x362_valid),
    .io_in_x362_bits_addr(x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_in_x362_bits_addr),
    .io_in_x362_bits_size(x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_in_x362_bits_size),
    .io_in_x207_outdram_number(x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_in_x207_outdram_number),
    .io_sigsIn_backpressure(x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_rr)
  );
  x371_ctrchain x371_ctrchain ( // @[SpatialBlocks.scala 37:22:@38559.4]
    .clock(x371_ctrchain_clock),
    .reset(x371_ctrchain_reset),
    .io_input_reset(x371_ctrchain_io_input_reset),
    .io_input_enable(x371_ctrchain_io_input_enable),
    .io_output_counts_0(x371_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x371_ctrchain_io_output_oobs_0),
    .io_output_done(x371_ctrchain_io_output_done)
  );
  x378_inr_Foreach_sm x378_inr_Foreach_sm ( // @[sm_x378_inr_Foreach.scala 33:18:@38612.4]
    .clock(x378_inr_Foreach_sm_clock),
    .reset(x378_inr_Foreach_sm_reset),
    .io_enable(x378_inr_Foreach_sm_io_enable),
    .io_done(x378_inr_Foreach_sm_io_done),
    .io_doneLatch(x378_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x378_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x378_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x378_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x378_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x378_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x378_inr_Foreach_sm_io_backpressure),
    .io_break(x378_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@38640.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@38680.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@38688.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x378_inr_Foreach_kernelx378_inr_Foreach_concrete1 x378_inr_Foreach_kernelx378_inr_Foreach_concrete1 ( // @[sm_x378_inr_Foreach.scala 78:24:@38723.4]
    .clock(x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_clock),
    .reset(x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_reset),
    .io_in_x211_outbuf_0_rPort_0_ofs_0(x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x211_outbuf_0_rPort_0_ofs_0),
    .io_in_x211_outbuf_0_rPort_0_en_0(x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x211_outbuf_0_rPort_0_en_0),
    .io_in_x211_outbuf_0_rPort_0_backpressure(x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x211_outbuf_0_rPort_0_backpressure),
    .io_in_x211_outbuf_0_rPort_0_output_0(x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x211_outbuf_0_rPort_0_output_0),
    .io_in_x363_valid(x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x363_valid),
    .io_in_x363_bits_wdata_0(x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x363_bits_wdata_0),
    .io_in_x363_bits_wstrb(x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x363_bits_wstrb),
    .io_sigsIn_backpressure(x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_rr)
  );
  x382_inr_UnitPipe_sm x382_inr_UnitPipe_sm ( // @[sm_x382_inr_UnitPipe.scala 32:18:@38843.4]
    .clock(x382_inr_UnitPipe_sm_clock),
    .reset(x382_inr_UnitPipe_sm_reset),
    .io_enable(x382_inr_UnitPipe_sm_io_enable),
    .io_done(x382_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x382_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x382_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x382_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x382_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x382_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@38900.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@38908.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x382_inr_UnitPipe_kernelx382_inr_UnitPipe_concrete1 x382_inr_UnitPipe_kernelx382_inr_UnitPipe_concrete1 ( // @[sm_x382_inr_UnitPipe.scala 60:24:@38938.4]
    .io_in_x364_ready(x382_inr_UnitPipe_kernelx382_inr_UnitPipe_concrete1_io_in_x364_ready),
    .io_sigsIn_datapathEn(x382_inr_UnitPipe_kernelx382_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x369_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@38424.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@38458.4 package.scala 96:25:@38459.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@38466.4 package.scala 96:25:@38467.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@38469.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@38645.4 package.scala 96:25:@38646.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@38685.4 package.scala 96:25:@38686.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@38693.4 package.scala 96:25:@38694.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@38696.4]
  assign _T_479 = x378_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@38705.4]
  assign _T_480 = ~ x378_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@38706.4]
  assign _T_547 = x382_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@38871.4]
  assign x382_inr_UnitPipe_sigsIn_forwardpressure = io_in_x364_valid | x382_inr_UnitPipe_sm_io_doneLatch; // @[sm_x383_outr_UnitPipe.scala 101:55:@38878.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@38905.4 package.scala 96:25:@38906.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@38913.4 package.scala 96:25:@38914.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@38916.4]
  assign x382_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@38917.4]
  assign io_in_x211_outbuf_0_rPort_0_ofs_0 = x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x211_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@38774.4]
  assign io_in_x211_outbuf_0_rPort_0_en_0 = x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x211_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@38773.4]
  assign io_in_x211_outbuf_0_rPort_0_backpressure = x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x211_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@38772.4]
  assign io_in_x362_valid = x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_in_x362_valid; // @[sm_x369_inr_UnitPipe.scala 49:23:@38529.4]
  assign io_in_x362_bits_addr = x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_in_x362_bits_addr; // @[sm_x369_inr_UnitPipe.scala 49:23:@38528.4]
  assign io_in_x362_bits_size = x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_in_x362_bits_size; // @[sm_x369_inr_UnitPipe.scala 49:23:@38527.4]
  assign io_in_x363_valid = x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x363_valid; // @[sm_x378_inr_Foreach.scala 50:23:@38778.4]
  assign io_in_x363_bits_wdata_0 = x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x363_bits_wdata_0; // @[sm_x378_inr_Foreach.scala 50:23:@38777.4]
  assign io_in_x363_bits_wstrb = x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x363_bits_wstrb; // @[sm_x378_inr_Foreach.scala 50:23:@38776.4]
  assign io_in_x364_ready = x382_inr_UnitPipe_kernelx382_inr_UnitPipe_concrete1_io_in_x364_ready; // @[sm_x382_inr_UnitPipe.scala 46:23:@38974.4]
  assign io_sigsOut_smDoneIn_0 = x369_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@38476.4]
  assign io_sigsOut_smDoneIn_1 = x378_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@38703.4]
  assign io_sigsOut_smDoneIn_2 = x382_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@38923.4]
  assign io_sigsOut_smCtrCopyDone_0 = x369_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@38490.4]
  assign io_sigsOut_smCtrCopyDone_1 = x378_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@38722.4]
  assign io_sigsOut_smCtrCopyDone_2 = x382_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@38937.4]
  assign x369_inr_UnitPipe_sm_clock = clock; // @[:@38397.4]
  assign x369_inr_UnitPipe_sm_reset = reset; // @[:@38398.4]
  assign x369_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@38473.4]
  assign x369_inr_UnitPipe_sm_io_ctrDone = x369_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x383_outr_UnitPipe.scala 77:39:@38428.4]
  assign x369_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@38475.4]
  assign x369_inr_UnitPipe_sm_io_backpressure = io_in_x362_ready | x369_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@38447.4]
  assign RetimeWrapper_clock = clock; // @[:@38454.4]
  assign RetimeWrapper_reset = reset; // @[:@38455.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@38457.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@38456.4]
  assign RetimeWrapper_1_clock = clock; // @[:@38462.4]
  assign RetimeWrapper_1_reset = reset; // @[:@38463.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@38465.4]
  assign RetimeWrapper_1_io_in = x369_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@38464.4]
  assign x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_in_x207_outdram_number = io_in_x207_outdram_number; // @[sm_x369_inr_UnitPipe.scala 50:31:@38531.4]
  assign x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x362_ready | x369_inr_UnitPipe_sm_io_doneLatch; // @[sm_x369_inr_UnitPipe.scala 74:22:@38546.4]
  assign x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x369_inr_UnitPipe_sm_io_datapathEn; // @[sm_x369_inr_UnitPipe.scala 74:22:@38544.4]
  assign x369_inr_UnitPipe_kernelx369_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x369_inr_UnitPipe.scala 73:18:@38532.4]
  assign x371_ctrchain_clock = clock; // @[:@38560.4]
  assign x371_ctrchain_reset = reset; // @[:@38561.4]
  assign x371_ctrchain_io_input_reset = x378_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@38721.4]
  assign x371_ctrchain_io_input_enable = x378_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@38673.4 SpatialBlocks.scala 159:42:@38720.4]
  assign x378_inr_Foreach_sm_clock = clock; // @[:@38613.4]
  assign x378_inr_Foreach_sm_reset = reset; // @[:@38614.4]
  assign x378_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@38700.4]
  assign x378_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x383_outr_UnitPipe.scala 90:38:@38648.4]
  assign x378_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@38702.4]
  assign x378_inr_Foreach_sm_io_backpressure = io_in_x363_ready | x378_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@38674.4]
  assign x378_inr_Foreach_sm_io_break = 1'h0; // @[sm_x383_outr_UnitPipe.scala 94:36:@38654.4]
  assign RetimeWrapper_2_clock = clock; // @[:@38641.4]
  assign RetimeWrapper_2_reset = reset; // @[:@38642.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@38644.4]
  assign RetimeWrapper_2_io_in = x371_ctrchain_io_output_done; // @[package.scala 94:16:@38643.4]
  assign RetimeWrapper_3_clock = clock; // @[:@38681.4]
  assign RetimeWrapper_3_reset = reset; // @[:@38682.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@38684.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@38683.4]
  assign RetimeWrapper_4_clock = clock; // @[:@38689.4]
  assign RetimeWrapper_4_reset = reset; // @[:@38690.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@38692.4]
  assign RetimeWrapper_4_io_in = x378_inr_Foreach_sm_io_done; // @[package.scala 94:16:@38691.4]
  assign x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_clock = clock; // @[:@38724.4]
  assign x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_reset = reset; // @[:@38725.4]
  assign x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_in_x211_outbuf_0_rPort_0_output_0 = io_in_x211_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@38771.4]
  assign x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x363_ready | x378_inr_Foreach_sm_io_doneLatch; // @[sm_x378_inr_Foreach.scala 83:22:@38794.4]
  assign x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x378_inr_Foreach.scala 83:22:@38792.4]
  assign x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_sigsIn_break = x378_inr_Foreach_sm_io_break; // @[sm_x378_inr_Foreach.scala 83:22:@38790.4]
  assign x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x371_ctrchain_io_output_counts_0[22]}},x371_ctrchain_io_output_counts_0}; // @[sm_x378_inr_Foreach.scala 83:22:@38785.4]
  assign x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x371_ctrchain_io_output_oobs_0; // @[sm_x378_inr_Foreach.scala 83:22:@38784.4]
  assign x378_inr_Foreach_kernelx378_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x378_inr_Foreach.scala 82:18:@38780.4]
  assign x382_inr_UnitPipe_sm_clock = clock; // @[:@38844.4]
  assign x382_inr_UnitPipe_sm_reset = reset; // @[:@38845.4]
  assign x382_inr_UnitPipe_sm_io_enable = x382_inr_UnitPipe_sigsIn_baseEn & x382_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@38920.4]
  assign x382_inr_UnitPipe_sm_io_ctrDone = x382_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x383_outr_UnitPipe.scala 99:39:@38875.4]
  assign x382_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@38922.4]
  assign RetimeWrapper_5_clock = clock; // @[:@38901.4]
  assign RetimeWrapper_5_reset = reset; // @[:@38902.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@38904.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@38903.4]
  assign RetimeWrapper_6_clock = clock; // @[:@38909.4]
  assign RetimeWrapper_6_reset = reset; // @[:@38910.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@38912.4]
  assign RetimeWrapper_6_io_in = x382_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@38911.4]
  assign x382_inr_UnitPipe_kernelx382_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x382_inr_UnitPipe_sm_io_datapathEn; // @[sm_x382_inr_UnitPipe.scala 65:22:@38987.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x493_kernelx493_concrete1( // @[:@39003.2]
  input          clock, // @[:@39004.4]
  input          reset, // @[:@39005.4]
  output [20:0]  io_in_x211_outbuf_0_rPort_0_ofs_0, // @[:@39006.4]
  output         io_in_x211_outbuf_0_rPort_0_en_0, // @[:@39006.4]
  output         io_in_x211_outbuf_0_rPort_0_backpressure, // @[:@39006.4]
  input  [31:0]  io_in_x211_outbuf_0_rPort_0_output_0, // @[:@39006.4]
  input          io_in_x362_ready, // @[:@39006.4]
  output         io_in_x362_valid, // @[:@39006.4]
  output [63:0]  io_in_x362_bits_addr, // @[:@39006.4]
  output [31:0]  io_in_x362_bits_size, // @[:@39006.4]
  input          io_in_x209_TVALID, // @[:@39006.4]
  output         io_in_x209_TREADY, // @[:@39006.4]
  input  [255:0] io_in_x209_TDATA, // @[:@39006.4]
  input  [7:0]   io_in_x209_TID, // @[:@39006.4]
  input  [7:0]   io_in_x209_TDEST, // @[:@39006.4]
  input          io_in_x363_ready, // @[:@39006.4]
  output         io_in_x363_valid, // @[:@39006.4]
  output [31:0]  io_in_x363_bits_wdata_0, // @[:@39006.4]
  output         io_in_x363_bits_wstrb, // @[:@39006.4]
  input  [63:0]  io_in_x207_outdram_number, // @[:@39006.4]
  output         io_in_x210_TVALID, // @[:@39006.4]
  input          io_in_x210_TREADY, // @[:@39006.4]
  output [255:0] io_in_x210_TDATA, // @[:@39006.4]
  output         io_in_x364_ready, // @[:@39006.4]
  input          io_in_x364_valid, // @[:@39006.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@39006.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@39006.4]
  input          io_sigsIn_smChildAcks_0, // @[:@39006.4]
  input          io_sigsIn_smChildAcks_1, // @[:@39006.4]
  output         io_sigsOut_smDoneIn_0, // @[:@39006.4]
  output         io_sigsOut_smDoneIn_1, // @[:@39006.4]
  input          io_rr // @[:@39006.4]
);
  wire  x361_outr_UnitPipe_sm_clock; // @[sm_x361_outr_UnitPipe.scala 32:18:@39079.4]
  wire  x361_outr_UnitPipe_sm_reset; // @[sm_x361_outr_UnitPipe.scala 32:18:@39079.4]
  wire  x361_outr_UnitPipe_sm_io_enable; // @[sm_x361_outr_UnitPipe.scala 32:18:@39079.4]
  wire  x361_outr_UnitPipe_sm_io_done; // @[sm_x361_outr_UnitPipe.scala 32:18:@39079.4]
  wire  x361_outr_UnitPipe_sm_io_parentAck; // @[sm_x361_outr_UnitPipe.scala 32:18:@39079.4]
  wire  x361_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x361_outr_UnitPipe.scala 32:18:@39079.4]
  wire  x361_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x361_outr_UnitPipe.scala 32:18:@39079.4]
  wire  x361_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x361_outr_UnitPipe.scala 32:18:@39079.4]
  wire  x361_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x361_outr_UnitPipe.scala 32:18:@39079.4]
  wire  x361_outr_UnitPipe_sm_io_childAck_0; // @[sm_x361_outr_UnitPipe.scala 32:18:@39079.4]
  wire  x361_outr_UnitPipe_sm_io_childAck_1; // @[sm_x361_outr_UnitPipe.scala 32:18:@39079.4]
  wire  x361_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x361_outr_UnitPipe.scala 32:18:@39079.4]
  wire  x361_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x361_outr_UnitPipe.scala 32:18:@39079.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@39141.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@39141.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@39141.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@39141.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@39141.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@39149.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@39149.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@39149.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@39149.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@39149.4]
  wire  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_clock; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_reset; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x209_TVALID; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x209_TREADY; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire [255:0] x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x209_TDATA; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire [7:0] x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x209_TID; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire [7:0] x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x209_TDEST; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x210_TVALID; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x210_TREADY; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire [255:0] x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x210_TDATA; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_rr; // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
  wire  x383_outr_UnitPipe_sm_clock; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_reset; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_io_enable; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_io_done; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_io_parentAck; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_io_childAck_0; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_io_childAck_1; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_io_childAck_2; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  x383_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@39430.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@39430.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@39430.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@39430.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@39430.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@39438.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@39438.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@39438.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@39438.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@39438.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_clock; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_reset; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire [20:0] x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x211_outbuf_0_rPort_0_ofs_0; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x211_outbuf_0_rPort_0_en_0; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x211_outbuf_0_rPort_0_backpressure; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire [31:0] x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x211_outbuf_0_rPort_0_output_0; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x362_ready; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x362_valid; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire [63:0] x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x362_bits_addr; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire [31:0] x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x362_bits_size; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x363_ready; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x363_valid; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire [31:0] x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x363_bits_wdata_0; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x363_bits_wstrb; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire [63:0] x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x207_outdram_number; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x364_ready; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x364_valid; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_rr; // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
  wire  _T_408; // @[package.scala 96:25:@39146.4 package.scala 96:25:@39147.4]
  wire  _T_414; // @[package.scala 96:25:@39154.4 package.scala 96:25:@39155.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@39157.4]
  wire  _T_508; // @[package.scala 96:25:@39435.4 package.scala 96:25:@39436.4]
  wire  _T_514; // @[package.scala 96:25:@39443.4 package.scala 96:25:@39444.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@39446.4]
  x361_outr_UnitPipe_sm x361_outr_UnitPipe_sm ( // @[sm_x361_outr_UnitPipe.scala 32:18:@39079.4]
    .clock(x361_outr_UnitPipe_sm_clock),
    .reset(x361_outr_UnitPipe_sm_reset),
    .io_enable(x361_outr_UnitPipe_sm_io_enable),
    .io_done(x361_outr_UnitPipe_sm_io_done),
    .io_parentAck(x361_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x361_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x361_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x361_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x361_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x361_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x361_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x361_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x361_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@39141.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@39149.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1 x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1 ( // @[sm_x361_outr_UnitPipe.scala 87:24:@39180.4]
    .clock(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_clock),
    .reset(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_reset),
    .io_in_x209_TVALID(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x209_TVALID),
    .io_in_x209_TREADY(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x209_TREADY),
    .io_in_x209_TDATA(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x209_TDATA),
    .io_in_x209_TID(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x209_TID),
    .io_in_x209_TDEST(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x209_TDEST),
    .io_in_x210_TVALID(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x210_TVALID),
    .io_in_x210_TREADY(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x210_TREADY),
    .io_in_x210_TDATA(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x210_TDATA),
    .io_sigsIn_smEnableOuts_0(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_rr)
  );
  x383_outr_UnitPipe_sm x383_outr_UnitPipe_sm ( // @[sm_x383_outr_UnitPipe.scala 36:18:@39358.4]
    .clock(x383_outr_UnitPipe_sm_clock),
    .reset(x383_outr_UnitPipe_sm_reset),
    .io_enable(x383_outr_UnitPipe_sm_io_enable),
    .io_done(x383_outr_UnitPipe_sm_io_done),
    .io_parentAck(x383_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x383_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x383_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x383_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x383_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x383_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x383_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x383_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x383_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x383_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x383_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x383_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x383_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@39430.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@39438.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1 x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1 ( // @[sm_x383_outr_UnitPipe.scala 108:24:@39470.4]
    .clock(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_clock),
    .reset(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_reset),
    .io_in_x211_outbuf_0_rPort_0_ofs_0(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x211_outbuf_0_rPort_0_ofs_0),
    .io_in_x211_outbuf_0_rPort_0_en_0(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x211_outbuf_0_rPort_0_en_0),
    .io_in_x211_outbuf_0_rPort_0_backpressure(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x211_outbuf_0_rPort_0_backpressure),
    .io_in_x211_outbuf_0_rPort_0_output_0(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x211_outbuf_0_rPort_0_output_0),
    .io_in_x362_ready(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x362_ready),
    .io_in_x362_valid(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x362_valid),
    .io_in_x362_bits_addr(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x362_bits_addr),
    .io_in_x362_bits_size(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x362_bits_size),
    .io_in_x363_ready(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x363_ready),
    .io_in_x363_valid(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x363_valid),
    .io_in_x363_bits_wdata_0(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x363_bits_wdata_0),
    .io_in_x363_bits_wstrb(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x363_bits_wstrb),
    .io_in_x207_outdram_number(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x207_outdram_number),
    .io_in_x364_ready(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x364_ready),
    .io_in_x364_valid(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x364_valid),
    .io_sigsIn_smEnableOuts_0(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@39146.4 package.scala 96:25:@39147.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@39154.4 package.scala 96:25:@39155.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@39157.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@39435.4 package.scala 96:25:@39436.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@39443.4 package.scala 96:25:@39444.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@39446.4]
  assign io_in_x211_outbuf_0_rPort_0_ofs_0 = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x211_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@39553.4]
  assign io_in_x211_outbuf_0_rPort_0_en_0 = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x211_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@39552.4]
  assign io_in_x211_outbuf_0_rPort_0_backpressure = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x211_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@39551.4]
  assign io_in_x362_valid = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x362_valid; // @[sm_x383_outr_UnitPipe.scala 59:23:@39557.4]
  assign io_in_x362_bits_addr = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x362_bits_addr; // @[sm_x383_outr_UnitPipe.scala 59:23:@39556.4]
  assign io_in_x362_bits_size = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x362_bits_size; // @[sm_x383_outr_UnitPipe.scala 59:23:@39555.4]
  assign io_in_x209_TREADY = x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x209_TREADY; // @[sm_x361_outr_UnitPipe.scala 48:23:@39248.4]
  assign io_in_x363_valid = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x363_valid; // @[sm_x383_outr_UnitPipe.scala 60:23:@39561.4]
  assign io_in_x363_bits_wdata_0 = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x363_bits_wdata_0; // @[sm_x383_outr_UnitPipe.scala 60:23:@39560.4]
  assign io_in_x363_bits_wstrb = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x363_bits_wstrb; // @[sm_x383_outr_UnitPipe.scala 60:23:@39559.4]
  assign io_in_x210_TVALID = x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x210_TVALID; // @[sm_x361_outr_UnitPipe.scala 49:23:@39258.4]
  assign io_in_x210_TDATA = x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x210_TDATA; // @[sm_x361_outr_UnitPipe.scala 49:23:@39256.4]
  assign io_in_x364_ready = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x364_ready; // @[sm_x383_outr_UnitPipe.scala 62:23:@39566.4]
  assign io_sigsOut_smDoneIn_0 = x361_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@39164.4]
  assign io_sigsOut_smDoneIn_1 = x383_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@39453.4]
  assign x361_outr_UnitPipe_sm_clock = clock; // @[:@39080.4]
  assign x361_outr_UnitPipe_sm_reset = reset; // @[:@39081.4]
  assign x361_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@39161.4]
  assign x361_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@39163.4]
  assign x361_outr_UnitPipe_sm_io_doneIn_0 = x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@39131.4]
  assign x361_outr_UnitPipe_sm_io_doneIn_1 = x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@39132.4]
  assign x361_outr_UnitPipe_sm_io_ctrCopyDone_0 = x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@39178.4]
  assign x361_outr_UnitPipe_sm_io_ctrCopyDone_1 = x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@39179.4]
  assign RetimeWrapper_clock = clock; // @[:@39142.4]
  assign RetimeWrapper_reset = reset; // @[:@39143.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@39145.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@39144.4]
  assign RetimeWrapper_1_clock = clock; // @[:@39150.4]
  assign RetimeWrapper_1_reset = reset; // @[:@39151.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@39153.4]
  assign RetimeWrapper_1_io_in = x361_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@39152.4]
  assign x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_clock = clock; // @[:@39181.4]
  assign x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_reset = reset; // @[:@39182.4]
  assign x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x209_TVALID = io_in_x209_TVALID; // @[sm_x361_outr_UnitPipe.scala 48:23:@39249.4]
  assign x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x209_TDATA = io_in_x209_TDATA; // @[sm_x361_outr_UnitPipe.scala 48:23:@39247.4]
  assign x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x209_TID = io_in_x209_TID; // @[sm_x361_outr_UnitPipe.scala 48:23:@39243.4]
  assign x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x209_TDEST = io_in_x209_TDEST; // @[sm_x361_outr_UnitPipe.scala 48:23:@39242.4]
  assign x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_in_x210_TREADY = io_in_x210_TREADY; // @[sm_x361_outr_UnitPipe.scala 49:23:@39257.4]
  assign x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x361_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x361_outr_UnitPipe.scala 92:22:@39274.4]
  assign x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x361_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x361_outr_UnitPipe.scala 92:22:@39275.4]
  assign x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x361_outr_UnitPipe_sm_io_childAck_0; // @[sm_x361_outr_UnitPipe.scala 92:22:@39270.4]
  assign x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x361_outr_UnitPipe_sm_io_childAck_1; // @[sm_x361_outr_UnitPipe.scala 92:22:@39271.4]
  assign x361_outr_UnitPipe_kernelx361_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x361_outr_UnitPipe.scala 91:18:@39259.4]
  assign x383_outr_UnitPipe_sm_clock = clock; // @[:@39359.4]
  assign x383_outr_UnitPipe_sm_reset = reset; // @[:@39360.4]
  assign x383_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@39450.4]
  assign x383_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@39452.4]
  assign x383_outr_UnitPipe_sm_io_doneIn_0 = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@39418.4]
  assign x383_outr_UnitPipe_sm_io_doneIn_1 = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@39419.4]
  assign x383_outr_UnitPipe_sm_io_doneIn_2 = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@39420.4]
  assign x383_outr_UnitPipe_sm_io_ctrCopyDone_0 = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@39467.4]
  assign x383_outr_UnitPipe_sm_io_ctrCopyDone_1 = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@39468.4]
  assign x383_outr_UnitPipe_sm_io_ctrCopyDone_2 = x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@39469.4]
  assign RetimeWrapper_2_clock = clock; // @[:@39431.4]
  assign RetimeWrapper_2_reset = reset; // @[:@39432.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@39434.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@39433.4]
  assign RetimeWrapper_3_clock = clock; // @[:@39439.4]
  assign RetimeWrapper_3_reset = reset; // @[:@39440.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@39442.4]
  assign RetimeWrapper_3_io_in = x383_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@39441.4]
  assign x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_clock = clock; // @[:@39471.4]
  assign x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_reset = reset; // @[:@39472.4]
  assign x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x211_outbuf_0_rPort_0_output_0 = io_in_x211_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@39550.4]
  assign x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x362_ready = io_in_x362_ready; // @[sm_x383_outr_UnitPipe.scala 59:23:@39558.4]
  assign x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x363_ready = io_in_x363_ready; // @[sm_x383_outr_UnitPipe.scala 60:23:@39562.4]
  assign x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x207_outdram_number = io_in_x207_outdram_number; // @[sm_x383_outr_UnitPipe.scala 61:31:@39563.4]
  assign x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_in_x364_valid = io_in_x364_valid; // @[sm_x383_outr_UnitPipe.scala 62:23:@39565.4]
  assign x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x383_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x383_outr_UnitPipe.scala 113:22:@39589.4]
  assign x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x383_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x383_outr_UnitPipe.scala 113:22:@39590.4]
  assign x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x383_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x383_outr_UnitPipe.scala 113:22:@39591.4]
  assign x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x383_outr_UnitPipe_sm_io_childAck_0; // @[sm_x383_outr_UnitPipe.scala 113:22:@39583.4]
  assign x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x383_outr_UnitPipe_sm_io_childAck_1; // @[sm_x383_outr_UnitPipe.scala 113:22:@39584.4]
  assign x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x383_outr_UnitPipe_sm_io_childAck_2; // @[sm_x383_outr_UnitPipe.scala 113:22:@39585.4]
  assign x383_outr_UnitPipe_kernelx383_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x383_outr_UnitPipe.scala 112:18:@39567.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@39619.2]
  input          clock, // @[:@39620.4]
  input          reset, // @[:@39621.4]
  input          io_in_x362_ready, // @[:@39622.4]
  output         io_in_x362_valid, // @[:@39622.4]
  output [63:0]  io_in_x362_bits_addr, // @[:@39622.4]
  output [31:0]  io_in_x362_bits_size, // @[:@39622.4]
  input          io_in_x209_TVALID, // @[:@39622.4]
  output         io_in_x209_TREADY, // @[:@39622.4]
  input  [255:0] io_in_x209_TDATA, // @[:@39622.4]
  input  [7:0]   io_in_x209_TID, // @[:@39622.4]
  input  [7:0]   io_in_x209_TDEST, // @[:@39622.4]
  input          io_in_x363_ready, // @[:@39622.4]
  output         io_in_x363_valid, // @[:@39622.4]
  output [31:0]  io_in_x363_bits_wdata_0, // @[:@39622.4]
  output         io_in_x363_bits_wstrb, // @[:@39622.4]
  input  [63:0]  io_in_x207_outdram_number, // @[:@39622.4]
  output         io_in_x210_TVALID, // @[:@39622.4]
  input          io_in_x210_TREADY, // @[:@39622.4]
  output [255:0] io_in_x210_TDATA, // @[:@39622.4]
  output         io_in_x364_ready, // @[:@39622.4]
  input          io_in_x364_valid, // @[:@39622.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@39622.4]
  input          io_sigsIn_smChildAcks_0, // @[:@39622.4]
  output         io_sigsOut_smDoneIn_0, // @[:@39622.4]
  input          io_rr // @[:@39622.4]
);
  wire  x211_outbuf_0_clock; // @[m_x211_outbuf_0.scala 27:17:@39632.4]
  wire  x211_outbuf_0_reset; // @[m_x211_outbuf_0.scala 27:17:@39632.4]
  wire [20:0] x211_outbuf_0_io_rPort_0_ofs_0; // @[m_x211_outbuf_0.scala 27:17:@39632.4]
  wire  x211_outbuf_0_io_rPort_0_en_0; // @[m_x211_outbuf_0.scala 27:17:@39632.4]
  wire  x211_outbuf_0_io_rPort_0_backpressure; // @[m_x211_outbuf_0.scala 27:17:@39632.4]
  wire [31:0] x211_outbuf_0_io_rPort_0_output_0; // @[m_x211_outbuf_0.scala 27:17:@39632.4]
  wire  x493_sm_clock; // @[sm_x493.scala 37:18:@39690.4]
  wire  x493_sm_reset; // @[sm_x493.scala 37:18:@39690.4]
  wire  x493_sm_io_enable; // @[sm_x493.scala 37:18:@39690.4]
  wire  x493_sm_io_done; // @[sm_x493.scala 37:18:@39690.4]
  wire  x493_sm_io_ctrDone; // @[sm_x493.scala 37:18:@39690.4]
  wire  x493_sm_io_ctrInc; // @[sm_x493.scala 37:18:@39690.4]
  wire  x493_sm_io_parentAck; // @[sm_x493.scala 37:18:@39690.4]
  wire  x493_sm_io_doneIn_0; // @[sm_x493.scala 37:18:@39690.4]
  wire  x493_sm_io_doneIn_1; // @[sm_x493.scala 37:18:@39690.4]
  wire  x493_sm_io_enableOut_0; // @[sm_x493.scala 37:18:@39690.4]
  wire  x493_sm_io_enableOut_1; // @[sm_x493.scala 37:18:@39690.4]
  wire  x493_sm_io_childAck_0; // @[sm_x493.scala 37:18:@39690.4]
  wire  x493_sm_io_childAck_1; // @[sm_x493.scala 37:18:@39690.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@39757.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@39757.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@39757.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@39757.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@39757.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@39765.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@39765.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@39765.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@39765.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@39765.4]
  wire  x493_kernelx493_concrete1_clock; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_reset; // @[sm_x493.scala 102:24:@39794.4]
  wire [20:0] x493_kernelx493_concrete1_io_in_x211_outbuf_0_rPort_0_ofs_0; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_in_x211_outbuf_0_rPort_0_en_0; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_in_x211_outbuf_0_rPort_0_backpressure; // @[sm_x493.scala 102:24:@39794.4]
  wire [31:0] x493_kernelx493_concrete1_io_in_x211_outbuf_0_rPort_0_output_0; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_in_x362_ready; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_in_x362_valid; // @[sm_x493.scala 102:24:@39794.4]
  wire [63:0] x493_kernelx493_concrete1_io_in_x362_bits_addr; // @[sm_x493.scala 102:24:@39794.4]
  wire [31:0] x493_kernelx493_concrete1_io_in_x362_bits_size; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_in_x209_TVALID; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_in_x209_TREADY; // @[sm_x493.scala 102:24:@39794.4]
  wire [255:0] x493_kernelx493_concrete1_io_in_x209_TDATA; // @[sm_x493.scala 102:24:@39794.4]
  wire [7:0] x493_kernelx493_concrete1_io_in_x209_TID; // @[sm_x493.scala 102:24:@39794.4]
  wire [7:0] x493_kernelx493_concrete1_io_in_x209_TDEST; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_in_x363_ready; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_in_x363_valid; // @[sm_x493.scala 102:24:@39794.4]
  wire [31:0] x493_kernelx493_concrete1_io_in_x363_bits_wdata_0; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_in_x363_bits_wstrb; // @[sm_x493.scala 102:24:@39794.4]
  wire [63:0] x493_kernelx493_concrete1_io_in_x207_outdram_number; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_in_x210_TVALID; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_in_x210_TREADY; // @[sm_x493.scala 102:24:@39794.4]
  wire [255:0] x493_kernelx493_concrete1_io_in_x210_TDATA; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_in_x364_ready; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_in_x364_valid; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x493.scala 102:24:@39794.4]
  wire  x493_kernelx493_concrete1_io_rr; // @[sm_x493.scala 102:24:@39794.4]
  wire  _T_266; // @[package.scala 100:49:@39723.4]
  reg  _T_269; // @[package.scala 48:56:@39724.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@39762.4 package.scala 96:25:@39763.4]
  wire  _T_289; // @[package.scala 96:25:@39770.4 package.scala 96:25:@39771.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@39773.4]
  x211_outbuf_0 x211_outbuf_0 ( // @[m_x211_outbuf_0.scala 27:17:@39632.4]
    .clock(x211_outbuf_0_clock),
    .reset(x211_outbuf_0_reset),
    .io_rPort_0_ofs_0(x211_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x211_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x211_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x211_outbuf_0_io_rPort_0_output_0)
  );
  x493_sm x493_sm ( // @[sm_x493.scala 37:18:@39690.4]
    .clock(x493_sm_clock),
    .reset(x493_sm_reset),
    .io_enable(x493_sm_io_enable),
    .io_done(x493_sm_io_done),
    .io_ctrDone(x493_sm_io_ctrDone),
    .io_ctrInc(x493_sm_io_ctrInc),
    .io_parentAck(x493_sm_io_parentAck),
    .io_doneIn_0(x493_sm_io_doneIn_0),
    .io_doneIn_1(x493_sm_io_doneIn_1),
    .io_enableOut_0(x493_sm_io_enableOut_0),
    .io_enableOut_1(x493_sm_io_enableOut_1),
    .io_childAck_0(x493_sm_io_childAck_0),
    .io_childAck_1(x493_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@39757.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@39765.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x493_kernelx493_concrete1 x493_kernelx493_concrete1 ( // @[sm_x493.scala 102:24:@39794.4]
    .clock(x493_kernelx493_concrete1_clock),
    .reset(x493_kernelx493_concrete1_reset),
    .io_in_x211_outbuf_0_rPort_0_ofs_0(x493_kernelx493_concrete1_io_in_x211_outbuf_0_rPort_0_ofs_0),
    .io_in_x211_outbuf_0_rPort_0_en_0(x493_kernelx493_concrete1_io_in_x211_outbuf_0_rPort_0_en_0),
    .io_in_x211_outbuf_0_rPort_0_backpressure(x493_kernelx493_concrete1_io_in_x211_outbuf_0_rPort_0_backpressure),
    .io_in_x211_outbuf_0_rPort_0_output_0(x493_kernelx493_concrete1_io_in_x211_outbuf_0_rPort_0_output_0),
    .io_in_x362_ready(x493_kernelx493_concrete1_io_in_x362_ready),
    .io_in_x362_valid(x493_kernelx493_concrete1_io_in_x362_valid),
    .io_in_x362_bits_addr(x493_kernelx493_concrete1_io_in_x362_bits_addr),
    .io_in_x362_bits_size(x493_kernelx493_concrete1_io_in_x362_bits_size),
    .io_in_x209_TVALID(x493_kernelx493_concrete1_io_in_x209_TVALID),
    .io_in_x209_TREADY(x493_kernelx493_concrete1_io_in_x209_TREADY),
    .io_in_x209_TDATA(x493_kernelx493_concrete1_io_in_x209_TDATA),
    .io_in_x209_TID(x493_kernelx493_concrete1_io_in_x209_TID),
    .io_in_x209_TDEST(x493_kernelx493_concrete1_io_in_x209_TDEST),
    .io_in_x363_ready(x493_kernelx493_concrete1_io_in_x363_ready),
    .io_in_x363_valid(x493_kernelx493_concrete1_io_in_x363_valid),
    .io_in_x363_bits_wdata_0(x493_kernelx493_concrete1_io_in_x363_bits_wdata_0),
    .io_in_x363_bits_wstrb(x493_kernelx493_concrete1_io_in_x363_bits_wstrb),
    .io_in_x207_outdram_number(x493_kernelx493_concrete1_io_in_x207_outdram_number),
    .io_in_x210_TVALID(x493_kernelx493_concrete1_io_in_x210_TVALID),
    .io_in_x210_TREADY(x493_kernelx493_concrete1_io_in_x210_TREADY),
    .io_in_x210_TDATA(x493_kernelx493_concrete1_io_in_x210_TDATA),
    .io_in_x364_ready(x493_kernelx493_concrete1_io_in_x364_ready),
    .io_in_x364_valid(x493_kernelx493_concrete1_io_in_x364_valid),
    .io_sigsIn_smEnableOuts_0(x493_kernelx493_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x493_kernelx493_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x493_kernelx493_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x493_kernelx493_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x493_kernelx493_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x493_kernelx493_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x493_kernelx493_concrete1_io_rr)
  );
  assign _T_266 = x493_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@39723.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@39762.4 package.scala 96:25:@39763.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@39770.4 package.scala 96:25:@39771.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@39773.4]
  assign io_in_x362_valid = x493_kernelx493_concrete1_io_in_x362_valid; // @[sm_x493.scala 64:23:@39880.4]
  assign io_in_x362_bits_addr = x493_kernelx493_concrete1_io_in_x362_bits_addr; // @[sm_x493.scala 64:23:@39879.4]
  assign io_in_x362_bits_size = x493_kernelx493_concrete1_io_in_x362_bits_size; // @[sm_x493.scala 64:23:@39878.4]
  assign io_in_x209_TREADY = x493_kernelx493_concrete1_io_in_x209_TREADY; // @[sm_x493.scala 65:23:@39889.4]
  assign io_in_x363_valid = x493_kernelx493_concrete1_io_in_x363_valid; // @[sm_x493.scala 66:23:@39893.4]
  assign io_in_x363_bits_wdata_0 = x493_kernelx493_concrete1_io_in_x363_bits_wdata_0; // @[sm_x493.scala 66:23:@39892.4]
  assign io_in_x363_bits_wstrb = x493_kernelx493_concrete1_io_in_x363_bits_wstrb; // @[sm_x493.scala 66:23:@39891.4]
  assign io_in_x210_TVALID = x493_kernelx493_concrete1_io_in_x210_TVALID; // @[sm_x493.scala 68:23:@39904.4]
  assign io_in_x210_TDATA = x493_kernelx493_concrete1_io_in_x210_TDATA; // @[sm_x493.scala 68:23:@39902.4]
  assign io_in_x364_ready = x493_kernelx493_concrete1_io_in_x364_ready; // @[sm_x493.scala 69:23:@39907.4]
  assign io_sigsOut_smDoneIn_0 = x493_sm_io_done; // @[SpatialBlocks.scala 156:53:@39780.4]
  assign x211_outbuf_0_clock = clock; // @[:@39633.4]
  assign x211_outbuf_0_reset = reset; // @[:@39634.4]
  assign x211_outbuf_0_io_rPort_0_ofs_0 = x493_kernelx493_concrete1_io_in_x211_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@39876.4]
  assign x211_outbuf_0_io_rPort_0_en_0 = x493_kernelx493_concrete1_io_in_x211_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@39875.4]
  assign x211_outbuf_0_io_rPort_0_backpressure = x493_kernelx493_concrete1_io_in_x211_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@39874.4]
  assign x493_sm_clock = clock; // @[:@39691.4]
  assign x493_sm_reset = reset; // @[:@39692.4]
  assign x493_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@39777.4]
  assign x493_sm_io_ctrDone = x493_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:26:@39727.4]
  assign x493_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@39779.4]
  assign x493_sm_io_doneIn_0 = x493_kernelx493_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@39747.4]
  assign x493_sm_io_doneIn_1 = x493_kernelx493_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@39748.4]
  assign RetimeWrapper_clock = clock; // @[:@39758.4]
  assign RetimeWrapper_reset = reset; // @[:@39759.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@39761.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@39760.4]
  assign RetimeWrapper_1_clock = clock; // @[:@39766.4]
  assign RetimeWrapper_1_reset = reset; // @[:@39767.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@39769.4]
  assign RetimeWrapper_1_io_in = x493_sm_io_done; // @[package.scala 94:16:@39768.4]
  assign x493_kernelx493_concrete1_clock = clock; // @[:@39795.4]
  assign x493_kernelx493_concrete1_reset = reset; // @[:@39796.4]
  assign x493_kernelx493_concrete1_io_in_x211_outbuf_0_rPort_0_output_0 = x211_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@39873.4]
  assign x493_kernelx493_concrete1_io_in_x362_ready = io_in_x362_ready; // @[sm_x493.scala 64:23:@39881.4]
  assign x493_kernelx493_concrete1_io_in_x209_TVALID = io_in_x209_TVALID; // @[sm_x493.scala 65:23:@39890.4]
  assign x493_kernelx493_concrete1_io_in_x209_TDATA = io_in_x209_TDATA; // @[sm_x493.scala 65:23:@39888.4]
  assign x493_kernelx493_concrete1_io_in_x209_TID = io_in_x209_TID; // @[sm_x493.scala 65:23:@39884.4]
  assign x493_kernelx493_concrete1_io_in_x209_TDEST = io_in_x209_TDEST; // @[sm_x493.scala 65:23:@39883.4]
  assign x493_kernelx493_concrete1_io_in_x363_ready = io_in_x363_ready; // @[sm_x493.scala 66:23:@39894.4]
  assign x493_kernelx493_concrete1_io_in_x207_outdram_number = io_in_x207_outdram_number; // @[sm_x493.scala 67:31:@39895.4]
  assign x493_kernelx493_concrete1_io_in_x210_TREADY = io_in_x210_TREADY; // @[sm_x493.scala 68:23:@39903.4]
  assign x493_kernelx493_concrete1_io_in_x364_valid = io_in_x364_valid; // @[sm_x493.scala 69:23:@39906.4]
  assign x493_kernelx493_concrete1_io_sigsIn_smEnableOuts_0 = x493_sm_io_enableOut_0; // @[sm_x493.scala 107:22:@39918.4]
  assign x493_kernelx493_concrete1_io_sigsIn_smEnableOuts_1 = x493_sm_io_enableOut_1; // @[sm_x493.scala 107:22:@39919.4]
  assign x493_kernelx493_concrete1_io_sigsIn_smChildAcks_0 = x493_sm_io_childAck_0; // @[sm_x493.scala 107:22:@39914.4]
  assign x493_kernelx493_concrete1_io_sigsIn_smChildAcks_1 = x493_sm_io_childAck_1; // @[sm_x493.scala 107:22:@39915.4]
  assign x493_kernelx493_concrete1_io_rr = io_rr; // @[sm_x493.scala 106:18:@39908.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@39941.2]
  input          clock, // @[:@39942.4]
  input          reset, // @[:@39943.4]
  input          io_enable, // @[:@39944.4]
  output         io_done, // @[:@39944.4]
  input          io_reset, // @[:@39944.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@39944.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@39944.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@39944.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@39944.4]
  output         io_memStreams_loads_0_data_ready, // @[:@39944.4]
  input          io_memStreams_loads_0_data_valid, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@39944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@39944.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@39944.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@39944.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@39944.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@39944.4]
  input          io_memStreams_stores_0_data_ready, // @[:@39944.4]
  output         io_memStreams_stores_0_data_valid, // @[:@39944.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@39944.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@39944.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@39944.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@39944.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@39944.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@39944.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@39944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@39944.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@39944.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@39944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@39944.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@39944.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@39944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@39944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@39944.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@39944.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@39944.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@39944.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@39944.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@39944.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@39944.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@39944.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@39944.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@39944.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@39944.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@39944.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@39944.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@39944.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@39944.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@39944.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@39944.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@39944.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@39944.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@39944.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@39944.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@39944.4]
  output         io_heap_0_req_valid, // @[:@39944.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@39944.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@39944.4]
  input          io_heap_0_resp_valid, // @[:@39944.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@39944.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@39944.4]
  input  [63:0]  io_argIns_0, // @[:@39944.4]
  input  [63:0]  io_argIns_1, // @[:@39944.4]
  input          io_argOuts_0_port_ready, // @[:@39944.4]
  output         io_argOuts_0_port_valid, // @[:@39944.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@39944.4]
  input  [63:0]  io_argOuts_0_echo // @[:@39944.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@40092.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@40092.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@40092.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@40092.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@40110.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@40110.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@40110.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@40110.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@40110.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@40119.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@40119.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@40119.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@40119.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@40119.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@40119.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@40158.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@40158.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@40158.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@40158.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@40158.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@40158.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@40158.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@40158.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@40158.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@40158.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@40158.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@40190.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@40190.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@40190.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@40190.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@40190.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x362_ready; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x362_valid; // @[sm_RootController.scala 91:24:@40252.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x362_bits_addr; // @[sm_RootController.scala 91:24:@40252.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x362_bits_size; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x209_TVALID; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x209_TREADY; // @[sm_RootController.scala 91:24:@40252.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x209_TDATA; // @[sm_RootController.scala 91:24:@40252.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x209_TID; // @[sm_RootController.scala 91:24:@40252.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x209_TDEST; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x363_ready; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x363_valid; // @[sm_RootController.scala 91:24:@40252.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x363_bits_wdata_0; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x363_bits_wstrb; // @[sm_RootController.scala 91:24:@40252.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x207_outdram_number; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x210_TVALID; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x210_TREADY; // @[sm_RootController.scala 91:24:@40252.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x210_TDATA; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x364_ready; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x364_valid; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@40252.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@40252.4]
  wire  _T_599; // @[package.scala 96:25:@40115.4 package.scala 96:25:@40116.4]
  wire  _T_664; // @[Main.scala 46:50:@40186.4]
  wire  _T_665; // @[Main.scala 46:59:@40187.4]
  wire  _T_677; // @[package.scala 100:49:@40207.4]
  reg  _T_680; // @[package.scala 48:56:@40208.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@40092.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@40110.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@40119.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@40158.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@40190.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@40252.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x362_ready(RootController_kernelRootController_concrete1_io_in_x362_ready),
    .io_in_x362_valid(RootController_kernelRootController_concrete1_io_in_x362_valid),
    .io_in_x362_bits_addr(RootController_kernelRootController_concrete1_io_in_x362_bits_addr),
    .io_in_x362_bits_size(RootController_kernelRootController_concrete1_io_in_x362_bits_size),
    .io_in_x209_TVALID(RootController_kernelRootController_concrete1_io_in_x209_TVALID),
    .io_in_x209_TREADY(RootController_kernelRootController_concrete1_io_in_x209_TREADY),
    .io_in_x209_TDATA(RootController_kernelRootController_concrete1_io_in_x209_TDATA),
    .io_in_x209_TID(RootController_kernelRootController_concrete1_io_in_x209_TID),
    .io_in_x209_TDEST(RootController_kernelRootController_concrete1_io_in_x209_TDEST),
    .io_in_x363_ready(RootController_kernelRootController_concrete1_io_in_x363_ready),
    .io_in_x363_valid(RootController_kernelRootController_concrete1_io_in_x363_valid),
    .io_in_x363_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x363_bits_wdata_0),
    .io_in_x363_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x363_bits_wstrb),
    .io_in_x207_outdram_number(RootController_kernelRootController_concrete1_io_in_x207_outdram_number),
    .io_in_x210_TVALID(RootController_kernelRootController_concrete1_io_in_x210_TVALID),
    .io_in_x210_TREADY(RootController_kernelRootController_concrete1_io_in_x210_TREADY),
    .io_in_x210_TDATA(RootController_kernelRootController_concrete1_io_in_x210_TDATA),
    .io_in_x364_ready(RootController_kernelRootController_concrete1_io_in_x364_ready),
    .io_in_x364_valid(RootController_kernelRootController_concrete1_io_in_x364_valid),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@40115.4 package.scala 96:25:@40116.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@40186.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@40187.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@40207.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@40206.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x362_valid; // @[sm_RootController.scala 60:23:@40315.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x362_bits_addr; // @[sm_RootController.scala 60:23:@40314.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x362_bits_size; // @[sm_RootController.scala 60:23:@40313.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x363_valid; // @[sm_RootController.scala 62:23:@40328.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x363_bits_wdata_0; // @[sm_RootController.scala 62:23:@40327.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x363_bits_wstrb; // @[sm_RootController.scala 62:23:@40326.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x364_ready; // @[sm_RootController.scala 65:23:@40342.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x209_TREADY; // @[sm_RootController.scala 61:23:@40324.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x210_TVALID; // @[sm_RootController.scala 64:23:@40339.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x210_TDATA; // @[sm_RootController.scala 64:23:@40337.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 64:23:@40336.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 64:23:@40335.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 64:23:@40334.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 64:23:@40333.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 64:23:@40332.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 64:23:@40331.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@40093.4]
  assign SingleCounter_reset = reset; // @[:@40094.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@40108.4]
  assign RetimeWrapper_clock = clock; // @[:@40111.4]
  assign RetimeWrapper_reset = reset; // @[:@40112.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@40114.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@40113.4]
  assign SRFF_clock = clock; // @[:@40120.4]
  assign SRFF_reset = reset; // @[:@40121.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@40370.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@40204.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@40205.4]
  assign RootController_sm_clock = clock; // @[:@40159.4]
  assign RootController_sm_reset = reset; // @[:@40160.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@40203.4 SpatialBlocks.scala 140:18:@40237.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@40231.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@40211.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@40199.4 SpatialBlocks.scala 142:21:@40239.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@40228.4]
  assign RetimeWrapper_1_clock = clock; // @[:@40191.4]
  assign RetimeWrapper_1_reset = reset; // @[:@40192.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@40194.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@40193.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@40253.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@40254.4]
  assign RootController_kernelRootController_concrete1_io_in_x362_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 60:23:@40316.4]
  assign RootController_kernelRootController_concrete1_io_in_x209_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 61:23:@40325.4]
  assign RootController_kernelRootController_concrete1_io_in_x209_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 61:23:@40323.4]
  assign RootController_kernelRootController_concrete1_io_in_x209_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 61:23:@40319.4]
  assign RootController_kernelRootController_concrete1_io_in_x209_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 61:23:@40318.4]
  assign RootController_kernelRootController_concrete1_io_in_x363_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 62:23:@40329.4]
  assign RootController_kernelRootController_concrete1_io_in_x207_outdram_number = io_argIns_1; // @[sm_RootController.scala 63:31:@40330.4]
  assign RootController_kernelRootController_concrete1_io_in_x210_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 64:23:@40338.4]
  assign RootController_kernelRootController_concrete1_io_in_x364_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 65:23:@40341.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@40351.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@40349.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@40343.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module Counter( // @[:@40372.2]
  input        clock, // @[:@40373.4]
  input        reset, // @[:@40374.4]
  input        io_enable, // @[:@40375.4]
  output [5:0] io_out, // @[:@40375.4]
  output [5:0] io_next // @[:@40375.4]
);
  reg [5:0] count; // @[Counter.scala 15:22:@40377.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_17; // @[Counter.scala 17:24:@40378.4]
  wire [5:0] newCount; // @[Counter.scala 17:24:@40379.4]
  wire [5:0] _GEN_0; // @[Counter.scala 21:26:@40384.6]
  assign _T_17 = count + 6'h1; // @[Counter.scala 17:24:@40378.4]
  assign newCount = count + 6'h1; // @[Counter.scala 17:24:@40379.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@40384.6]
  assign io_out = count; // @[Counter.scala 25:10:@40387.4]
  assign io_next = count + 6'h1; // @[Counter.scala 26:11:@40388.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module SRAM_25( // @[:@40424.2]
  input         clock, // @[:@40425.4]
  input         reset, // @[:@40426.4]
  input  [5:0]  io_raddr, // @[:@40427.4]
  input         io_wen, // @[:@40427.4]
  input  [5:0]  io_waddr, // @[:@40427.4]
  input  [63:0] io_wdata_addr, // @[:@40427.4]
  input  [31:0] io_wdata_size, // @[:@40427.4]
  output [63:0] io_rdata_addr, // @[:@40427.4]
  output [31:0] io_rdata_size // @[:@40427.4]
);
  wire [95:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@40429.4]
  wire [95:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@40429.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@40429.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@40429.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@40429.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@40429.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@40429.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@40429.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@40429.4]
  wire [95:0] _T_17; // @[SRAM.scala 175:38:@40443.4]
  wire  _T_20; // @[SRAM.scala 182:49:@40448.4]
  wire  _T_21; // @[SRAM.scala 182:37:@40449.4]
  reg  _T_24; // @[SRAM.scala 182:29:@40450.4]
  reg [31:0] _RAND_0;
  reg [95:0] _T_28; // @[SRAM.scala 183:29:@40453.4]
  reg [95:0] _RAND_1;
  wire [95:0] _T_29; // @[SRAM.scala 184:22:@40455.4]
  SRAMVerilogAWS #(.DWIDTH(96), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@40429.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_17 = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:38:@40443.4]
  assign _T_20 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@40448.4]
  assign _T_21 = io_wen & _T_20; // @[SRAM.scala 182:37:@40449.4]
  assign _T_29 = _T_24 ? _T_28 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:22:@40455.4]
  assign io_rdata_addr = _T_29[95:32]; // @[SRAM.scala 184:16:@40464.4]
  assign io_rdata_size = _T_29[31:0]; // @[SRAM.scala 184:16:@40463.4]
  assign SRAMVerilogAWS_wdata = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:20:@40444.4]
  assign SRAMVerilogAWS_backpressure = 1'h1; // @[SRAM.scala 176:27:@40445.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@40441.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@40447.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@40446.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@40442.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@40440.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@40439.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_24 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _T_28 = _RAND_1[95:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_21;
    end
    if (reset) begin
      _T_28 <= 96'h0;
    end else begin
      _T_28 <= _T_17;
    end
  end
endmodule
module FIFO( // @[:@40466.2]
  input         clock, // @[:@40467.4]
  input         reset, // @[:@40468.4]
  output        io_in_ready, // @[:@40469.4]
  input         io_in_valid, // @[:@40469.4]
  input  [63:0] io_in_bits_addr, // @[:@40469.4]
  input  [31:0] io_in_bits_size, // @[:@40469.4]
  input         io_out_ready, // @[:@40469.4]
  output        io_out_valid, // @[:@40469.4]
  output [63:0] io_out_bits_addr, // @[:@40469.4]
  output [31:0] io_out_bits_size // @[:@40469.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@40865.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@40865.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@40865.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@40865.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@40865.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@40875.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@40875.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@40875.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@40875.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@40875.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@40890.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@40890.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@40890.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@40890.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@40890.4]
  wire [63:0] SRAM_io_wdata_addr; // @[FIFO.scala 73:19:@40890.4]
  wire [31:0] SRAM_io_wdata_size; // @[FIFO.scala 73:19:@40890.4]
  wire [63:0] SRAM_io_rdata_addr; // @[FIFO.scala 73:19:@40890.4]
  wire [31:0] SRAM_io_rdata_size; // @[FIFO.scala 73:19:@40890.4]
  wire  writeEn; // @[FIFO.scala 30:29:@40863.4]
  wire  readEn; // @[FIFO.scala 31:29:@40864.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@40885.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@40886.4]
  wire  _T_824; // @[FIFO.scala 45:27:@40887.4]
  wire  empty; // @[FIFO.scala 45:24:@40888.4]
  wire  full; // @[FIFO.scala 46:23:@40889.4]
  wire  _T_827; // @[FIFO.scala 83:17:@40902.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@40903.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@40865.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@40875.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_25 SRAM ( // @[FIFO.scala 73:19:@40890.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata_addr(SRAM_io_wdata_addr),
    .io_wdata_size(SRAM_io_wdata_size),
    .io_rdata_addr(SRAM_io_rdata_addr),
    .io_rdata_size(SRAM_io_rdata_size)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@40863.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@40864.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@40886.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@40887.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@40888.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@40889.4]
  assign _T_827 = writeEn != readEn; // @[FIFO.scala 83:17:@40902.4]
  assign _GEN_0 = _T_827 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@40903.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@40909.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@40907.4]
  assign io_out_bits_addr = SRAM_io_rdata_addr; // @[FIFO.scala 79:17:@40900.4]
  assign io_out_bits_size = SRAM_io_rdata_size; // @[FIFO.scala 79:17:@40899.4]
  assign enqCounter_clock = clock; // @[:@40866.4]
  assign enqCounter_reset = reset; // @[:@40867.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@40873.4]
  assign deqCounter_clock = clock; // @[:@40876.4]
  assign deqCounter_reset = reset; // @[:@40877.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@40883.4]
  assign SRAM_clock = clock; // @[:@40891.4]
  assign SRAM_reset = reset; // @[:@40892.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@40894.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@40895.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@40896.4]
  assign SRAM_io_wdata_addr = io_in_bits_addr; // @[FIFO.scala 78:16:@40898.4]
  assign SRAM_io_wdata_size = io_in_bits_size; // @[FIFO.scala 78:16:@40897.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_827) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module Counter_2( // @[:@40911.2]
  input        clock, // @[:@40912.4]
  input        reset, // @[:@40913.4]
  input        io_enable, // @[:@40914.4]
  output [3:0] io_out // @[:@40914.4]
);
  reg [3:0] count; // @[Counter.scala 15:22:@40916.4]
  reg [31:0] _RAND_0;
  wire [4:0] _T_17; // @[Counter.scala 17:24:@40917.4]
  wire [3:0] newCount; // @[Counter.scala 17:24:@40918.4]
  wire [3:0] _GEN_0; // @[Counter.scala 21:26:@40923.6]
  assign _T_17 = count + 4'h1; // @[Counter.scala 17:24:@40917.4]
  assign newCount = count + 4'h1; // @[Counter.scala 17:24:@40918.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@40923.6]
  assign io_out = count; // @[Counter.scala 25:10:@40926.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module Counter_4( // @[:@40947.2]
  input        clock, // @[:@40948.4]
  input        reset, // @[:@40949.4]
  input        io_reset, // @[:@40950.4]
  input        io_enable, // @[:@40950.4]
  input  [1:0] io_stride, // @[:@40950.4]
  output [1:0] io_out, // @[:@40950.4]
  output [1:0] io_next // @[:@40950.4]
);
  reg [1:0] count; // @[Counter.scala 15:22:@40952.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_17; // @[Counter.scala 17:24:@40953.4]
  wire [1:0] newCount; // @[Counter.scala 17:24:@40954.4]
  wire [1:0] _GEN_0; // @[Counter.scala 21:26:@40959.6]
  wire [1:0] _GEN_1; // @[Counter.scala 19:18:@40955.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@40953.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@40954.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@40959.6]
  assign _GEN_1 = io_reset ? 2'h0 : _GEN_0; // @[Counter.scala 19:18:@40955.4]
  assign io_out = count; // @[Counter.scala 25:10:@40962.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@40963.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 2'h0;
    end else begin
      if (io_reset) begin
        count <= 2'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_26( // @[:@40999.2]
  input         clock, // @[:@41000.4]
  input         reset, // @[:@41001.4]
  input  [1:0]  io_raddr, // @[:@41002.4]
  input         io_wen, // @[:@41002.4]
  input  [1:0]  io_waddr, // @[:@41002.4]
  input  [31:0] io_wdata, // @[:@41002.4]
  output [31:0] io_rdata, // @[:@41002.4]
  input         io_backpressure // @[:@41002.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@41004.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@41004.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@41004.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@41004.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@41004.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@41004.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@41004.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@41004.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@41004.4]
  wire  _T_19; // @[SRAM.scala 182:49:@41022.4]
  wire  _T_20; // @[SRAM.scala 182:37:@41023.4]
  reg  _T_23; // @[SRAM.scala 182:29:@41024.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@41026.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(4), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@41004.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@41022.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@41023.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@41031.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@41018.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@41019.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@41016.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@41021.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@41020.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@41017.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@41015.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@41014.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module FIFO_1( // @[:@41033.2]
  input         clock, // @[:@41034.4]
  input         reset, // @[:@41035.4]
  output        io_in_ready, // @[:@41036.4]
  input         io_in_valid, // @[:@41036.4]
  input  [31:0] io_in_bits, // @[:@41036.4]
  input         io_out_ready, // @[:@41036.4]
  output        io_out_valid, // @[:@41036.4]
  output [31:0] io_out_bits // @[:@41036.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@41062.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@41062.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@41062.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@41062.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@41062.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@41062.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@41062.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@41072.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@41072.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@41072.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@41072.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@41072.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@41072.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@41072.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@41087.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@41087.4]
  wire [1:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@41087.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@41087.4]
  wire [1:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@41087.4]
  wire [31:0] SRAM_io_wdata; // @[FIFO.scala 73:19:@41087.4]
  wire [31:0] SRAM_io_rdata; // @[FIFO.scala 73:19:@41087.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@41087.4]
  wire  writeEn; // @[FIFO.scala 30:29:@41060.4]
  wire  readEn; // @[FIFO.scala 31:29:@41061.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@41082.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@41083.4]
  wire  _T_104; // @[FIFO.scala 45:27:@41084.4]
  wire  empty; // @[FIFO.scala 45:24:@41085.4]
  wire  full; // @[FIFO.scala 46:23:@41086.4]
  wire  _T_107; // @[FIFO.scala 83:17:@41097.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@41098.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@41062.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@41072.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_26 SRAM ( // @[FIFO.scala 73:19:@41087.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@41060.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@41061.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@41083.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@41084.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@41085.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@41086.4]
  assign _T_107 = writeEn != readEn; // @[FIFO.scala 83:17:@41097.4]
  assign _GEN_0 = _T_107 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@41098.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@41104.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@41102.4]
  assign io_out_bits = SRAM_io_rdata; // @[FIFO.scala 79:17:@41095.4]
  assign enqCounter_clock = clock; // @[:@41063.4]
  assign enqCounter_reset = reset; // @[:@41064.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@41070.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@41071.4]
  assign deqCounter_clock = clock; // @[:@41073.4]
  assign deqCounter_reset = reset; // @[:@41074.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@41080.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@41081.4]
  assign SRAM_clock = clock; // @[:@41088.4]
  assign SRAM_reset = reset; // @[:@41089.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@41091.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@41092.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@41093.4]
  assign SRAM_io_wdata = io_in_bits; // @[FIFO.scala 78:16:@41094.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@41096.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_107) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec( // @[:@43491.2]
  input         clock, // @[:@43492.4]
  input         reset, // @[:@43493.4]
  output        io_in_ready, // @[:@43494.4]
  input         io_in_valid, // @[:@43494.4]
  input  [31:0] io_in_bits_0, // @[:@43494.4]
  input         io_out_ready, // @[:@43494.4]
  output        io_out_valid, // @[:@43494.4]
  output [31:0] io_out_bits_0, // @[:@43494.4]
  output [31:0] io_out_bits_1, // @[:@43494.4]
  output [31:0] io_out_bits_2, // @[:@43494.4]
  output [31:0] io_out_bits_3, // @[:@43494.4]
  output [31:0] io_out_bits_4, // @[:@43494.4]
  output [31:0] io_out_bits_5, // @[:@43494.4]
  output [31:0] io_out_bits_6, // @[:@43494.4]
  output [31:0] io_out_bits_7, // @[:@43494.4]
  output [31:0] io_out_bits_8, // @[:@43494.4]
  output [31:0] io_out_bits_9, // @[:@43494.4]
  output [31:0] io_out_bits_10, // @[:@43494.4]
  output [31:0] io_out_bits_11, // @[:@43494.4]
  output [31:0] io_out_bits_12, // @[:@43494.4]
  output [31:0] io_out_bits_13, // @[:@43494.4]
  output [31:0] io_out_bits_14, // @[:@43494.4]
  output [31:0] io_out_bits_15 // @[:@43494.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@43498.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@43498.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@43498.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@43498.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@43509.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@43509.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@43509.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@43509.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@43522.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@43522.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@43522.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@43522.4]
  wire [31:0] fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@43522.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@43522.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@43522.4]
  wire [31:0] fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@43522.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@43557.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@43557.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@43557.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@43557.4]
  wire [31:0] fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@43557.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@43557.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@43557.4]
  wire [31:0] fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@43557.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@43592.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@43592.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@43592.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@43592.4]
  wire [31:0] fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@43592.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@43592.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@43592.4]
  wire [31:0] fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@43592.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@43627.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@43627.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@43627.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@43627.4]
  wire [31:0] fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@43627.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@43627.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@43627.4]
  wire [31:0] fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@43627.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@43662.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@43662.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@43662.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@43662.4]
  wire [31:0] fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@43662.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@43662.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@43662.4]
  wire [31:0] fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@43662.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@43697.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@43697.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@43697.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@43697.4]
  wire [31:0] fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@43697.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@43697.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@43697.4]
  wire [31:0] fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@43697.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@43732.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@43732.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@43732.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@43732.4]
  wire [31:0] fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@43732.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@43732.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@43732.4]
  wire [31:0] fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@43732.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@43767.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@43767.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@43767.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@43767.4]
  wire [31:0] fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@43767.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@43767.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@43767.4]
  wire [31:0] fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@43767.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@43802.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@43802.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@43802.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@43802.4]
  wire [31:0] fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@43802.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@43802.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@43802.4]
  wire [31:0] fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@43802.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@43837.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@43837.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@43837.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@43837.4]
  wire [31:0] fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@43837.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@43837.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@43837.4]
  wire [31:0] fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@43837.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@43872.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@43872.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@43872.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@43872.4]
  wire [31:0] fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@43872.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@43872.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@43872.4]
  wire [31:0] fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@43872.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@43907.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@43907.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@43907.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@43907.4]
  wire [31:0] fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@43907.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@43907.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@43907.4]
  wire [31:0] fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@43907.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@43942.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@43942.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@43942.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@43942.4]
  wire [31:0] fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@43942.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@43942.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@43942.4]
  wire [31:0] fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@43942.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@43977.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@43977.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@43977.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@43977.4]
  wire [31:0] fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@43977.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@43977.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@43977.4]
  wire [31:0] fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@43977.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@44012.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@44012.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@44012.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@44012.4]
  wire [31:0] fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@44012.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@44012.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@44012.4]
  wire [31:0] fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@44012.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@44047.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@44047.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@44047.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@44047.4]
  wire [31:0] fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@44047.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@44047.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@44047.4]
  wire [31:0] fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@44047.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@43497.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@43520.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@43547.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@43582.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@43617.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@43652.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@43687.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@43722.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@43757.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@43792.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@43827.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@43862.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@43897.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@43932.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@43967.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@44002.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@44037.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@44072.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44083.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44084.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@44114.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44085.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@44114.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44086.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@44114.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44087.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@44114.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44088.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@44114.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44089.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@44114.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44090.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@44114.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44091.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@44114.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44092.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@44114.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44093.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@44114.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44094.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@44114.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44095.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@44114.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44096.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@44114.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44097.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@44114.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44098.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@44133.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@44134.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@44135.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@44136.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@44137.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@44138.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@44139.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@44140.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@44141.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@44142.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@44143.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@44144.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@44145.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@44146.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@43498.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@43509.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_1 fifos_0 ( // @[FIFOVec.scala 40:19:@43522.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_1 fifos_1 ( // @[FIFOVec.scala 40:19:@43557.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_1 fifos_2 ( // @[FIFOVec.scala 40:19:@43592.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_1 fifos_3 ( // @[FIFOVec.scala 40:19:@43627.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_1 fifos_4 ( // @[FIFOVec.scala 40:19:@43662.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_1 fifos_5 ( // @[FIFOVec.scala 40:19:@43697.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_1 fifos_6 ( // @[FIFOVec.scala 40:19:@43732.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_1 fifos_7 ( // @[FIFOVec.scala 40:19:@43767.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_1 fifos_8 ( // @[FIFOVec.scala 40:19:@43802.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_1 fifos_9 ( // @[FIFOVec.scala 40:19:@43837.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_1 fifos_10 ( // @[FIFOVec.scala 40:19:@43872.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_1 fifos_11 ( // @[FIFOVec.scala 40:19:@43907.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_1 fifos_12 ( // @[FIFOVec.scala 40:19:@43942.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_1 fifos_13 ( // @[FIFOVec.scala 40:19:@43977.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_1 fifos_14 ( // @[FIFOVec.scala 40:19:@44012.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_1 fifos_15 ( // @[FIFOVec.scala 40:19:@44047.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@43497.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@43520.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@43547.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@43582.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@43617.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@43652.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@43687.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@43722.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@43757.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@43792.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@43827.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@43862.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@43897.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@43932.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@43967.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@44002.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@44037.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@44072.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44083.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44084.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@44114.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44085.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@44114.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44086.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@44114.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44087.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@44114.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44088.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@44114.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44089.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@44114.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44090.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@44114.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44091.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@44114.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44092.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@44114.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44093.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@44114.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44094.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@44114.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44095.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@44114.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44096.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@44114.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44097.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@44114.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@44082.4 FIFOVec.scala 49:42:@44098.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@44133.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@44134.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@44135.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@44136.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@44137.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@44138.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@44139.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@44140.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@44141.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@44142.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@44143.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@44144.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@44145.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@44146.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@44115.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@44149.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@44457.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@44458.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@44459.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@44460.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@44461.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@44462.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@44463.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@44464.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@44465.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@44466.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@44467.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@44468.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@44469.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@44470.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@44471.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@44472.4]
  assign enqCounter_clock = clock; // @[:@43499.4]
  assign enqCounter_reset = reset; // @[:@43500.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@43507.4]
  assign deqCounter_clock = clock; // @[:@43510.4]
  assign deqCounter_reset = reset; // @[:@43511.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@43518.4]
  assign fifos_0_clock = clock; // @[:@43523.4]
  assign fifos_0_reset = reset; // @[:@43524.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@43550.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43552.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43556.4]
  assign fifos_1_clock = clock; // @[:@43558.4]
  assign fifos_1_reset = reset; // @[:@43559.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@43585.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43587.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43591.4]
  assign fifos_2_clock = clock; // @[:@43593.4]
  assign fifos_2_reset = reset; // @[:@43594.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@43620.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43622.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43626.4]
  assign fifos_3_clock = clock; // @[:@43628.4]
  assign fifos_3_reset = reset; // @[:@43629.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@43655.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43657.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43661.4]
  assign fifos_4_clock = clock; // @[:@43663.4]
  assign fifos_4_reset = reset; // @[:@43664.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@43690.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43692.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43696.4]
  assign fifos_5_clock = clock; // @[:@43698.4]
  assign fifos_5_reset = reset; // @[:@43699.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@43725.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43727.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43731.4]
  assign fifos_6_clock = clock; // @[:@43733.4]
  assign fifos_6_reset = reset; // @[:@43734.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@43760.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43762.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43766.4]
  assign fifos_7_clock = clock; // @[:@43768.4]
  assign fifos_7_reset = reset; // @[:@43769.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@43795.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43797.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43801.4]
  assign fifos_8_clock = clock; // @[:@43803.4]
  assign fifos_8_reset = reset; // @[:@43804.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@43830.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43832.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43836.4]
  assign fifos_9_clock = clock; // @[:@43838.4]
  assign fifos_9_reset = reset; // @[:@43839.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@43865.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43867.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43871.4]
  assign fifos_10_clock = clock; // @[:@43873.4]
  assign fifos_10_reset = reset; // @[:@43874.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@43900.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43902.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43906.4]
  assign fifos_11_clock = clock; // @[:@43908.4]
  assign fifos_11_reset = reset; // @[:@43909.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@43935.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43937.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43941.4]
  assign fifos_12_clock = clock; // @[:@43943.4]
  assign fifos_12_reset = reset; // @[:@43944.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@43970.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43972.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43976.4]
  assign fifos_13_clock = clock; // @[:@43978.4]
  assign fifos_13_reset = reset; // @[:@43979.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@44005.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44007.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44011.4]
  assign fifos_14_clock = clock; // @[:@44013.4]
  assign fifos_14_reset = reset; // @[:@44014.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@44040.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44042.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44046.4]
  assign fifos_15_clock = clock; // @[:@44048.4]
  assign fifos_15_reset = reset; // @[:@44049.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@44075.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44077.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44081.4]
endmodule
module FFRAM( // @[:@44546.2]
  input        clock, // @[:@44547.4]
  input        reset, // @[:@44548.4]
  input  [1:0] io_raddr, // @[:@44549.4]
  input        io_wen, // @[:@44549.4]
  input  [1:0] io_waddr, // @[:@44549.4]
  input        io_wdata, // @[:@44549.4]
  output       io_rdata, // @[:@44549.4]
  input        io_banks_0_wdata_valid, // @[:@44549.4]
  input        io_banks_0_wdata_bits, // @[:@44549.4]
  input        io_banks_1_wdata_valid, // @[:@44549.4]
  input        io_banks_1_wdata_bits, // @[:@44549.4]
  input        io_banks_2_wdata_valid, // @[:@44549.4]
  input        io_banks_2_wdata_bits, // @[:@44549.4]
  input        io_banks_3_wdata_valid, // @[:@44549.4]
  input        io_banks_3_wdata_bits // @[:@44549.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@44553.4]
  reg [31:0] _RAND_0;
  wire  _T_88; // @[SRAM.scala 148:37:@44554.4]
  wire  _T_89; // @[SRAM.scala 148:25:@44555.4]
  wire  _T_90; // @[SRAM.scala 148:15:@44556.4]
  wire  _T_91; // @[SRAM.scala 149:15:@44558.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@44557.4]
  reg  regs_1; // @[SRAM.scala 145:20:@44564.4]
  reg [31:0] _RAND_1;
  wire  _T_97; // @[SRAM.scala 148:37:@44565.4]
  wire  _T_98; // @[SRAM.scala 148:25:@44566.4]
  wire  _T_99; // @[SRAM.scala 148:15:@44567.4]
  wire  _T_100; // @[SRAM.scala 149:15:@44569.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@44568.4]
  reg  regs_2; // @[SRAM.scala 145:20:@44575.4]
  reg [31:0] _RAND_2;
  wire  _T_106; // @[SRAM.scala 148:37:@44576.4]
  wire  _T_107; // @[SRAM.scala 148:25:@44577.4]
  wire  _T_108; // @[SRAM.scala 148:15:@44578.4]
  wire  _T_109; // @[SRAM.scala 149:15:@44580.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@44579.4]
  reg  regs_3; // @[SRAM.scala 145:20:@44586.4]
  reg [31:0] _RAND_3;
  wire  _T_115; // @[SRAM.scala 148:37:@44587.4]
  wire  _T_116; // @[SRAM.scala 148:25:@44588.4]
  wire  _T_117; // @[SRAM.scala 148:15:@44589.4]
  wire  _T_118; // @[SRAM.scala 149:15:@44591.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@44590.4]
  wire  _GEN_5; // @[SRAM.scala 155:12:@44600.4]
  wire  _GEN_6; // @[SRAM.scala 155:12:@44600.4]
  assign _T_88 = io_waddr == 2'h0; // @[SRAM.scala 148:37:@44554.4]
  assign _T_89 = io_wen & _T_88; // @[SRAM.scala 148:25:@44555.4]
  assign _T_90 = io_banks_0_wdata_valid | _T_89; // @[SRAM.scala 148:15:@44556.4]
  assign _T_91 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44558.6]
  assign _GEN_0 = _T_90 ? _T_91 : regs_0; // @[SRAM.scala 148:48:@44557.4]
  assign _T_97 = io_waddr == 2'h1; // @[SRAM.scala 148:37:@44565.4]
  assign _T_98 = io_wen & _T_97; // @[SRAM.scala 148:25:@44566.4]
  assign _T_99 = io_banks_1_wdata_valid | _T_98; // @[SRAM.scala 148:15:@44567.4]
  assign _T_100 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44569.6]
  assign _GEN_1 = _T_99 ? _T_100 : regs_1; // @[SRAM.scala 148:48:@44568.4]
  assign _T_106 = io_waddr == 2'h2; // @[SRAM.scala 148:37:@44576.4]
  assign _T_107 = io_wen & _T_106; // @[SRAM.scala 148:25:@44577.4]
  assign _T_108 = io_banks_2_wdata_valid | _T_107; // @[SRAM.scala 148:15:@44578.4]
  assign _T_109 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44580.6]
  assign _GEN_2 = _T_108 ? _T_109 : regs_2; // @[SRAM.scala 148:48:@44579.4]
  assign _T_115 = io_waddr == 2'h3; // @[SRAM.scala 148:37:@44587.4]
  assign _T_116 = io_wen & _T_115; // @[SRAM.scala 148:25:@44588.4]
  assign _T_117 = io_banks_3_wdata_valid | _T_116; // @[SRAM.scala 148:15:@44589.4]
  assign _T_118 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44591.6]
  assign _GEN_3 = _T_117 ? _T_118 : regs_3; // @[SRAM.scala 148:48:@44590.4]
  assign _GEN_5 = 2'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@44600.4]
  assign _GEN_6 = 2'h2 == io_raddr ? regs_2 : _GEN_5; // @[SRAM.scala 155:12:@44600.4]
  assign io_rdata = 2'h3 == io_raddr ? regs_3 : _GEN_6; // @[SRAM.scala 155:12:@44600.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_90) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_99) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_108) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_117) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_17( // @[:@44602.2]
  input   clock, // @[:@44603.4]
  input   reset, // @[:@44604.4]
  output  io_in_ready, // @[:@44605.4]
  input   io_in_valid, // @[:@44605.4]
  input   io_in_bits, // @[:@44605.4]
  input   io_out_ready, // @[:@44605.4]
  output  io_out_valid, // @[:@44605.4]
  output  io_out_bits // @[:@44605.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@44631.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@44631.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@44631.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@44631.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@44631.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@44631.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@44631.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@44641.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@44641.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@44641.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@44641.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@44641.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@44641.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@44641.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@44656.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@44656.4]
  wire [1:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@44656.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@44656.4]
  wire [1:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@44656.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@44656.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@44656.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@44656.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@44656.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@44656.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@44656.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@44656.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@44656.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@44656.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@44656.4]
  wire  writeEn; // @[FIFO.scala 30:29:@44629.4]
  wire  readEn; // @[FIFO.scala 31:29:@44630.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@44651.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@44652.4]
  wire  _T_104; // @[FIFO.scala 45:27:@44653.4]
  wire  empty; // @[FIFO.scala 45:24:@44654.4]
  wire  full; // @[FIFO.scala 46:23:@44655.4]
  wire  _T_157; // @[FIFO.scala 83:17:@44742.4]
  wire  _GEN_4; // @[FIFO.scala 83:29:@44743.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@44631.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@44641.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM FFRAM ( // @[FIFO.scala 49:19:@44656.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@44629.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@44630.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@44652.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@44653.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@44654.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@44655.4]
  assign _T_157 = writeEn != readEn; // @[FIFO.scala 83:17:@44742.4]
  assign _GEN_4 = _T_157 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@44743.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@44749.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@44747.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@44681.4]
  assign enqCounter_clock = clock; // @[:@44632.4]
  assign enqCounter_reset = reset; // @[:@44633.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@44639.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@44640.4]
  assign deqCounter_clock = clock; // @[:@44642.4]
  assign deqCounter_reset = reset; // @[:@44643.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@44649.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@44650.4]
  assign FFRAM_clock = clock; // @[:@44657.4]
  assign FFRAM_reset = reset; // @[:@44658.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@44677.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@44678.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@44679.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@44680.4]
  assign FFRAM_io_banks_0_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@44683.4]
  assign FFRAM_io_banks_0_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@44682.4]
  assign FFRAM_io_banks_1_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@44686.4]
  assign FFRAM_io_banks_1_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@44685.4]
  assign FFRAM_io_banks_2_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@44689.4]
  assign FFRAM_io_banks_2_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@44688.4]
  assign FFRAM_io_banks_3_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@44692.4]
  assign FFRAM_io_banks_3_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@44691.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_157) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_1( // @[:@48366.2]
  input   clock, // @[:@48367.4]
  input   reset, // @[:@48368.4]
  output  io_in_ready, // @[:@48369.4]
  input   io_in_valid, // @[:@48369.4]
  input   io_in_bits_0, // @[:@48369.4]
  input   io_out_ready, // @[:@48369.4]
  output  io_out_valid, // @[:@48369.4]
  output  io_out_bits_0, // @[:@48369.4]
  output  io_out_bits_1, // @[:@48369.4]
  output  io_out_bits_2, // @[:@48369.4]
  output  io_out_bits_3, // @[:@48369.4]
  output  io_out_bits_4, // @[:@48369.4]
  output  io_out_bits_5, // @[:@48369.4]
  output  io_out_bits_6, // @[:@48369.4]
  output  io_out_bits_7, // @[:@48369.4]
  output  io_out_bits_8, // @[:@48369.4]
  output  io_out_bits_9, // @[:@48369.4]
  output  io_out_bits_10, // @[:@48369.4]
  output  io_out_bits_11, // @[:@48369.4]
  output  io_out_bits_12, // @[:@48369.4]
  output  io_out_bits_13, // @[:@48369.4]
  output  io_out_bits_14, // @[:@48369.4]
  output  io_out_bits_15 // @[:@48369.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@48373.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@48373.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@48373.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@48373.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@48384.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@48384.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@48384.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@48384.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@48397.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@48397.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@48397.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@48397.4]
  wire  fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@48397.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@48397.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@48397.4]
  wire  fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@48397.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@48432.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@48432.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@48432.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@48432.4]
  wire  fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@48432.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@48432.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@48432.4]
  wire  fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@48432.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@48467.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@48467.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@48467.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@48467.4]
  wire  fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@48467.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@48467.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@48467.4]
  wire  fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@48467.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@48502.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@48502.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@48502.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@48502.4]
  wire  fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@48502.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@48502.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@48502.4]
  wire  fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@48502.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@48537.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@48537.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@48537.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@48537.4]
  wire  fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@48537.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@48537.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@48537.4]
  wire  fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@48537.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@48572.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@48572.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@48572.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@48572.4]
  wire  fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@48572.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@48572.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@48572.4]
  wire  fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@48572.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@48607.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@48607.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@48607.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@48607.4]
  wire  fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@48607.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@48607.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@48607.4]
  wire  fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@48607.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@48642.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@48642.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@48642.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@48642.4]
  wire  fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@48642.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@48642.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@48642.4]
  wire  fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@48642.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@48677.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@48677.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@48677.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@48677.4]
  wire  fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@48677.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@48677.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@48677.4]
  wire  fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@48677.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@48712.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@48712.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@48712.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@48712.4]
  wire  fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@48712.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@48712.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@48712.4]
  wire  fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@48712.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@48747.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@48747.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@48747.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@48747.4]
  wire  fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@48747.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@48747.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@48747.4]
  wire  fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@48747.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@48782.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@48782.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@48782.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@48782.4]
  wire  fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@48782.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@48782.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@48782.4]
  wire  fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@48782.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@48817.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@48817.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@48817.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@48817.4]
  wire  fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@48817.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@48817.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@48817.4]
  wire  fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@48817.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@48852.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@48852.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@48852.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@48852.4]
  wire  fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@48852.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@48852.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@48852.4]
  wire  fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@48852.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@48887.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@48887.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@48887.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@48887.4]
  wire  fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@48887.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@48887.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@48887.4]
  wire  fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@48887.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@48922.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@48922.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@48922.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@48922.4]
  wire  fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@48922.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@48922.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@48922.4]
  wire  fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@48922.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@48372.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@48395.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@48422.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@48457.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@48492.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@48527.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@48562.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@48597.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@48632.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@48667.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@48702.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@48737.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@48772.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@48807.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@48842.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@48877.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@48912.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@48947.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48958.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48959.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@48989.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48960.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@48989.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48961.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@48989.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48962.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@48989.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48963.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@48989.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48964.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@48989.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48965.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@48989.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48966.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@48989.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48967.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@48989.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48968.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@48989.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48969.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@48989.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48970.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@48989.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48971.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@48989.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48972.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@48989.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48973.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@49008.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@49009.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@49010.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@49011.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@49012.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@49013.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@49014.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@49015.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@49016.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@49017.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@49018.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@49019.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@49020.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@49021.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@48373.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@48384.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_17 fifos_0 ( // @[FIFOVec.scala 40:19:@48397.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_17 fifos_1 ( // @[FIFOVec.scala 40:19:@48432.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_17 fifos_2 ( // @[FIFOVec.scala 40:19:@48467.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_17 fifos_3 ( // @[FIFOVec.scala 40:19:@48502.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_17 fifos_4 ( // @[FIFOVec.scala 40:19:@48537.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_17 fifos_5 ( // @[FIFOVec.scala 40:19:@48572.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_17 fifos_6 ( // @[FIFOVec.scala 40:19:@48607.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_17 fifos_7 ( // @[FIFOVec.scala 40:19:@48642.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_17 fifos_8 ( // @[FIFOVec.scala 40:19:@48677.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_17 fifos_9 ( // @[FIFOVec.scala 40:19:@48712.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_17 fifos_10 ( // @[FIFOVec.scala 40:19:@48747.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_17 fifos_11 ( // @[FIFOVec.scala 40:19:@48782.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_17 fifos_12 ( // @[FIFOVec.scala 40:19:@48817.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_17 fifos_13 ( // @[FIFOVec.scala 40:19:@48852.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_17 fifos_14 ( // @[FIFOVec.scala 40:19:@48887.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_17 fifos_15 ( // @[FIFOVec.scala 40:19:@48922.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@48372.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@48395.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@48422.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@48457.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@48492.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@48527.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@48562.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@48597.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@48632.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@48667.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@48702.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@48737.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@48772.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@48807.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@48842.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@48877.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@48912.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@48947.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48958.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48959.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@48989.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48960.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@48989.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48961.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@48989.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48962.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@48989.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48963.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@48989.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48964.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@48989.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48965.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@48989.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48966.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@48989.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48967.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@48989.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48968.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@48989.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48969.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@48989.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48970.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@48989.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48971.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@48989.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48972.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@48989.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@48957.4 FIFOVec.scala 49:42:@48973.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@49008.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@49009.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@49010.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@49011.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@49012.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@49013.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@49014.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@49015.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@49016.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@49017.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@49018.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@49019.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@49020.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@49021.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@48990.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@49024.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@49332.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@49333.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@49334.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@49335.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@49336.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@49337.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@49338.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@49339.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@49340.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@49341.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@49342.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@49343.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@49344.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@49345.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@49346.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@49347.4]
  assign enqCounter_clock = clock; // @[:@48374.4]
  assign enqCounter_reset = reset; // @[:@48375.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@48382.4]
  assign deqCounter_clock = clock; // @[:@48385.4]
  assign deqCounter_reset = reset; // @[:@48386.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@48393.4]
  assign fifos_0_clock = clock; // @[:@48398.4]
  assign fifos_0_reset = reset; // @[:@48399.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@48425.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48427.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48431.4]
  assign fifos_1_clock = clock; // @[:@48433.4]
  assign fifos_1_reset = reset; // @[:@48434.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@48460.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48462.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48466.4]
  assign fifos_2_clock = clock; // @[:@48468.4]
  assign fifos_2_reset = reset; // @[:@48469.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@48495.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48497.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48501.4]
  assign fifos_3_clock = clock; // @[:@48503.4]
  assign fifos_3_reset = reset; // @[:@48504.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@48530.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48532.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48536.4]
  assign fifos_4_clock = clock; // @[:@48538.4]
  assign fifos_4_reset = reset; // @[:@48539.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@48565.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48567.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48571.4]
  assign fifos_5_clock = clock; // @[:@48573.4]
  assign fifos_5_reset = reset; // @[:@48574.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@48600.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48602.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48606.4]
  assign fifos_6_clock = clock; // @[:@48608.4]
  assign fifos_6_reset = reset; // @[:@48609.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@48635.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48637.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48641.4]
  assign fifos_7_clock = clock; // @[:@48643.4]
  assign fifos_7_reset = reset; // @[:@48644.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@48670.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48672.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48676.4]
  assign fifos_8_clock = clock; // @[:@48678.4]
  assign fifos_8_reset = reset; // @[:@48679.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@48705.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48707.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48711.4]
  assign fifos_9_clock = clock; // @[:@48713.4]
  assign fifos_9_reset = reset; // @[:@48714.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@48740.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48742.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48746.4]
  assign fifos_10_clock = clock; // @[:@48748.4]
  assign fifos_10_reset = reset; // @[:@48749.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@48775.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48777.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48781.4]
  assign fifos_11_clock = clock; // @[:@48783.4]
  assign fifos_11_reset = reset; // @[:@48784.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@48810.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48812.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48816.4]
  assign fifos_12_clock = clock; // @[:@48818.4]
  assign fifos_12_reset = reset; // @[:@48819.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@48845.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48847.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48851.4]
  assign fifos_13_clock = clock; // @[:@48853.4]
  assign fifos_13_reset = reset; // @[:@48854.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@48880.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48882.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48886.4]
  assign fifos_14_clock = clock; // @[:@48888.4]
  assign fifos_14_reset = reset; // @[:@48889.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@48915.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48917.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48921.4]
  assign fifos_15_clock = clock; // @[:@48923.4]
  assign fifos_15_reset = reset; // @[:@48924.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@48950.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48952.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48956.4]
endmodule
module FIFOWidthConvert( // @[:@49349.2]
  input         clock, // @[:@49350.4]
  input         reset, // @[:@49351.4]
  output        io_in_ready, // @[:@49352.4]
  input         io_in_valid, // @[:@49352.4]
  input  [31:0] io_in_bits_data_0, // @[:@49352.4]
  input         io_in_bits_strobe, // @[:@49352.4]
  input         io_out_ready, // @[:@49352.4]
  output        io_out_valid, // @[:@49352.4]
  output [31:0] io_out_bits_data_0, // @[:@49352.4]
  output [31:0] io_out_bits_data_1, // @[:@49352.4]
  output [31:0] io_out_bits_data_2, // @[:@49352.4]
  output [31:0] io_out_bits_data_3, // @[:@49352.4]
  output [31:0] io_out_bits_data_4, // @[:@49352.4]
  output [31:0] io_out_bits_data_5, // @[:@49352.4]
  output [31:0] io_out_bits_data_6, // @[:@49352.4]
  output [31:0] io_out_bits_data_7, // @[:@49352.4]
  output [31:0] io_out_bits_data_8, // @[:@49352.4]
  output [31:0] io_out_bits_data_9, // @[:@49352.4]
  output [31:0] io_out_bits_data_10, // @[:@49352.4]
  output [31:0] io_out_bits_data_11, // @[:@49352.4]
  output [31:0] io_out_bits_data_12, // @[:@49352.4]
  output [31:0] io_out_bits_data_13, // @[:@49352.4]
  output [31:0] io_out_bits_data_14, // @[:@49352.4]
  output [31:0] io_out_bits_data_15, // @[:@49352.4]
  output [63:0] io_out_bits_strobe // @[:@49352.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 61:22:@49354.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_in_bits_0; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_ready; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_valid; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_0; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_1; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_2; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_3; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_4; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_5; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_6; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_7; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_8; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_9; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_10; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_11; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_12; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_13; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_14; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire  FIFOVec_1_io_out_bits_15; // @[FIFOWidthConvert.scala 62:26:@49395.4]
  wire [319:0] _T_55; // @[Cat.scala 30:58:@49454.4]
  wire [511:0] _T_61; // @[Cat.scala 30:58:@49460.4]
  wire [9:0] _T_108; // @[Cat.scala 30:58:@49518.4]
  wire [15:0] _T_114; // @[Cat.scala 30:58:@49524.4]
  wire  _T_115; // @[FIFOWidthConvert.scala 36:14:@49525.4]
  wire  _T_119; // @[FIFOWidthConvert.scala 36:14:@49529.4]
  wire  _T_123; // @[FIFOWidthConvert.scala 36:14:@49533.4]
  wire  _T_127; // @[FIFOWidthConvert.scala 36:14:@49537.4]
  wire  _T_131; // @[FIFOWidthConvert.scala 36:14:@49541.4]
  wire  _T_135; // @[FIFOWidthConvert.scala 36:14:@49545.4]
  wire  _T_139; // @[FIFOWidthConvert.scala 36:14:@49549.4]
  wire  _T_143; // @[FIFOWidthConvert.scala 36:14:@49553.4]
  wire  _T_147; // @[FIFOWidthConvert.scala 36:14:@49557.4]
  wire  _T_151; // @[FIFOWidthConvert.scala 36:14:@49561.4]
  wire  _T_155; // @[FIFOWidthConvert.scala 36:14:@49565.4]
  wire  _T_159; // @[FIFOWidthConvert.scala 36:14:@49569.4]
  wire  _T_163; // @[FIFOWidthConvert.scala 36:14:@49573.4]
  wire  _T_167; // @[FIFOWidthConvert.scala 36:14:@49577.4]
  wire  _T_171; // @[FIFOWidthConvert.scala 36:14:@49581.4]
  wire  _T_175; // @[FIFOWidthConvert.scala 36:14:@49585.4]
  wire [9:0] _T_257; // @[Cat.scala 30:58:@49662.4]
  wire [18:0] _T_266; // @[Cat.scala 30:58:@49671.4]
  wire [27:0] _T_275; // @[Cat.scala 30:58:@49680.4]
  wire [36:0] _T_284; // @[Cat.scala 30:58:@49689.4]
  wire [45:0] _T_293; // @[Cat.scala 30:58:@49698.4]
  wire [54:0] _T_302; // @[Cat.scala 30:58:@49707.4]
  wire [62:0] _T_310; // @[Cat.scala 30:58:@49715.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 61:22:@49354.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15)
  );
  FIFOVec_1 FIFOVec_1 ( // @[FIFOWidthConvert.scala 62:26:@49395.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid),
    .io_in_bits_0(FIFOVec_1_io_in_bits_0),
    .io_out_ready(FIFOVec_1_io_out_ready),
    .io_out_valid(FIFOVec_1_io_out_valid),
    .io_out_bits_0(FIFOVec_1_io_out_bits_0),
    .io_out_bits_1(FIFOVec_1_io_out_bits_1),
    .io_out_bits_2(FIFOVec_1_io_out_bits_2),
    .io_out_bits_3(FIFOVec_1_io_out_bits_3),
    .io_out_bits_4(FIFOVec_1_io_out_bits_4),
    .io_out_bits_5(FIFOVec_1_io_out_bits_5),
    .io_out_bits_6(FIFOVec_1_io_out_bits_6),
    .io_out_bits_7(FIFOVec_1_io_out_bits_7),
    .io_out_bits_8(FIFOVec_1_io_out_bits_8),
    .io_out_bits_9(FIFOVec_1_io_out_bits_9),
    .io_out_bits_10(FIFOVec_1_io_out_bits_10),
    .io_out_bits_11(FIFOVec_1_io_out_bits_11),
    .io_out_bits_12(FIFOVec_1_io_out_bits_12),
    .io_out_bits_13(FIFOVec_1_io_out_bits_13),
    .io_out_bits_14(FIFOVec_1_io_out_bits_14),
    .io_out_bits_15(FIFOVec_1_io_out_bits_15)
  );
  assign _T_55 = {FIFOVec_io_out_bits_15,FIFOVec_io_out_bits_14,FIFOVec_io_out_bits_13,FIFOVec_io_out_bits_12,FIFOVec_io_out_bits_11,FIFOVec_io_out_bits_10,FIFOVec_io_out_bits_9,FIFOVec_io_out_bits_8,FIFOVec_io_out_bits_7,FIFOVec_io_out_bits_6}; // @[Cat.scala 30:58:@49454.4]
  assign _T_61 = {_T_55,FIFOVec_io_out_bits_5,FIFOVec_io_out_bits_4,FIFOVec_io_out_bits_3,FIFOVec_io_out_bits_2,FIFOVec_io_out_bits_1,FIFOVec_io_out_bits_0}; // @[Cat.scala 30:58:@49460.4]
  assign _T_108 = {FIFOVec_1_io_out_bits_0,FIFOVec_1_io_out_bits_1,FIFOVec_1_io_out_bits_2,FIFOVec_1_io_out_bits_3,FIFOVec_1_io_out_bits_4,FIFOVec_1_io_out_bits_5,FIFOVec_1_io_out_bits_6,FIFOVec_1_io_out_bits_7,FIFOVec_1_io_out_bits_8,FIFOVec_1_io_out_bits_9}; // @[Cat.scala 30:58:@49518.4]
  assign _T_114 = {_T_108,FIFOVec_1_io_out_bits_10,FIFOVec_1_io_out_bits_11,FIFOVec_1_io_out_bits_12,FIFOVec_1_io_out_bits_13,FIFOVec_1_io_out_bits_14,FIFOVec_1_io_out_bits_15}; // @[Cat.scala 30:58:@49524.4]
  assign _T_115 = _T_114[0]; // @[FIFOWidthConvert.scala 36:14:@49525.4]
  assign _T_119 = _T_114[1]; // @[FIFOWidthConvert.scala 36:14:@49529.4]
  assign _T_123 = _T_114[2]; // @[FIFOWidthConvert.scala 36:14:@49533.4]
  assign _T_127 = _T_114[3]; // @[FIFOWidthConvert.scala 36:14:@49537.4]
  assign _T_131 = _T_114[4]; // @[FIFOWidthConvert.scala 36:14:@49541.4]
  assign _T_135 = _T_114[5]; // @[FIFOWidthConvert.scala 36:14:@49545.4]
  assign _T_139 = _T_114[6]; // @[FIFOWidthConvert.scala 36:14:@49549.4]
  assign _T_143 = _T_114[7]; // @[FIFOWidthConvert.scala 36:14:@49553.4]
  assign _T_147 = _T_114[8]; // @[FIFOWidthConvert.scala 36:14:@49557.4]
  assign _T_151 = _T_114[9]; // @[FIFOWidthConvert.scala 36:14:@49561.4]
  assign _T_155 = _T_114[10]; // @[FIFOWidthConvert.scala 36:14:@49565.4]
  assign _T_159 = _T_114[11]; // @[FIFOWidthConvert.scala 36:14:@49569.4]
  assign _T_163 = _T_114[12]; // @[FIFOWidthConvert.scala 36:14:@49573.4]
  assign _T_167 = _T_114[13]; // @[FIFOWidthConvert.scala 36:14:@49577.4]
  assign _T_171 = _T_114[14]; // @[FIFOWidthConvert.scala 36:14:@49581.4]
  assign _T_175 = _T_114[15]; // @[FIFOWidthConvert.scala 36:14:@49585.4]
  assign _T_257 = {_T_175,_T_175,_T_175,_T_175,_T_171,_T_171,_T_171,_T_171,_T_167,_T_167}; // @[Cat.scala 30:58:@49662.4]
  assign _T_266 = {_T_257,_T_167,_T_167,_T_163,_T_163,_T_163,_T_163,_T_159,_T_159,_T_159}; // @[Cat.scala 30:58:@49671.4]
  assign _T_275 = {_T_266,_T_159,_T_155,_T_155,_T_155,_T_155,_T_151,_T_151,_T_151,_T_151}; // @[Cat.scala 30:58:@49680.4]
  assign _T_284 = {_T_275,_T_147,_T_147,_T_147,_T_147,_T_143,_T_143,_T_143,_T_143,_T_139}; // @[Cat.scala 30:58:@49689.4]
  assign _T_293 = {_T_284,_T_139,_T_139,_T_139,_T_135,_T_135,_T_135,_T_135,_T_131,_T_131}; // @[Cat.scala 30:58:@49698.4]
  assign _T_302 = {_T_293,_T_131,_T_131,_T_127,_T_127,_T_127,_T_127,_T_123,_T_123,_T_123}; // @[Cat.scala 30:58:@49707.4]
  assign _T_310 = {_T_302,_T_123,_T_119,_T_119,_T_119,_T_119,_T_115,_T_115,_T_115}; // @[Cat.scala 30:58:@49715.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 71:17:@49444.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 72:18:@49445.4]
  assign io_out_bits_data_0 = _T_61[31:0]; // @[FIFOWidthConvert.scala 73:22:@49494.4]
  assign io_out_bits_data_1 = _T_61[63:32]; // @[FIFOWidthConvert.scala 73:22:@49495.4]
  assign io_out_bits_data_2 = _T_61[95:64]; // @[FIFOWidthConvert.scala 73:22:@49496.4]
  assign io_out_bits_data_3 = _T_61[127:96]; // @[FIFOWidthConvert.scala 73:22:@49497.4]
  assign io_out_bits_data_4 = _T_61[159:128]; // @[FIFOWidthConvert.scala 73:22:@49498.4]
  assign io_out_bits_data_5 = _T_61[191:160]; // @[FIFOWidthConvert.scala 73:22:@49499.4]
  assign io_out_bits_data_6 = _T_61[223:192]; // @[FIFOWidthConvert.scala 73:22:@49500.4]
  assign io_out_bits_data_7 = _T_61[255:224]; // @[FIFOWidthConvert.scala 73:22:@49501.4]
  assign io_out_bits_data_8 = _T_61[287:256]; // @[FIFOWidthConvert.scala 73:22:@49502.4]
  assign io_out_bits_data_9 = _T_61[319:288]; // @[FIFOWidthConvert.scala 73:22:@49503.4]
  assign io_out_bits_data_10 = _T_61[351:320]; // @[FIFOWidthConvert.scala 73:22:@49504.4]
  assign io_out_bits_data_11 = _T_61[383:352]; // @[FIFOWidthConvert.scala 73:22:@49505.4]
  assign io_out_bits_data_12 = _T_61[415:384]; // @[FIFOWidthConvert.scala 73:22:@49506.4]
  assign io_out_bits_data_13 = _T_61[447:416]; // @[FIFOWidthConvert.scala 73:22:@49507.4]
  assign io_out_bits_data_14 = _T_61[479:448]; // @[FIFOWidthConvert.scala 73:22:@49508.4]
  assign io_out_bits_data_15 = _T_61[511:480]; // @[FIFOWidthConvert.scala 73:22:@49509.4]
  assign io_out_bits_strobe = {_T_310,_T_115}; // @[FIFOWidthConvert.scala 74:24:@49717.4]
  assign FIFOVec_clock = clock; // @[:@49355.4]
  assign FIFOVec_reset = reset; // @[:@49356.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 68:22:@49441.4]
  assign FIFOVec_io_in_bits_0 = io_in_bits_data_0; // @[FIFOWidthConvert.scala 67:24:@49440.4]
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 75:23:@49718.4]
  assign FIFOVec_1_clock = clock; // @[:@49396.4]
  assign FIFOVec_1_reset = reset; // @[:@49397.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 70:26:@49443.4]
  assign FIFOVec_1_io_in_bits_0 = io_in_bits_strobe; // @[FIFOWidthConvert.scala 69:28:@49442.4]
  assign FIFOVec_1_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 76:27:@49719.4]
endmodule
module FFRAM_16( // @[:@49757.2]
  input        clock, // @[:@49758.4]
  input        reset, // @[:@49759.4]
  input  [5:0] io_raddr, // @[:@49760.4]
  input        io_wen, // @[:@49760.4]
  input  [5:0] io_waddr, // @[:@49760.4]
  input        io_wdata, // @[:@49760.4]
  output       io_rdata, // @[:@49760.4]
  input        io_banks_0_wdata_valid, // @[:@49760.4]
  input        io_banks_0_wdata_bits, // @[:@49760.4]
  input        io_banks_1_wdata_valid, // @[:@49760.4]
  input        io_banks_1_wdata_bits, // @[:@49760.4]
  input        io_banks_2_wdata_valid, // @[:@49760.4]
  input        io_banks_2_wdata_bits, // @[:@49760.4]
  input        io_banks_3_wdata_valid, // @[:@49760.4]
  input        io_banks_3_wdata_bits, // @[:@49760.4]
  input        io_banks_4_wdata_valid, // @[:@49760.4]
  input        io_banks_4_wdata_bits, // @[:@49760.4]
  input        io_banks_5_wdata_valid, // @[:@49760.4]
  input        io_banks_5_wdata_bits, // @[:@49760.4]
  input        io_banks_6_wdata_valid, // @[:@49760.4]
  input        io_banks_6_wdata_bits, // @[:@49760.4]
  input        io_banks_7_wdata_valid, // @[:@49760.4]
  input        io_banks_7_wdata_bits, // @[:@49760.4]
  input        io_banks_8_wdata_valid, // @[:@49760.4]
  input        io_banks_8_wdata_bits, // @[:@49760.4]
  input        io_banks_9_wdata_valid, // @[:@49760.4]
  input        io_banks_9_wdata_bits, // @[:@49760.4]
  input        io_banks_10_wdata_valid, // @[:@49760.4]
  input        io_banks_10_wdata_bits, // @[:@49760.4]
  input        io_banks_11_wdata_valid, // @[:@49760.4]
  input        io_banks_11_wdata_bits, // @[:@49760.4]
  input        io_banks_12_wdata_valid, // @[:@49760.4]
  input        io_banks_12_wdata_bits, // @[:@49760.4]
  input        io_banks_13_wdata_valid, // @[:@49760.4]
  input        io_banks_13_wdata_bits, // @[:@49760.4]
  input        io_banks_14_wdata_valid, // @[:@49760.4]
  input        io_banks_14_wdata_bits, // @[:@49760.4]
  input        io_banks_15_wdata_valid, // @[:@49760.4]
  input        io_banks_15_wdata_bits, // @[:@49760.4]
  input        io_banks_16_wdata_valid, // @[:@49760.4]
  input        io_banks_16_wdata_bits, // @[:@49760.4]
  input        io_banks_17_wdata_valid, // @[:@49760.4]
  input        io_banks_17_wdata_bits, // @[:@49760.4]
  input        io_banks_18_wdata_valid, // @[:@49760.4]
  input        io_banks_18_wdata_bits, // @[:@49760.4]
  input        io_banks_19_wdata_valid, // @[:@49760.4]
  input        io_banks_19_wdata_bits, // @[:@49760.4]
  input        io_banks_20_wdata_valid, // @[:@49760.4]
  input        io_banks_20_wdata_bits, // @[:@49760.4]
  input        io_banks_21_wdata_valid, // @[:@49760.4]
  input        io_banks_21_wdata_bits, // @[:@49760.4]
  input        io_banks_22_wdata_valid, // @[:@49760.4]
  input        io_banks_22_wdata_bits, // @[:@49760.4]
  input        io_banks_23_wdata_valid, // @[:@49760.4]
  input        io_banks_23_wdata_bits, // @[:@49760.4]
  input        io_banks_24_wdata_valid, // @[:@49760.4]
  input        io_banks_24_wdata_bits, // @[:@49760.4]
  input        io_banks_25_wdata_valid, // @[:@49760.4]
  input        io_banks_25_wdata_bits, // @[:@49760.4]
  input        io_banks_26_wdata_valid, // @[:@49760.4]
  input        io_banks_26_wdata_bits, // @[:@49760.4]
  input        io_banks_27_wdata_valid, // @[:@49760.4]
  input        io_banks_27_wdata_bits, // @[:@49760.4]
  input        io_banks_28_wdata_valid, // @[:@49760.4]
  input        io_banks_28_wdata_bits, // @[:@49760.4]
  input        io_banks_29_wdata_valid, // @[:@49760.4]
  input        io_banks_29_wdata_bits, // @[:@49760.4]
  input        io_banks_30_wdata_valid, // @[:@49760.4]
  input        io_banks_30_wdata_bits, // @[:@49760.4]
  input        io_banks_31_wdata_valid, // @[:@49760.4]
  input        io_banks_31_wdata_bits, // @[:@49760.4]
  input        io_banks_32_wdata_valid, // @[:@49760.4]
  input        io_banks_32_wdata_bits, // @[:@49760.4]
  input        io_banks_33_wdata_valid, // @[:@49760.4]
  input        io_banks_33_wdata_bits, // @[:@49760.4]
  input        io_banks_34_wdata_valid, // @[:@49760.4]
  input        io_banks_34_wdata_bits, // @[:@49760.4]
  input        io_banks_35_wdata_valid, // @[:@49760.4]
  input        io_banks_35_wdata_bits, // @[:@49760.4]
  input        io_banks_36_wdata_valid, // @[:@49760.4]
  input        io_banks_36_wdata_bits, // @[:@49760.4]
  input        io_banks_37_wdata_valid, // @[:@49760.4]
  input        io_banks_37_wdata_bits, // @[:@49760.4]
  input        io_banks_38_wdata_valid, // @[:@49760.4]
  input        io_banks_38_wdata_bits, // @[:@49760.4]
  input        io_banks_39_wdata_valid, // @[:@49760.4]
  input        io_banks_39_wdata_bits, // @[:@49760.4]
  input        io_banks_40_wdata_valid, // @[:@49760.4]
  input        io_banks_40_wdata_bits, // @[:@49760.4]
  input        io_banks_41_wdata_valid, // @[:@49760.4]
  input        io_banks_41_wdata_bits, // @[:@49760.4]
  input        io_banks_42_wdata_valid, // @[:@49760.4]
  input        io_banks_42_wdata_bits, // @[:@49760.4]
  input        io_banks_43_wdata_valid, // @[:@49760.4]
  input        io_banks_43_wdata_bits, // @[:@49760.4]
  input        io_banks_44_wdata_valid, // @[:@49760.4]
  input        io_banks_44_wdata_bits, // @[:@49760.4]
  input        io_banks_45_wdata_valid, // @[:@49760.4]
  input        io_banks_45_wdata_bits, // @[:@49760.4]
  input        io_banks_46_wdata_valid, // @[:@49760.4]
  input        io_banks_46_wdata_bits, // @[:@49760.4]
  input        io_banks_47_wdata_valid, // @[:@49760.4]
  input        io_banks_47_wdata_bits, // @[:@49760.4]
  input        io_banks_48_wdata_valid, // @[:@49760.4]
  input        io_banks_48_wdata_bits, // @[:@49760.4]
  input        io_banks_49_wdata_valid, // @[:@49760.4]
  input        io_banks_49_wdata_bits, // @[:@49760.4]
  input        io_banks_50_wdata_valid, // @[:@49760.4]
  input        io_banks_50_wdata_bits, // @[:@49760.4]
  input        io_banks_51_wdata_valid, // @[:@49760.4]
  input        io_banks_51_wdata_bits, // @[:@49760.4]
  input        io_banks_52_wdata_valid, // @[:@49760.4]
  input        io_banks_52_wdata_bits, // @[:@49760.4]
  input        io_banks_53_wdata_valid, // @[:@49760.4]
  input        io_banks_53_wdata_bits, // @[:@49760.4]
  input        io_banks_54_wdata_valid, // @[:@49760.4]
  input        io_banks_54_wdata_bits, // @[:@49760.4]
  input        io_banks_55_wdata_valid, // @[:@49760.4]
  input        io_banks_55_wdata_bits, // @[:@49760.4]
  input        io_banks_56_wdata_valid, // @[:@49760.4]
  input        io_banks_56_wdata_bits, // @[:@49760.4]
  input        io_banks_57_wdata_valid, // @[:@49760.4]
  input        io_banks_57_wdata_bits, // @[:@49760.4]
  input        io_banks_58_wdata_valid, // @[:@49760.4]
  input        io_banks_58_wdata_bits, // @[:@49760.4]
  input        io_banks_59_wdata_valid, // @[:@49760.4]
  input        io_banks_59_wdata_bits, // @[:@49760.4]
  input        io_banks_60_wdata_valid, // @[:@49760.4]
  input        io_banks_60_wdata_bits, // @[:@49760.4]
  input        io_banks_61_wdata_valid, // @[:@49760.4]
  input        io_banks_61_wdata_bits, // @[:@49760.4]
  input        io_banks_62_wdata_valid, // @[:@49760.4]
  input        io_banks_62_wdata_bits, // @[:@49760.4]
  input        io_banks_63_wdata_valid, // @[:@49760.4]
  input        io_banks_63_wdata_bits // @[:@49760.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@49764.4]
  reg [31:0] _RAND_0;
  wire  _T_688; // @[SRAM.scala 148:37:@49765.4]
  wire  _T_689; // @[SRAM.scala 148:25:@49766.4]
  wire  _T_690; // @[SRAM.scala 148:15:@49767.4]
  wire  _T_691; // @[SRAM.scala 149:15:@49769.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@49768.4]
  reg  regs_1; // @[SRAM.scala 145:20:@49775.4]
  reg [31:0] _RAND_1;
  wire  _T_697; // @[SRAM.scala 148:37:@49776.4]
  wire  _T_698; // @[SRAM.scala 148:25:@49777.4]
  wire  _T_699; // @[SRAM.scala 148:15:@49778.4]
  wire  _T_700; // @[SRAM.scala 149:15:@49780.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@49779.4]
  reg  regs_2; // @[SRAM.scala 145:20:@49786.4]
  reg [31:0] _RAND_2;
  wire  _T_706; // @[SRAM.scala 148:37:@49787.4]
  wire  _T_707; // @[SRAM.scala 148:25:@49788.4]
  wire  _T_708; // @[SRAM.scala 148:15:@49789.4]
  wire  _T_709; // @[SRAM.scala 149:15:@49791.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@49790.4]
  reg  regs_3; // @[SRAM.scala 145:20:@49797.4]
  reg [31:0] _RAND_3;
  wire  _T_715; // @[SRAM.scala 148:37:@49798.4]
  wire  _T_716; // @[SRAM.scala 148:25:@49799.4]
  wire  _T_717; // @[SRAM.scala 148:15:@49800.4]
  wire  _T_718; // @[SRAM.scala 149:15:@49802.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@49801.4]
  reg  regs_4; // @[SRAM.scala 145:20:@49808.4]
  reg [31:0] _RAND_4;
  wire  _T_724; // @[SRAM.scala 148:37:@49809.4]
  wire  _T_725; // @[SRAM.scala 148:25:@49810.4]
  wire  _T_726; // @[SRAM.scala 148:15:@49811.4]
  wire  _T_727; // @[SRAM.scala 149:15:@49813.6]
  wire  _GEN_4; // @[SRAM.scala 148:48:@49812.4]
  reg  regs_5; // @[SRAM.scala 145:20:@49819.4]
  reg [31:0] _RAND_5;
  wire  _T_733; // @[SRAM.scala 148:37:@49820.4]
  wire  _T_734; // @[SRAM.scala 148:25:@49821.4]
  wire  _T_735; // @[SRAM.scala 148:15:@49822.4]
  wire  _T_736; // @[SRAM.scala 149:15:@49824.6]
  wire  _GEN_5; // @[SRAM.scala 148:48:@49823.4]
  reg  regs_6; // @[SRAM.scala 145:20:@49830.4]
  reg [31:0] _RAND_6;
  wire  _T_742; // @[SRAM.scala 148:37:@49831.4]
  wire  _T_743; // @[SRAM.scala 148:25:@49832.4]
  wire  _T_744; // @[SRAM.scala 148:15:@49833.4]
  wire  _T_745; // @[SRAM.scala 149:15:@49835.6]
  wire  _GEN_6; // @[SRAM.scala 148:48:@49834.4]
  reg  regs_7; // @[SRAM.scala 145:20:@49841.4]
  reg [31:0] _RAND_7;
  wire  _T_751; // @[SRAM.scala 148:37:@49842.4]
  wire  _T_752; // @[SRAM.scala 148:25:@49843.4]
  wire  _T_753; // @[SRAM.scala 148:15:@49844.4]
  wire  _T_754; // @[SRAM.scala 149:15:@49846.6]
  wire  _GEN_7; // @[SRAM.scala 148:48:@49845.4]
  reg  regs_8; // @[SRAM.scala 145:20:@49852.4]
  reg [31:0] _RAND_8;
  wire  _T_760; // @[SRAM.scala 148:37:@49853.4]
  wire  _T_761; // @[SRAM.scala 148:25:@49854.4]
  wire  _T_762; // @[SRAM.scala 148:15:@49855.4]
  wire  _T_763; // @[SRAM.scala 149:15:@49857.6]
  wire  _GEN_8; // @[SRAM.scala 148:48:@49856.4]
  reg  regs_9; // @[SRAM.scala 145:20:@49863.4]
  reg [31:0] _RAND_9;
  wire  _T_769; // @[SRAM.scala 148:37:@49864.4]
  wire  _T_770; // @[SRAM.scala 148:25:@49865.4]
  wire  _T_771; // @[SRAM.scala 148:15:@49866.4]
  wire  _T_772; // @[SRAM.scala 149:15:@49868.6]
  wire  _GEN_9; // @[SRAM.scala 148:48:@49867.4]
  reg  regs_10; // @[SRAM.scala 145:20:@49874.4]
  reg [31:0] _RAND_10;
  wire  _T_778; // @[SRAM.scala 148:37:@49875.4]
  wire  _T_779; // @[SRAM.scala 148:25:@49876.4]
  wire  _T_780; // @[SRAM.scala 148:15:@49877.4]
  wire  _T_781; // @[SRAM.scala 149:15:@49879.6]
  wire  _GEN_10; // @[SRAM.scala 148:48:@49878.4]
  reg  regs_11; // @[SRAM.scala 145:20:@49885.4]
  reg [31:0] _RAND_11;
  wire  _T_787; // @[SRAM.scala 148:37:@49886.4]
  wire  _T_788; // @[SRAM.scala 148:25:@49887.4]
  wire  _T_789; // @[SRAM.scala 148:15:@49888.4]
  wire  _T_790; // @[SRAM.scala 149:15:@49890.6]
  wire  _GEN_11; // @[SRAM.scala 148:48:@49889.4]
  reg  regs_12; // @[SRAM.scala 145:20:@49896.4]
  reg [31:0] _RAND_12;
  wire  _T_796; // @[SRAM.scala 148:37:@49897.4]
  wire  _T_797; // @[SRAM.scala 148:25:@49898.4]
  wire  _T_798; // @[SRAM.scala 148:15:@49899.4]
  wire  _T_799; // @[SRAM.scala 149:15:@49901.6]
  wire  _GEN_12; // @[SRAM.scala 148:48:@49900.4]
  reg  regs_13; // @[SRAM.scala 145:20:@49907.4]
  reg [31:0] _RAND_13;
  wire  _T_805; // @[SRAM.scala 148:37:@49908.4]
  wire  _T_806; // @[SRAM.scala 148:25:@49909.4]
  wire  _T_807; // @[SRAM.scala 148:15:@49910.4]
  wire  _T_808; // @[SRAM.scala 149:15:@49912.6]
  wire  _GEN_13; // @[SRAM.scala 148:48:@49911.4]
  reg  regs_14; // @[SRAM.scala 145:20:@49918.4]
  reg [31:0] _RAND_14;
  wire  _T_814; // @[SRAM.scala 148:37:@49919.4]
  wire  _T_815; // @[SRAM.scala 148:25:@49920.4]
  wire  _T_816; // @[SRAM.scala 148:15:@49921.4]
  wire  _T_817; // @[SRAM.scala 149:15:@49923.6]
  wire  _GEN_14; // @[SRAM.scala 148:48:@49922.4]
  reg  regs_15; // @[SRAM.scala 145:20:@49929.4]
  reg [31:0] _RAND_15;
  wire  _T_823; // @[SRAM.scala 148:37:@49930.4]
  wire  _T_824; // @[SRAM.scala 148:25:@49931.4]
  wire  _T_825; // @[SRAM.scala 148:15:@49932.4]
  wire  _T_826; // @[SRAM.scala 149:15:@49934.6]
  wire  _GEN_15; // @[SRAM.scala 148:48:@49933.4]
  reg  regs_16; // @[SRAM.scala 145:20:@49940.4]
  reg [31:0] _RAND_16;
  wire  _T_832; // @[SRAM.scala 148:37:@49941.4]
  wire  _T_833; // @[SRAM.scala 148:25:@49942.4]
  wire  _T_834; // @[SRAM.scala 148:15:@49943.4]
  wire  _T_835; // @[SRAM.scala 149:15:@49945.6]
  wire  _GEN_16; // @[SRAM.scala 148:48:@49944.4]
  reg  regs_17; // @[SRAM.scala 145:20:@49951.4]
  reg [31:0] _RAND_17;
  wire  _T_841; // @[SRAM.scala 148:37:@49952.4]
  wire  _T_842; // @[SRAM.scala 148:25:@49953.4]
  wire  _T_843; // @[SRAM.scala 148:15:@49954.4]
  wire  _T_844; // @[SRAM.scala 149:15:@49956.6]
  wire  _GEN_17; // @[SRAM.scala 148:48:@49955.4]
  reg  regs_18; // @[SRAM.scala 145:20:@49962.4]
  reg [31:0] _RAND_18;
  wire  _T_850; // @[SRAM.scala 148:37:@49963.4]
  wire  _T_851; // @[SRAM.scala 148:25:@49964.4]
  wire  _T_852; // @[SRAM.scala 148:15:@49965.4]
  wire  _T_853; // @[SRAM.scala 149:15:@49967.6]
  wire  _GEN_18; // @[SRAM.scala 148:48:@49966.4]
  reg  regs_19; // @[SRAM.scala 145:20:@49973.4]
  reg [31:0] _RAND_19;
  wire  _T_859; // @[SRAM.scala 148:37:@49974.4]
  wire  _T_860; // @[SRAM.scala 148:25:@49975.4]
  wire  _T_861; // @[SRAM.scala 148:15:@49976.4]
  wire  _T_862; // @[SRAM.scala 149:15:@49978.6]
  wire  _GEN_19; // @[SRAM.scala 148:48:@49977.4]
  reg  regs_20; // @[SRAM.scala 145:20:@49984.4]
  reg [31:0] _RAND_20;
  wire  _T_868; // @[SRAM.scala 148:37:@49985.4]
  wire  _T_869; // @[SRAM.scala 148:25:@49986.4]
  wire  _T_870; // @[SRAM.scala 148:15:@49987.4]
  wire  _T_871; // @[SRAM.scala 149:15:@49989.6]
  wire  _GEN_20; // @[SRAM.scala 148:48:@49988.4]
  reg  regs_21; // @[SRAM.scala 145:20:@49995.4]
  reg [31:0] _RAND_21;
  wire  _T_877; // @[SRAM.scala 148:37:@49996.4]
  wire  _T_878; // @[SRAM.scala 148:25:@49997.4]
  wire  _T_879; // @[SRAM.scala 148:15:@49998.4]
  wire  _T_880; // @[SRAM.scala 149:15:@50000.6]
  wire  _GEN_21; // @[SRAM.scala 148:48:@49999.4]
  reg  regs_22; // @[SRAM.scala 145:20:@50006.4]
  reg [31:0] _RAND_22;
  wire  _T_886; // @[SRAM.scala 148:37:@50007.4]
  wire  _T_887; // @[SRAM.scala 148:25:@50008.4]
  wire  _T_888; // @[SRAM.scala 148:15:@50009.4]
  wire  _T_889; // @[SRAM.scala 149:15:@50011.6]
  wire  _GEN_22; // @[SRAM.scala 148:48:@50010.4]
  reg  regs_23; // @[SRAM.scala 145:20:@50017.4]
  reg [31:0] _RAND_23;
  wire  _T_895; // @[SRAM.scala 148:37:@50018.4]
  wire  _T_896; // @[SRAM.scala 148:25:@50019.4]
  wire  _T_897; // @[SRAM.scala 148:15:@50020.4]
  wire  _T_898; // @[SRAM.scala 149:15:@50022.6]
  wire  _GEN_23; // @[SRAM.scala 148:48:@50021.4]
  reg  regs_24; // @[SRAM.scala 145:20:@50028.4]
  reg [31:0] _RAND_24;
  wire  _T_904; // @[SRAM.scala 148:37:@50029.4]
  wire  _T_905; // @[SRAM.scala 148:25:@50030.4]
  wire  _T_906; // @[SRAM.scala 148:15:@50031.4]
  wire  _T_907; // @[SRAM.scala 149:15:@50033.6]
  wire  _GEN_24; // @[SRAM.scala 148:48:@50032.4]
  reg  regs_25; // @[SRAM.scala 145:20:@50039.4]
  reg [31:0] _RAND_25;
  wire  _T_913; // @[SRAM.scala 148:37:@50040.4]
  wire  _T_914; // @[SRAM.scala 148:25:@50041.4]
  wire  _T_915; // @[SRAM.scala 148:15:@50042.4]
  wire  _T_916; // @[SRAM.scala 149:15:@50044.6]
  wire  _GEN_25; // @[SRAM.scala 148:48:@50043.4]
  reg  regs_26; // @[SRAM.scala 145:20:@50050.4]
  reg [31:0] _RAND_26;
  wire  _T_922; // @[SRAM.scala 148:37:@50051.4]
  wire  _T_923; // @[SRAM.scala 148:25:@50052.4]
  wire  _T_924; // @[SRAM.scala 148:15:@50053.4]
  wire  _T_925; // @[SRAM.scala 149:15:@50055.6]
  wire  _GEN_26; // @[SRAM.scala 148:48:@50054.4]
  reg  regs_27; // @[SRAM.scala 145:20:@50061.4]
  reg [31:0] _RAND_27;
  wire  _T_931; // @[SRAM.scala 148:37:@50062.4]
  wire  _T_932; // @[SRAM.scala 148:25:@50063.4]
  wire  _T_933; // @[SRAM.scala 148:15:@50064.4]
  wire  _T_934; // @[SRAM.scala 149:15:@50066.6]
  wire  _GEN_27; // @[SRAM.scala 148:48:@50065.4]
  reg  regs_28; // @[SRAM.scala 145:20:@50072.4]
  reg [31:0] _RAND_28;
  wire  _T_940; // @[SRAM.scala 148:37:@50073.4]
  wire  _T_941; // @[SRAM.scala 148:25:@50074.4]
  wire  _T_942; // @[SRAM.scala 148:15:@50075.4]
  wire  _T_943; // @[SRAM.scala 149:15:@50077.6]
  wire  _GEN_28; // @[SRAM.scala 148:48:@50076.4]
  reg  regs_29; // @[SRAM.scala 145:20:@50083.4]
  reg [31:0] _RAND_29;
  wire  _T_949; // @[SRAM.scala 148:37:@50084.4]
  wire  _T_950; // @[SRAM.scala 148:25:@50085.4]
  wire  _T_951; // @[SRAM.scala 148:15:@50086.4]
  wire  _T_952; // @[SRAM.scala 149:15:@50088.6]
  wire  _GEN_29; // @[SRAM.scala 148:48:@50087.4]
  reg  regs_30; // @[SRAM.scala 145:20:@50094.4]
  reg [31:0] _RAND_30;
  wire  _T_958; // @[SRAM.scala 148:37:@50095.4]
  wire  _T_959; // @[SRAM.scala 148:25:@50096.4]
  wire  _T_960; // @[SRAM.scala 148:15:@50097.4]
  wire  _T_961; // @[SRAM.scala 149:15:@50099.6]
  wire  _GEN_30; // @[SRAM.scala 148:48:@50098.4]
  reg  regs_31; // @[SRAM.scala 145:20:@50105.4]
  reg [31:0] _RAND_31;
  wire  _T_967; // @[SRAM.scala 148:37:@50106.4]
  wire  _T_968; // @[SRAM.scala 148:25:@50107.4]
  wire  _T_969; // @[SRAM.scala 148:15:@50108.4]
  wire  _T_970; // @[SRAM.scala 149:15:@50110.6]
  wire  _GEN_31; // @[SRAM.scala 148:48:@50109.4]
  reg  regs_32; // @[SRAM.scala 145:20:@50116.4]
  reg [31:0] _RAND_32;
  wire  _T_976; // @[SRAM.scala 148:37:@50117.4]
  wire  _T_977; // @[SRAM.scala 148:25:@50118.4]
  wire  _T_978; // @[SRAM.scala 148:15:@50119.4]
  wire  _T_979; // @[SRAM.scala 149:15:@50121.6]
  wire  _GEN_32; // @[SRAM.scala 148:48:@50120.4]
  reg  regs_33; // @[SRAM.scala 145:20:@50127.4]
  reg [31:0] _RAND_33;
  wire  _T_985; // @[SRAM.scala 148:37:@50128.4]
  wire  _T_986; // @[SRAM.scala 148:25:@50129.4]
  wire  _T_987; // @[SRAM.scala 148:15:@50130.4]
  wire  _T_988; // @[SRAM.scala 149:15:@50132.6]
  wire  _GEN_33; // @[SRAM.scala 148:48:@50131.4]
  reg  regs_34; // @[SRAM.scala 145:20:@50138.4]
  reg [31:0] _RAND_34;
  wire  _T_994; // @[SRAM.scala 148:37:@50139.4]
  wire  _T_995; // @[SRAM.scala 148:25:@50140.4]
  wire  _T_996; // @[SRAM.scala 148:15:@50141.4]
  wire  _T_997; // @[SRAM.scala 149:15:@50143.6]
  wire  _GEN_34; // @[SRAM.scala 148:48:@50142.4]
  reg  regs_35; // @[SRAM.scala 145:20:@50149.4]
  reg [31:0] _RAND_35;
  wire  _T_1003; // @[SRAM.scala 148:37:@50150.4]
  wire  _T_1004; // @[SRAM.scala 148:25:@50151.4]
  wire  _T_1005; // @[SRAM.scala 148:15:@50152.4]
  wire  _T_1006; // @[SRAM.scala 149:15:@50154.6]
  wire  _GEN_35; // @[SRAM.scala 148:48:@50153.4]
  reg  regs_36; // @[SRAM.scala 145:20:@50160.4]
  reg [31:0] _RAND_36;
  wire  _T_1012; // @[SRAM.scala 148:37:@50161.4]
  wire  _T_1013; // @[SRAM.scala 148:25:@50162.4]
  wire  _T_1014; // @[SRAM.scala 148:15:@50163.4]
  wire  _T_1015; // @[SRAM.scala 149:15:@50165.6]
  wire  _GEN_36; // @[SRAM.scala 148:48:@50164.4]
  reg  regs_37; // @[SRAM.scala 145:20:@50171.4]
  reg [31:0] _RAND_37;
  wire  _T_1021; // @[SRAM.scala 148:37:@50172.4]
  wire  _T_1022; // @[SRAM.scala 148:25:@50173.4]
  wire  _T_1023; // @[SRAM.scala 148:15:@50174.4]
  wire  _T_1024; // @[SRAM.scala 149:15:@50176.6]
  wire  _GEN_37; // @[SRAM.scala 148:48:@50175.4]
  reg  regs_38; // @[SRAM.scala 145:20:@50182.4]
  reg [31:0] _RAND_38;
  wire  _T_1030; // @[SRAM.scala 148:37:@50183.4]
  wire  _T_1031; // @[SRAM.scala 148:25:@50184.4]
  wire  _T_1032; // @[SRAM.scala 148:15:@50185.4]
  wire  _T_1033; // @[SRAM.scala 149:15:@50187.6]
  wire  _GEN_38; // @[SRAM.scala 148:48:@50186.4]
  reg  regs_39; // @[SRAM.scala 145:20:@50193.4]
  reg [31:0] _RAND_39;
  wire  _T_1039; // @[SRAM.scala 148:37:@50194.4]
  wire  _T_1040; // @[SRAM.scala 148:25:@50195.4]
  wire  _T_1041; // @[SRAM.scala 148:15:@50196.4]
  wire  _T_1042; // @[SRAM.scala 149:15:@50198.6]
  wire  _GEN_39; // @[SRAM.scala 148:48:@50197.4]
  reg  regs_40; // @[SRAM.scala 145:20:@50204.4]
  reg [31:0] _RAND_40;
  wire  _T_1048; // @[SRAM.scala 148:37:@50205.4]
  wire  _T_1049; // @[SRAM.scala 148:25:@50206.4]
  wire  _T_1050; // @[SRAM.scala 148:15:@50207.4]
  wire  _T_1051; // @[SRAM.scala 149:15:@50209.6]
  wire  _GEN_40; // @[SRAM.scala 148:48:@50208.4]
  reg  regs_41; // @[SRAM.scala 145:20:@50215.4]
  reg [31:0] _RAND_41;
  wire  _T_1057; // @[SRAM.scala 148:37:@50216.4]
  wire  _T_1058; // @[SRAM.scala 148:25:@50217.4]
  wire  _T_1059; // @[SRAM.scala 148:15:@50218.4]
  wire  _T_1060; // @[SRAM.scala 149:15:@50220.6]
  wire  _GEN_41; // @[SRAM.scala 148:48:@50219.4]
  reg  regs_42; // @[SRAM.scala 145:20:@50226.4]
  reg [31:0] _RAND_42;
  wire  _T_1066; // @[SRAM.scala 148:37:@50227.4]
  wire  _T_1067; // @[SRAM.scala 148:25:@50228.4]
  wire  _T_1068; // @[SRAM.scala 148:15:@50229.4]
  wire  _T_1069; // @[SRAM.scala 149:15:@50231.6]
  wire  _GEN_42; // @[SRAM.scala 148:48:@50230.4]
  reg  regs_43; // @[SRAM.scala 145:20:@50237.4]
  reg [31:0] _RAND_43;
  wire  _T_1075; // @[SRAM.scala 148:37:@50238.4]
  wire  _T_1076; // @[SRAM.scala 148:25:@50239.4]
  wire  _T_1077; // @[SRAM.scala 148:15:@50240.4]
  wire  _T_1078; // @[SRAM.scala 149:15:@50242.6]
  wire  _GEN_43; // @[SRAM.scala 148:48:@50241.4]
  reg  regs_44; // @[SRAM.scala 145:20:@50248.4]
  reg [31:0] _RAND_44;
  wire  _T_1084; // @[SRAM.scala 148:37:@50249.4]
  wire  _T_1085; // @[SRAM.scala 148:25:@50250.4]
  wire  _T_1086; // @[SRAM.scala 148:15:@50251.4]
  wire  _T_1087; // @[SRAM.scala 149:15:@50253.6]
  wire  _GEN_44; // @[SRAM.scala 148:48:@50252.4]
  reg  regs_45; // @[SRAM.scala 145:20:@50259.4]
  reg [31:0] _RAND_45;
  wire  _T_1093; // @[SRAM.scala 148:37:@50260.4]
  wire  _T_1094; // @[SRAM.scala 148:25:@50261.4]
  wire  _T_1095; // @[SRAM.scala 148:15:@50262.4]
  wire  _T_1096; // @[SRAM.scala 149:15:@50264.6]
  wire  _GEN_45; // @[SRAM.scala 148:48:@50263.4]
  reg  regs_46; // @[SRAM.scala 145:20:@50270.4]
  reg [31:0] _RAND_46;
  wire  _T_1102; // @[SRAM.scala 148:37:@50271.4]
  wire  _T_1103; // @[SRAM.scala 148:25:@50272.4]
  wire  _T_1104; // @[SRAM.scala 148:15:@50273.4]
  wire  _T_1105; // @[SRAM.scala 149:15:@50275.6]
  wire  _GEN_46; // @[SRAM.scala 148:48:@50274.4]
  reg  regs_47; // @[SRAM.scala 145:20:@50281.4]
  reg [31:0] _RAND_47;
  wire  _T_1111; // @[SRAM.scala 148:37:@50282.4]
  wire  _T_1112; // @[SRAM.scala 148:25:@50283.4]
  wire  _T_1113; // @[SRAM.scala 148:15:@50284.4]
  wire  _T_1114; // @[SRAM.scala 149:15:@50286.6]
  wire  _GEN_47; // @[SRAM.scala 148:48:@50285.4]
  reg  regs_48; // @[SRAM.scala 145:20:@50292.4]
  reg [31:0] _RAND_48;
  wire  _T_1120; // @[SRAM.scala 148:37:@50293.4]
  wire  _T_1121; // @[SRAM.scala 148:25:@50294.4]
  wire  _T_1122; // @[SRAM.scala 148:15:@50295.4]
  wire  _T_1123; // @[SRAM.scala 149:15:@50297.6]
  wire  _GEN_48; // @[SRAM.scala 148:48:@50296.4]
  reg  regs_49; // @[SRAM.scala 145:20:@50303.4]
  reg [31:0] _RAND_49;
  wire  _T_1129; // @[SRAM.scala 148:37:@50304.4]
  wire  _T_1130; // @[SRAM.scala 148:25:@50305.4]
  wire  _T_1131; // @[SRAM.scala 148:15:@50306.4]
  wire  _T_1132; // @[SRAM.scala 149:15:@50308.6]
  wire  _GEN_49; // @[SRAM.scala 148:48:@50307.4]
  reg  regs_50; // @[SRAM.scala 145:20:@50314.4]
  reg [31:0] _RAND_50;
  wire  _T_1138; // @[SRAM.scala 148:37:@50315.4]
  wire  _T_1139; // @[SRAM.scala 148:25:@50316.4]
  wire  _T_1140; // @[SRAM.scala 148:15:@50317.4]
  wire  _T_1141; // @[SRAM.scala 149:15:@50319.6]
  wire  _GEN_50; // @[SRAM.scala 148:48:@50318.4]
  reg  regs_51; // @[SRAM.scala 145:20:@50325.4]
  reg [31:0] _RAND_51;
  wire  _T_1147; // @[SRAM.scala 148:37:@50326.4]
  wire  _T_1148; // @[SRAM.scala 148:25:@50327.4]
  wire  _T_1149; // @[SRAM.scala 148:15:@50328.4]
  wire  _T_1150; // @[SRAM.scala 149:15:@50330.6]
  wire  _GEN_51; // @[SRAM.scala 148:48:@50329.4]
  reg  regs_52; // @[SRAM.scala 145:20:@50336.4]
  reg [31:0] _RAND_52;
  wire  _T_1156; // @[SRAM.scala 148:37:@50337.4]
  wire  _T_1157; // @[SRAM.scala 148:25:@50338.4]
  wire  _T_1158; // @[SRAM.scala 148:15:@50339.4]
  wire  _T_1159; // @[SRAM.scala 149:15:@50341.6]
  wire  _GEN_52; // @[SRAM.scala 148:48:@50340.4]
  reg  regs_53; // @[SRAM.scala 145:20:@50347.4]
  reg [31:0] _RAND_53;
  wire  _T_1165; // @[SRAM.scala 148:37:@50348.4]
  wire  _T_1166; // @[SRAM.scala 148:25:@50349.4]
  wire  _T_1167; // @[SRAM.scala 148:15:@50350.4]
  wire  _T_1168; // @[SRAM.scala 149:15:@50352.6]
  wire  _GEN_53; // @[SRAM.scala 148:48:@50351.4]
  reg  regs_54; // @[SRAM.scala 145:20:@50358.4]
  reg [31:0] _RAND_54;
  wire  _T_1174; // @[SRAM.scala 148:37:@50359.4]
  wire  _T_1175; // @[SRAM.scala 148:25:@50360.4]
  wire  _T_1176; // @[SRAM.scala 148:15:@50361.4]
  wire  _T_1177; // @[SRAM.scala 149:15:@50363.6]
  wire  _GEN_54; // @[SRAM.scala 148:48:@50362.4]
  reg  regs_55; // @[SRAM.scala 145:20:@50369.4]
  reg [31:0] _RAND_55;
  wire  _T_1183; // @[SRAM.scala 148:37:@50370.4]
  wire  _T_1184; // @[SRAM.scala 148:25:@50371.4]
  wire  _T_1185; // @[SRAM.scala 148:15:@50372.4]
  wire  _T_1186; // @[SRAM.scala 149:15:@50374.6]
  wire  _GEN_55; // @[SRAM.scala 148:48:@50373.4]
  reg  regs_56; // @[SRAM.scala 145:20:@50380.4]
  reg [31:0] _RAND_56;
  wire  _T_1192; // @[SRAM.scala 148:37:@50381.4]
  wire  _T_1193; // @[SRAM.scala 148:25:@50382.4]
  wire  _T_1194; // @[SRAM.scala 148:15:@50383.4]
  wire  _T_1195; // @[SRAM.scala 149:15:@50385.6]
  wire  _GEN_56; // @[SRAM.scala 148:48:@50384.4]
  reg  regs_57; // @[SRAM.scala 145:20:@50391.4]
  reg [31:0] _RAND_57;
  wire  _T_1201; // @[SRAM.scala 148:37:@50392.4]
  wire  _T_1202; // @[SRAM.scala 148:25:@50393.4]
  wire  _T_1203; // @[SRAM.scala 148:15:@50394.4]
  wire  _T_1204; // @[SRAM.scala 149:15:@50396.6]
  wire  _GEN_57; // @[SRAM.scala 148:48:@50395.4]
  reg  regs_58; // @[SRAM.scala 145:20:@50402.4]
  reg [31:0] _RAND_58;
  wire  _T_1210; // @[SRAM.scala 148:37:@50403.4]
  wire  _T_1211; // @[SRAM.scala 148:25:@50404.4]
  wire  _T_1212; // @[SRAM.scala 148:15:@50405.4]
  wire  _T_1213; // @[SRAM.scala 149:15:@50407.6]
  wire  _GEN_58; // @[SRAM.scala 148:48:@50406.4]
  reg  regs_59; // @[SRAM.scala 145:20:@50413.4]
  reg [31:0] _RAND_59;
  wire  _T_1219; // @[SRAM.scala 148:37:@50414.4]
  wire  _T_1220; // @[SRAM.scala 148:25:@50415.4]
  wire  _T_1221; // @[SRAM.scala 148:15:@50416.4]
  wire  _T_1222; // @[SRAM.scala 149:15:@50418.6]
  wire  _GEN_59; // @[SRAM.scala 148:48:@50417.4]
  reg  regs_60; // @[SRAM.scala 145:20:@50424.4]
  reg [31:0] _RAND_60;
  wire  _T_1228; // @[SRAM.scala 148:37:@50425.4]
  wire  _T_1229; // @[SRAM.scala 148:25:@50426.4]
  wire  _T_1230; // @[SRAM.scala 148:15:@50427.4]
  wire  _T_1231; // @[SRAM.scala 149:15:@50429.6]
  wire  _GEN_60; // @[SRAM.scala 148:48:@50428.4]
  reg  regs_61; // @[SRAM.scala 145:20:@50435.4]
  reg [31:0] _RAND_61;
  wire  _T_1237; // @[SRAM.scala 148:37:@50436.4]
  wire  _T_1238; // @[SRAM.scala 148:25:@50437.4]
  wire  _T_1239; // @[SRAM.scala 148:15:@50438.4]
  wire  _T_1240; // @[SRAM.scala 149:15:@50440.6]
  wire  _GEN_61; // @[SRAM.scala 148:48:@50439.4]
  reg  regs_62; // @[SRAM.scala 145:20:@50446.4]
  reg [31:0] _RAND_62;
  wire  _T_1246; // @[SRAM.scala 148:37:@50447.4]
  wire  _T_1247; // @[SRAM.scala 148:25:@50448.4]
  wire  _T_1248; // @[SRAM.scala 148:15:@50449.4]
  wire  _T_1249; // @[SRAM.scala 149:15:@50451.6]
  wire  _GEN_62; // @[SRAM.scala 148:48:@50450.4]
  reg  regs_63; // @[SRAM.scala 145:20:@50457.4]
  reg [31:0] _RAND_63;
  wire  _T_1255; // @[SRAM.scala 148:37:@50458.4]
  wire  _T_1256; // @[SRAM.scala 148:25:@50459.4]
  wire  _T_1257; // @[SRAM.scala 148:15:@50460.4]
  wire  _T_1258; // @[SRAM.scala 149:15:@50462.6]
  wire  _GEN_63; // @[SRAM.scala 148:48:@50461.4]
  wire  _GEN_65; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_66; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_67; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_68; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_69; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_70; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_71; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_72; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_73; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_74; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_75; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_76; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_77; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_78; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_79; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_80; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_81; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_82; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_83; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_84; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_85; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_86; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_87; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_88; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_89; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_90; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_91; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_92; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_93; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_94; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_95; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_96; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_97; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_98; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_99; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_100; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_101; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_102; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_103; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_104; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_105; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_106; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_107; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_108; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_109; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_110; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_111; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_112; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_113; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_114; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_115; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_116; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_117; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_118; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_119; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_120; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_121; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_122; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_123; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_124; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_125; // @[SRAM.scala 155:12:@50531.4]
  wire  _GEN_126; // @[SRAM.scala 155:12:@50531.4]
  assign _T_688 = io_waddr == 6'h0; // @[SRAM.scala 148:37:@49765.4]
  assign _T_689 = io_wen & _T_688; // @[SRAM.scala 148:25:@49766.4]
  assign _T_690 = io_banks_0_wdata_valid | _T_689; // @[SRAM.scala 148:15:@49767.4]
  assign _T_691 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49769.6]
  assign _GEN_0 = _T_690 ? _T_691 : regs_0; // @[SRAM.scala 148:48:@49768.4]
  assign _T_697 = io_waddr == 6'h1; // @[SRAM.scala 148:37:@49776.4]
  assign _T_698 = io_wen & _T_697; // @[SRAM.scala 148:25:@49777.4]
  assign _T_699 = io_banks_1_wdata_valid | _T_698; // @[SRAM.scala 148:15:@49778.4]
  assign _T_700 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49780.6]
  assign _GEN_1 = _T_699 ? _T_700 : regs_1; // @[SRAM.scala 148:48:@49779.4]
  assign _T_706 = io_waddr == 6'h2; // @[SRAM.scala 148:37:@49787.4]
  assign _T_707 = io_wen & _T_706; // @[SRAM.scala 148:25:@49788.4]
  assign _T_708 = io_banks_2_wdata_valid | _T_707; // @[SRAM.scala 148:15:@49789.4]
  assign _T_709 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49791.6]
  assign _GEN_2 = _T_708 ? _T_709 : regs_2; // @[SRAM.scala 148:48:@49790.4]
  assign _T_715 = io_waddr == 6'h3; // @[SRAM.scala 148:37:@49798.4]
  assign _T_716 = io_wen & _T_715; // @[SRAM.scala 148:25:@49799.4]
  assign _T_717 = io_banks_3_wdata_valid | _T_716; // @[SRAM.scala 148:15:@49800.4]
  assign _T_718 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49802.6]
  assign _GEN_3 = _T_717 ? _T_718 : regs_3; // @[SRAM.scala 148:48:@49801.4]
  assign _T_724 = io_waddr == 6'h4; // @[SRAM.scala 148:37:@49809.4]
  assign _T_725 = io_wen & _T_724; // @[SRAM.scala 148:25:@49810.4]
  assign _T_726 = io_banks_4_wdata_valid | _T_725; // @[SRAM.scala 148:15:@49811.4]
  assign _T_727 = io_banks_4_wdata_valid ? io_banks_4_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49813.6]
  assign _GEN_4 = _T_726 ? _T_727 : regs_4; // @[SRAM.scala 148:48:@49812.4]
  assign _T_733 = io_waddr == 6'h5; // @[SRAM.scala 148:37:@49820.4]
  assign _T_734 = io_wen & _T_733; // @[SRAM.scala 148:25:@49821.4]
  assign _T_735 = io_banks_5_wdata_valid | _T_734; // @[SRAM.scala 148:15:@49822.4]
  assign _T_736 = io_banks_5_wdata_valid ? io_banks_5_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49824.6]
  assign _GEN_5 = _T_735 ? _T_736 : regs_5; // @[SRAM.scala 148:48:@49823.4]
  assign _T_742 = io_waddr == 6'h6; // @[SRAM.scala 148:37:@49831.4]
  assign _T_743 = io_wen & _T_742; // @[SRAM.scala 148:25:@49832.4]
  assign _T_744 = io_banks_6_wdata_valid | _T_743; // @[SRAM.scala 148:15:@49833.4]
  assign _T_745 = io_banks_6_wdata_valid ? io_banks_6_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49835.6]
  assign _GEN_6 = _T_744 ? _T_745 : regs_6; // @[SRAM.scala 148:48:@49834.4]
  assign _T_751 = io_waddr == 6'h7; // @[SRAM.scala 148:37:@49842.4]
  assign _T_752 = io_wen & _T_751; // @[SRAM.scala 148:25:@49843.4]
  assign _T_753 = io_banks_7_wdata_valid | _T_752; // @[SRAM.scala 148:15:@49844.4]
  assign _T_754 = io_banks_7_wdata_valid ? io_banks_7_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49846.6]
  assign _GEN_7 = _T_753 ? _T_754 : regs_7; // @[SRAM.scala 148:48:@49845.4]
  assign _T_760 = io_waddr == 6'h8; // @[SRAM.scala 148:37:@49853.4]
  assign _T_761 = io_wen & _T_760; // @[SRAM.scala 148:25:@49854.4]
  assign _T_762 = io_banks_8_wdata_valid | _T_761; // @[SRAM.scala 148:15:@49855.4]
  assign _T_763 = io_banks_8_wdata_valid ? io_banks_8_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49857.6]
  assign _GEN_8 = _T_762 ? _T_763 : regs_8; // @[SRAM.scala 148:48:@49856.4]
  assign _T_769 = io_waddr == 6'h9; // @[SRAM.scala 148:37:@49864.4]
  assign _T_770 = io_wen & _T_769; // @[SRAM.scala 148:25:@49865.4]
  assign _T_771 = io_banks_9_wdata_valid | _T_770; // @[SRAM.scala 148:15:@49866.4]
  assign _T_772 = io_banks_9_wdata_valid ? io_banks_9_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49868.6]
  assign _GEN_9 = _T_771 ? _T_772 : regs_9; // @[SRAM.scala 148:48:@49867.4]
  assign _T_778 = io_waddr == 6'ha; // @[SRAM.scala 148:37:@49875.4]
  assign _T_779 = io_wen & _T_778; // @[SRAM.scala 148:25:@49876.4]
  assign _T_780 = io_banks_10_wdata_valid | _T_779; // @[SRAM.scala 148:15:@49877.4]
  assign _T_781 = io_banks_10_wdata_valid ? io_banks_10_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49879.6]
  assign _GEN_10 = _T_780 ? _T_781 : regs_10; // @[SRAM.scala 148:48:@49878.4]
  assign _T_787 = io_waddr == 6'hb; // @[SRAM.scala 148:37:@49886.4]
  assign _T_788 = io_wen & _T_787; // @[SRAM.scala 148:25:@49887.4]
  assign _T_789 = io_banks_11_wdata_valid | _T_788; // @[SRAM.scala 148:15:@49888.4]
  assign _T_790 = io_banks_11_wdata_valid ? io_banks_11_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49890.6]
  assign _GEN_11 = _T_789 ? _T_790 : regs_11; // @[SRAM.scala 148:48:@49889.4]
  assign _T_796 = io_waddr == 6'hc; // @[SRAM.scala 148:37:@49897.4]
  assign _T_797 = io_wen & _T_796; // @[SRAM.scala 148:25:@49898.4]
  assign _T_798 = io_banks_12_wdata_valid | _T_797; // @[SRAM.scala 148:15:@49899.4]
  assign _T_799 = io_banks_12_wdata_valid ? io_banks_12_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49901.6]
  assign _GEN_12 = _T_798 ? _T_799 : regs_12; // @[SRAM.scala 148:48:@49900.4]
  assign _T_805 = io_waddr == 6'hd; // @[SRAM.scala 148:37:@49908.4]
  assign _T_806 = io_wen & _T_805; // @[SRAM.scala 148:25:@49909.4]
  assign _T_807 = io_banks_13_wdata_valid | _T_806; // @[SRAM.scala 148:15:@49910.4]
  assign _T_808 = io_banks_13_wdata_valid ? io_banks_13_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49912.6]
  assign _GEN_13 = _T_807 ? _T_808 : regs_13; // @[SRAM.scala 148:48:@49911.4]
  assign _T_814 = io_waddr == 6'he; // @[SRAM.scala 148:37:@49919.4]
  assign _T_815 = io_wen & _T_814; // @[SRAM.scala 148:25:@49920.4]
  assign _T_816 = io_banks_14_wdata_valid | _T_815; // @[SRAM.scala 148:15:@49921.4]
  assign _T_817 = io_banks_14_wdata_valid ? io_banks_14_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49923.6]
  assign _GEN_14 = _T_816 ? _T_817 : regs_14; // @[SRAM.scala 148:48:@49922.4]
  assign _T_823 = io_waddr == 6'hf; // @[SRAM.scala 148:37:@49930.4]
  assign _T_824 = io_wen & _T_823; // @[SRAM.scala 148:25:@49931.4]
  assign _T_825 = io_banks_15_wdata_valid | _T_824; // @[SRAM.scala 148:15:@49932.4]
  assign _T_826 = io_banks_15_wdata_valid ? io_banks_15_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49934.6]
  assign _GEN_15 = _T_825 ? _T_826 : regs_15; // @[SRAM.scala 148:48:@49933.4]
  assign _T_832 = io_waddr == 6'h10; // @[SRAM.scala 148:37:@49941.4]
  assign _T_833 = io_wen & _T_832; // @[SRAM.scala 148:25:@49942.4]
  assign _T_834 = io_banks_16_wdata_valid | _T_833; // @[SRAM.scala 148:15:@49943.4]
  assign _T_835 = io_banks_16_wdata_valid ? io_banks_16_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49945.6]
  assign _GEN_16 = _T_834 ? _T_835 : regs_16; // @[SRAM.scala 148:48:@49944.4]
  assign _T_841 = io_waddr == 6'h11; // @[SRAM.scala 148:37:@49952.4]
  assign _T_842 = io_wen & _T_841; // @[SRAM.scala 148:25:@49953.4]
  assign _T_843 = io_banks_17_wdata_valid | _T_842; // @[SRAM.scala 148:15:@49954.4]
  assign _T_844 = io_banks_17_wdata_valid ? io_banks_17_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49956.6]
  assign _GEN_17 = _T_843 ? _T_844 : regs_17; // @[SRAM.scala 148:48:@49955.4]
  assign _T_850 = io_waddr == 6'h12; // @[SRAM.scala 148:37:@49963.4]
  assign _T_851 = io_wen & _T_850; // @[SRAM.scala 148:25:@49964.4]
  assign _T_852 = io_banks_18_wdata_valid | _T_851; // @[SRAM.scala 148:15:@49965.4]
  assign _T_853 = io_banks_18_wdata_valid ? io_banks_18_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49967.6]
  assign _GEN_18 = _T_852 ? _T_853 : regs_18; // @[SRAM.scala 148:48:@49966.4]
  assign _T_859 = io_waddr == 6'h13; // @[SRAM.scala 148:37:@49974.4]
  assign _T_860 = io_wen & _T_859; // @[SRAM.scala 148:25:@49975.4]
  assign _T_861 = io_banks_19_wdata_valid | _T_860; // @[SRAM.scala 148:15:@49976.4]
  assign _T_862 = io_banks_19_wdata_valid ? io_banks_19_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49978.6]
  assign _GEN_19 = _T_861 ? _T_862 : regs_19; // @[SRAM.scala 148:48:@49977.4]
  assign _T_868 = io_waddr == 6'h14; // @[SRAM.scala 148:37:@49985.4]
  assign _T_869 = io_wen & _T_868; // @[SRAM.scala 148:25:@49986.4]
  assign _T_870 = io_banks_20_wdata_valid | _T_869; // @[SRAM.scala 148:15:@49987.4]
  assign _T_871 = io_banks_20_wdata_valid ? io_banks_20_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49989.6]
  assign _GEN_20 = _T_870 ? _T_871 : regs_20; // @[SRAM.scala 148:48:@49988.4]
  assign _T_877 = io_waddr == 6'h15; // @[SRAM.scala 148:37:@49996.4]
  assign _T_878 = io_wen & _T_877; // @[SRAM.scala 148:25:@49997.4]
  assign _T_879 = io_banks_21_wdata_valid | _T_878; // @[SRAM.scala 148:15:@49998.4]
  assign _T_880 = io_banks_21_wdata_valid ? io_banks_21_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50000.6]
  assign _GEN_21 = _T_879 ? _T_880 : regs_21; // @[SRAM.scala 148:48:@49999.4]
  assign _T_886 = io_waddr == 6'h16; // @[SRAM.scala 148:37:@50007.4]
  assign _T_887 = io_wen & _T_886; // @[SRAM.scala 148:25:@50008.4]
  assign _T_888 = io_banks_22_wdata_valid | _T_887; // @[SRAM.scala 148:15:@50009.4]
  assign _T_889 = io_banks_22_wdata_valid ? io_banks_22_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50011.6]
  assign _GEN_22 = _T_888 ? _T_889 : regs_22; // @[SRAM.scala 148:48:@50010.4]
  assign _T_895 = io_waddr == 6'h17; // @[SRAM.scala 148:37:@50018.4]
  assign _T_896 = io_wen & _T_895; // @[SRAM.scala 148:25:@50019.4]
  assign _T_897 = io_banks_23_wdata_valid | _T_896; // @[SRAM.scala 148:15:@50020.4]
  assign _T_898 = io_banks_23_wdata_valid ? io_banks_23_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50022.6]
  assign _GEN_23 = _T_897 ? _T_898 : regs_23; // @[SRAM.scala 148:48:@50021.4]
  assign _T_904 = io_waddr == 6'h18; // @[SRAM.scala 148:37:@50029.4]
  assign _T_905 = io_wen & _T_904; // @[SRAM.scala 148:25:@50030.4]
  assign _T_906 = io_banks_24_wdata_valid | _T_905; // @[SRAM.scala 148:15:@50031.4]
  assign _T_907 = io_banks_24_wdata_valid ? io_banks_24_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50033.6]
  assign _GEN_24 = _T_906 ? _T_907 : regs_24; // @[SRAM.scala 148:48:@50032.4]
  assign _T_913 = io_waddr == 6'h19; // @[SRAM.scala 148:37:@50040.4]
  assign _T_914 = io_wen & _T_913; // @[SRAM.scala 148:25:@50041.4]
  assign _T_915 = io_banks_25_wdata_valid | _T_914; // @[SRAM.scala 148:15:@50042.4]
  assign _T_916 = io_banks_25_wdata_valid ? io_banks_25_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50044.6]
  assign _GEN_25 = _T_915 ? _T_916 : regs_25; // @[SRAM.scala 148:48:@50043.4]
  assign _T_922 = io_waddr == 6'h1a; // @[SRAM.scala 148:37:@50051.4]
  assign _T_923 = io_wen & _T_922; // @[SRAM.scala 148:25:@50052.4]
  assign _T_924 = io_banks_26_wdata_valid | _T_923; // @[SRAM.scala 148:15:@50053.4]
  assign _T_925 = io_banks_26_wdata_valid ? io_banks_26_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50055.6]
  assign _GEN_26 = _T_924 ? _T_925 : regs_26; // @[SRAM.scala 148:48:@50054.4]
  assign _T_931 = io_waddr == 6'h1b; // @[SRAM.scala 148:37:@50062.4]
  assign _T_932 = io_wen & _T_931; // @[SRAM.scala 148:25:@50063.4]
  assign _T_933 = io_banks_27_wdata_valid | _T_932; // @[SRAM.scala 148:15:@50064.4]
  assign _T_934 = io_banks_27_wdata_valid ? io_banks_27_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50066.6]
  assign _GEN_27 = _T_933 ? _T_934 : regs_27; // @[SRAM.scala 148:48:@50065.4]
  assign _T_940 = io_waddr == 6'h1c; // @[SRAM.scala 148:37:@50073.4]
  assign _T_941 = io_wen & _T_940; // @[SRAM.scala 148:25:@50074.4]
  assign _T_942 = io_banks_28_wdata_valid | _T_941; // @[SRAM.scala 148:15:@50075.4]
  assign _T_943 = io_banks_28_wdata_valid ? io_banks_28_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50077.6]
  assign _GEN_28 = _T_942 ? _T_943 : regs_28; // @[SRAM.scala 148:48:@50076.4]
  assign _T_949 = io_waddr == 6'h1d; // @[SRAM.scala 148:37:@50084.4]
  assign _T_950 = io_wen & _T_949; // @[SRAM.scala 148:25:@50085.4]
  assign _T_951 = io_banks_29_wdata_valid | _T_950; // @[SRAM.scala 148:15:@50086.4]
  assign _T_952 = io_banks_29_wdata_valid ? io_banks_29_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50088.6]
  assign _GEN_29 = _T_951 ? _T_952 : regs_29; // @[SRAM.scala 148:48:@50087.4]
  assign _T_958 = io_waddr == 6'h1e; // @[SRAM.scala 148:37:@50095.4]
  assign _T_959 = io_wen & _T_958; // @[SRAM.scala 148:25:@50096.4]
  assign _T_960 = io_banks_30_wdata_valid | _T_959; // @[SRAM.scala 148:15:@50097.4]
  assign _T_961 = io_banks_30_wdata_valid ? io_banks_30_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50099.6]
  assign _GEN_30 = _T_960 ? _T_961 : regs_30; // @[SRAM.scala 148:48:@50098.4]
  assign _T_967 = io_waddr == 6'h1f; // @[SRAM.scala 148:37:@50106.4]
  assign _T_968 = io_wen & _T_967; // @[SRAM.scala 148:25:@50107.4]
  assign _T_969 = io_banks_31_wdata_valid | _T_968; // @[SRAM.scala 148:15:@50108.4]
  assign _T_970 = io_banks_31_wdata_valid ? io_banks_31_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50110.6]
  assign _GEN_31 = _T_969 ? _T_970 : regs_31; // @[SRAM.scala 148:48:@50109.4]
  assign _T_976 = io_waddr == 6'h20; // @[SRAM.scala 148:37:@50117.4]
  assign _T_977 = io_wen & _T_976; // @[SRAM.scala 148:25:@50118.4]
  assign _T_978 = io_banks_32_wdata_valid | _T_977; // @[SRAM.scala 148:15:@50119.4]
  assign _T_979 = io_banks_32_wdata_valid ? io_banks_32_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50121.6]
  assign _GEN_32 = _T_978 ? _T_979 : regs_32; // @[SRAM.scala 148:48:@50120.4]
  assign _T_985 = io_waddr == 6'h21; // @[SRAM.scala 148:37:@50128.4]
  assign _T_986 = io_wen & _T_985; // @[SRAM.scala 148:25:@50129.4]
  assign _T_987 = io_banks_33_wdata_valid | _T_986; // @[SRAM.scala 148:15:@50130.4]
  assign _T_988 = io_banks_33_wdata_valid ? io_banks_33_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50132.6]
  assign _GEN_33 = _T_987 ? _T_988 : regs_33; // @[SRAM.scala 148:48:@50131.4]
  assign _T_994 = io_waddr == 6'h22; // @[SRAM.scala 148:37:@50139.4]
  assign _T_995 = io_wen & _T_994; // @[SRAM.scala 148:25:@50140.4]
  assign _T_996 = io_banks_34_wdata_valid | _T_995; // @[SRAM.scala 148:15:@50141.4]
  assign _T_997 = io_banks_34_wdata_valid ? io_banks_34_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50143.6]
  assign _GEN_34 = _T_996 ? _T_997 : regs_34; // @[SRAM.scala 148:48:@50142.4]
  assign _T_1003 = io_waddr == 6'h23; // @[SRAM.scala 148:37:@50150.4]
  assign _T_1004 = io_wen & _T_1003; // @[SRAM.scala 148:25:@50151.4]
  assign _T_1005 = io_banks_35_wdata_valid | _T_1004; // @[SRAM.scala 148:15:@50152.4]
  assign _T_1006 = io_banks_35_wdata_valid ? io_banks_35_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50154.6]
  assign _GEN_35 = _T_1005 ? _T_1006 : regs_35; // @[SRAM.scala 148:48:@50153.4]
  assign _T_1012 = io_waddr == 6'h24; // @[SRAM.scala 148:37:@50161.4]
  assign _T_1013 = io_wen & _T_1012; // @[SRAM.scala 148:25:@50162.4]
  assign _T_1014 = io_banks_36_wdata_valid | _T_1013; // @[SRAM.scala 148:15:@50163.4]
  assign _T_1015 = io_banks_36_wdata_valid ? io_banks_36_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50165.6]
  assign _GEN_36 = _T_1014 ? _T_1015 : regs_36; // @[SRAM.scala 148:48:@50164.4]
  assign _T_1021 = io_waddr == 6'h25; // @[SRAM.scala 148:37:@50172.4]
  assign _T_1022 = io_wen & _T_1021; // @[SRAM.scala 148:25:@50173.4]
  assign _T_1023 = io_banks_37_wdata_valid | _T_1022; // @[SRAM.scala 148:15:@50174.4]
  assign _T_1024 = io_banks_37_wdata_valid ? io_banks_37_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50176.6]
  assign _GEN_37 = _T_1023 ? _T_1024 : regs_37; // @[SRAM.scala 148:48:@50175.4]
  assign _T_1030 = io_waddr == 6'h26; // @[SRAM.scala 148:37:@50183.4]
  assign _T_1031 = io_wen & _T_1030; // @[SRAM.scala 148:25:@50184.4]
  assign _T_1032 = io_banks_38_wdata_valid | _T_1031; // @[SRAM.scala 148:15:@50185.4]
  assign _T_1033 = io_banks_38_wdata_valid ? io_banks_38_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50187.6]
  assign _GEN_38 = _T_1032 ? _T_1033 : regs_38; // @[SRAM.scala 148:48:@50186.4]
  assign _T_1039 = io_waddr == 6'h27; // @[SRAM.scala 148:37:@50194.4]
  assign _T_1040 = io_wen & _T_1039; // @[SRAM.scala 148:25:@50195.4]
  assign _T_1041 = io_banks_39_wdata_valid | _T_1040; // @[SRAM.scala 148:15:@50196.4]
  assign _T_1042 = io_banks_39_wdata_valid ? io_banks_39_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50198.6]
  assign _GEN_39 = _T_1041 ? _T_1042 : regs_39; // @[SRAM.scala 148:48:@50197.4]
  assign _T_1048 = io_waddr == 6'h28; // @[SRAM.scala 148:37:@50205.4]
  assign _T_1049 = io_wen & _T_1048; // @[SRAM.scala 148:25:@50206.4]
  assign _T_1050 = io_banks_40_wdata_valid | _T_1049; // @[SRAM.scala 148:15:@50207.4]
  assign _T_1051 = io_banks_40_wdata_valid ? io_banks_40_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50209.6]
  assign _GEN_40 = _T_1050 ? _T_1051 : regs_40; // @[SRAM.scala 148:48:@50208.4]
  assign _T_1057 = io_waddr == 6'h29; // @[SRAM.scala 148:37:@50216.4]
  assign _T_1058 = io_wen & _T_1057; // @[SRAM.scala 148:25:@50217.4]
  assign _T_1059 = io_banks_41_wdata_valid | _T_1058; // @[SRAM.scala 148:15:@50218.4]
  assign _T_1060 = io_banks_41_wdata_valid ? io_banks_41_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50220.6]
  assign _GEN_41 = _T_1059 ? _T_1060 : regs_41; // @[SRAM.scala 148:48:@50219.4]
  assign _T_1066 = io_waddr == 6'h2a; // @[SRAM.scala 148:37:@50227.4]
  assign _T_1067 = io_wen & _T_1066; // @[SRAM.scala 148:25:@50228.4]
  assign _T_1068 = io_banks_42_wdata_valid | _T_1067; // @[SRAM.scala 148:15:@50229.4]
  assign _T_1069 = io_banks_42_wdata_valid ? io_banks_42_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50231.6]
  assign _GEN_42 = _T_1068 ? _T_1069 : regs_42; // @[SRAM.scala 148:48:@50230.4]
  assign _T_1075 = io_waddr == 6'h2b; // @[SRAM.scala 148:37:@50238.4]
  assign _T_1076 = io_wen & _T_1075; // @[SRAM.scala 148:25:@50239.4]
  assign _T_1077 = io_banks_43_wdata_valid | _T_1076; // @[SRAM.scala 148:15:@50240.4]
  assign _T_1078 = io_banks_43_wdata_valid ? io_banks_43_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50242.6]
  assign _GEN_43 = _T_1077 ? _T_1078 : regs_43; // @[SRAM.scala 148:48:@50241.4]
  assign _T_1084 = io_waddr == 6'h2c; // @[SRAM.scala 148:37:@50249.4]
  assign _T_1085 = io_wen & _T_1084; // @[SRAM.scala 148:25:@50250.4]
  assign _T_1086 = io_banks_44_wdata_valid | _T_1085; // @[SRAM.scala 148:15:@50251.4]
  assign _T_1087 = io_banks_44_wdata_valid ? io_banks_44_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50253.6]
  assign _GEN_44 = _T_1086 ? _T_1087 : regs_44; // @[SRAM.scala 148:48:@50252.4]
  assign _T_1093 = io_waddr == 6'h2d; // @[SRAM.scala 148:37:@50260.4]
  assign _T_1094 = io_wen & _T_1093; // @[SRAM.scala 148:25:@50261.4]
  assign _T_1095 = io_banks_45_wdata_valid | _T_1094; // @[SRAM.scala 148:15:@50262.4]
  assign _T_1096 = io_banks_45_wdata_valid ? io_banks_45_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50264.6]
  assign _GEN_45 = _T_1095 ? _T_1096 : regs_45; // @[SRAM.scala 148:48:@50263.4]
  assign _T_1102 = io_waddr == 6'h2e; // @[SRAM.scala 148:37:@50271.4]
  assign _T_1103 = io_wen & _T_1102; // @[SRAM.scala 148:25:@50272.4]
  assign _T_1104 = io_banks_46_wdata_valid | _T_1103; // @[SRAM.scala 148:15:@50273.4]
  assign _T_1105 = io_banks_46_wdata_valid ? io_banks_46_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50275.6]
  assign _GEN_46 = _T_1104 ? _T_1105 : regs_46; // @[SRAM.scala 148:48:@50274.4]
  assign _T_1111 = io_waddr == 6'h2f; // @[SRAM.scala 148:37:@50282.4]
  assign _T_1112 = io_wen & _T_1111; // @[SRAM.scala 148:25:@50283.4]
  assign _T_1113 = io_banks_47_wdata_valid | _T_1112; // @[SRAM.scala 148:15:@50284.4]
  assign _T_1114 = io_banks_47_wdata_valid ? io_banks_47_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50286.6]
  assign _GEN_47 = _T_1113 ? _T_1114 : regs_47; // @[SRAM.scala 148:48:@50285.4]
  assign _T_1120 = io_waddr == 6'h30; // @[SRAM.scala 148:37:@50293.4]
  assign _T_1121 = io_wen & _T_1120; // @[SRAM.scala 148:25:@50294.4]
  assign _T_1122 = io_banks_48_wdata_valid | _T_1121; // @[SRAM.scala 148:15:@50295.4]
  assign _T_1123 = io_banks_48_wdata_valid ? io_banks_48_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50297.6]
  assign _GEN_48 = _T_1122 ? _T_1123 : regs_48; // @[SRAM.scala 148:48:@50296.4]
  assign _T_1129 = io_waddr == 6'h31; // @[SRAM.scala 148:37:@50304.4]
  assign _T_1130 = io_wen & _T_1129; // @[SRAM.scala 148:25:@50305.4]
  assign _T_1131 = io_banks_49_wdata_valid | _T_1130; // @[SRAM.scala 148:15:@50306.4]
  assign _T_1132 = io_banks_49_wdata_valid ? io_banks_49_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50308.6]
  assign _GEN_49 = _T_1131 ? _T_1132 : regs_49; // @[SRAM.scala 148:48:@50307.4]
  assign _T_1138 = io_waddr == 6'h32; // @[SRAM.scala 148:37:@50315.4]
  assign _T_1139 = io_wen & _T_1138; // @[SRAM.scala 148:25:@50316.4]
  assign _T_1140 = io_banks_50_wdata_valid | _T_1139; // @[SRAM.scala 148:15:@50317.4]
  assign _T_1141 = io_banks_50_wdata_valid ? io_banks_50_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50319.6]
  assign _GEN_50 = _T_1140 ? _T_1141 : regs_50; // @[SRAM.scala 148:48:@50318.4]
  assign _T_1147 = io_waddr == 6'h33; // @[SRAM.scala 148:37:@50326.4]
  assign _T_1148 = io_wen & _T_1147; // @[SRAM.scala 148:25:@50327.4]
  assign _T_1149 = io_banks_51_wdata_valid | _T_1148; // @[SRAM.scala 148:15:@50328.4]
  assign _T_1150 = io_banks_51_wdata_valid ? io_banks_51_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50330.6]
  assign _GEN_51 = _T_1149 ? _T_1150 : regs_51; // @[SRAM.scala 148:48:@50329.4]
  assign _T_1156 = io_waddr == 6'h34; // @[SRAM.scala 148:37:@50337.4]
  assign _T_1157 = io_wen & _T_1156; // @[SRAM.scala 148:25:@50338.4]
  assign _T_1158 = io_banks_52_wdata_valid | _T_1157; // @[SRAM.scala 148:15:@50339.4]
  assign _T_1159 = io_banks_52_wdata_valid ? io_banks_52_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50341.6]
  assign _GEN_52 = _T_1158 ? _T_1159 : regs_52; // @[SRAM.scala 148:48:@50340.4]
  assign _T_1165 = io_waddr == 6'h35; // @[SRAM.scala 148:37:@50348.4]
  assign _T_1166 = io_wen & _T_1165; // @[SRAM.scala 148:25:@50349.4]
  assign _T_1167 = io_banks_53_wdata_valid | _T_1166; // @[SRAM.scala 148:15:@50350.4]
  assign _T_1168 = io_banks_53_wdata_valid ? io_banks_53_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50352.6]
  assign _GEN_53 = _T_1167 ? _T_1168 : regs_53; // @[SRAM.scala 148:48:@50351.4]
  assign _T_1174 = io_waddr == 6'h36; // @[SRAM.scala 148:37:@50359.4]
  assign _T_1175 = io_wen & _T_1174; // @[SRAM.scala 148:25:@50360.4]
  assign _T_1176 = io_banks_54_wdata_valid | _T_1175; // @[SRAM.scala 148:15:@50361.4]
  assign _T_1177 = io_banks_54_wdata_valid ? io_banks_54_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50363.6]
  assign _GEN_54 = _T_1176 ? _T_1177 : regs_54; // @[SRAM.scala 148:48:@50362.4]
  assign _T_1183 = io_waddr == 6'h37; // @[SRAM.scala 148:37:@50370.4]
  assign _T_1184 = io_wen & _T_1183; // @[SRAM.scala 148:25:@50371.4]
  assign _T_1185 = io_banks_55_wdata_valid | _T_1184; // @[SRAM.scala 148:15:@50372.4]
  assign _T_1186 = io_banks_55_wdata_valid ? io_banks_55_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50374.6]
  assign _GEN_55 = _T_1185 ? _T_1186 : regs_55; // @[SRAM.scala 148:48:@50373.4]
  assign _T_1192 = io_waddr == 6'h38; // @[SRAM.scala 148:37:@50381.4]
  assign _T_1193 = io_wen & _T_1192; // @[SRAM.scala 148:25:@50382.4]
  assign _T_1194 = io_banks_56_wdata_valid | _T_1193; // @[SRAM.scala 148:15:@50383.4]
  assign _T_1195 = io_banks_56_wdata_valid ? io_banks_56_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50385.6]
  assign _GEN_56 = _T_1194 ? _T_1195 : regs_56; // @[SRAM.scala 148:48:@50384.4]
  assign _T_1201 = io_waddr == 6'h39; // @[SRAM.scala 148:37:@50392.4]
  assign _T_1202 = io_wen & _T_1201; // @[SRAM.scala 148:25:@50393.4]
  assign _T_1203 = io_banks_57_wdata_valid | _T_1202; // @[SRAM.scala 148:15:@50394.4]
  assign _T_1204 = io_banks_57_wdata_valid ? io_banks_57_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50396.6]
  assign _GEN_57 = _T_1203 ? _T_1204 : regs_57; // @[SRAM.scala 148:48:@50395.4]
  assign _T_1210 = io_waddr == 6'h3a; // @[SRAM.scala 148:37:@50403.4]
  assign _T_1211 = io_wen & _T_1210; // @[SRAM.scala 148:25:@50404.4]
  assign _T_1212 = io_banks_58_wdata_valid | _T_1211; // @[SRAM.scala 148:15:@50405.4]
  assign _T_1213 = io_banks_58_wdata_valid ? io_banks_58_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50407.6]
  assign _GEN_58 = _T_1212 ? _T_1213 : regs_58; // @[SRAM.scala 148:48:@50406.4]
  assign _T_1219 = io_waddr == 6'h3b; // @[SRAM.scala 148:37:@50414.4]
  assign _T_1220 = io_wen & _T_1219; // @[SRAM.scala 148:25:@50415.4]
  assign _T_1221 = io_banks_59_wdata_valid | _T_1220; // @[SRAM.scala 148:15:@50416.4]
  assign _T_1222 = io_banks_59_wdata_valid ? io_banks_59_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50418.6]
  assign _GEN_59 = _T_1221 ? _T_1222 : regs_59; // @[SRAM.scala 148:48:@50417.4]
  assign _T_1228 = io_waddr == 6'h3c; // @[SRAM.scala 148:37:@50425.4]
  assign _T_1229 = io_wen & _T_1228; // @[SRAM.scala 148:25:@50426.4]
  assign _T_1230 = io_banks_60_wdata_valid | _T_1229; // @[SRAM.scala 148:15:@50427.4]
  assign _T_1231 = io_banks_60_wdata_valid ? io_banks_60_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50429.6]
  assign _GEN_60 = _T_1230 ? _T_1231 : regs_60; // @[SRAM.scala 148:48:@50428.4]
  assign _T_1237 = io_waddr == 6'h3d; // @[SRAM.scala 148:37:@50436.4]
  assign _T_1238 = io_wen & _T_1237; // @[SRAM.scala 148:25:@50437.4]
  assign _T_1239 = io_banks_61_wdata_valid | _T_1238; // @[SRAM.scala 148:15:@50438.4]
  assign _T_1240 = io_banks_61_wdata_valid ? io_banks_61_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50440.6]
  assign _GEN_61 = _T_1239 ? _T_1240 : regs_61; // @[SRAM.scala 148:48:@50439.4]
  assign _T_1246 = io_waddr == 6'h3e; // @[SRAM.scala 148:37:@50447.4]
  assign _T_1247 = io_wen & _T_1246; // @[SRAM.scala 148:25:@50448.4]
  assign _T_1248 = io_banks_62_wdata_valid | _T_1247; // @[SRAM.scala 148:15:@50449.4]
  assign _T_1249 = io_banks_62_wdata_valid ? io_banks_62_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50451.6]
  assign _GEN_62 = _T_1248 ? _T_1249 : regs_62; // @[SRAM.scala 148:48:@50450.4]
  assign _T_1255 = io_waddr == 6'h3f; // @[SRAM.scala 148:37:@50458.4]
  assign _T_1256 = io_wen & _T_1255; // @[SRAM.scala 148:25:@50459.4]
  assign _T_1257 = io_banks_63_wdata_valid | _T_1256; // @[SRAM.scala 148:15:@50460.4]
  assign _T_1258 = io_banks_63_wdata_valid ? io_banks_63_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50462.6]
  assign _GEN_63 = _T_1257 ? _T_1258 : regs_63; // @[SRAM.scala 148:48:@50461.4]
  assign _GEN_65 = 6'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_66 = 6'h2 == io_raddr ? regs_2 : _GEN_65; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_67 = 6'h3 == io_raddr ? regs_3 : _GEN_66; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_68 = 6'h4 == io_raddr ? regs_4 : _GEN_67; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_69 = 6'h5 == io_raddr ? regs_5 : _GEN_68; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_70 = 6'h6 == io_raddr ? regs_6 : _GEN_69; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_71 = 6'h7 == io_raddr ? regs_7 : _GEN_70; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_72 = 6'h8 == io_raddr ? regs_8 : _GEN_71; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_73 = 6'h9 == io_raddr ? regs_9 : _GEN_72; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_74 = 6'ha == io_raddr ? regs_10 : _GEN_73; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_75 = 6'hb == io_raddr ? regs_11 : _GEN_74; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_76 = 6'hc == io_raddr ? regs_12 : _GEN_75; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_77 = 6'hd == io_raddr ? regs_13 : _GEN_76; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_78 = 6'he == io_raddr ? regs_14 : _GEN_77; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_79 = 6'hf == io_raddr ? regs_15 : _GEN_78; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_80 = 6'h10 == io_raddr ? regs_16 : _GEN_79; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_81 = 6'h11 == io_raddr ? regs_17 : _GEN_80; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_82 = 6'h12 == io_raddr ? regs_18 : _GEN_81; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_83 = 6'h13 == io_raddr ? regs_19 : _GEN_82; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_84 = 6'h14 == io_raddr ? regs_20 : _GEN_83; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_85 = 6'h15 == io_raddr ? regs_21 : _GEN_84; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_86 = 6'h16 == io_raddr ? regs_22 : _GEN_85; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_87 = 6'h17 == io_raddr ? regs_23 : _GEN_86; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_88 = 6'h18 == io_raddr ? regs_24 : _GEN_87; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_89 = 6'h19 == io_raddr ? regs_25 : _GEN_88; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_90 = 6'h1a == io_raddr ? regs_26 : _GEN_89; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_91 = 6'h1b == io_raddr ? regs_27 : _GEN_90; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_92 = 6'h1c == io_raddr ? regs_28 : _GEN_91; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_93 = 6'h1d == io_raddr ? regs_29 : _GEN_92; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_94 = 6'h1e == io_raddr ? regs_30 : _GEN_93; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_95 = 6'h1f == io_raddr ? regs_31 : _GEN_94; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_96 = 6'h20 == io_raddr ? regs_32 : _GEN_95; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_97 = 6'h21 == io_raddr ? regs_33 : _GEN_96; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_98 = 6'h22 == io_raddr ? regs_34 : _GEN_97; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_99 = 6'h23 == io_raddr ? regs_35 : _GEN_98; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_100 = 6'h24 == io_raddr ? regs_36 : _GEN_99; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_101 = 6'h25 == io_raddr ? regs_37 : _GEN_100; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_102 = 6'h26 == io_raddr ? regs_38 : _GEN_101; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_103 = 6'h27 == io_raddr ? regs_39 : _GEN_102; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_104 = 6'h28 == io_raddr ? regs_40 : _GEN_103; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_105 = 6'h29 == io_raddr ? regs_41 : _GEN_104; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_106 = 6'h2a == io_raddr ? regs_42 : _GEN_105; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_107 = 6'h2b == io_raddr ? regs_43 : _GEN_106; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_108 = 6'h2c == io_raddr ? regs_44 : _GEN_107; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_109 = 6'h2d == io_raddr ? regs_45 : _GEN_108; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_110 = 6'h2e == io_raddr ? regs_46 : _GEN_109; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_111 = 6'h2f == io_raddr ? regs_47 : _GEN_110; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_112 = 6'h30 == io_raddr ? regs_48 : _GEN_111; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_113 = 6'h31 == io_raddr ? regs_49 : _GEN_112; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_114 = 6'h32 == io_raddr ? regs_50 : _GEN_113; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_115 = 6'h33 == io_raddr ? regs_51 : _GEN_114; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_116 = 6'h34 == io_raddr ? regs_52 : _GEN_115; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_117 = 6'h35 == io_raddr ? regs_53 : _GEN_116; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_118 = 6'h36 == io_raddr ? regs_54 : _GEN_117; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_119 = 6'h37 == io_raddr ? regs_55 : _GEN_118; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_120 = 6'h38 == io_raddr ? regs_56 : _GEN_119; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_121 = 6'h39 == io_raddr ? regs_57 : _GEN_120; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_122 = 6'h3a == io_raddr ? regs_58 : _GEN_121; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_123 = 6'h3b == io_raddr ? regs_59 : _GEN_122; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_124 = 6'h3c == io_raddr ? regs_60 : _GEN_123; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_125 = 6'h3d == io_raddr ? regs_61 : _GEN_124; // @[SRAM.scala 155:12:@50531.4]
  assign _GEN_126 = 6'h3e == io_raddr ? regs_62 : _GEN_125; // @[SRAM.scala 155:12:@50531.4]
  assign io_rdata = 6'h3f == io_raddr ? regs_63 : _GEN_126; // @[SRAM.scala 155:12:@50531.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_690) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_699) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_708) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_717) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_4 <= 1'h0;
    end else begin
      if (_T_726) begin
        if (io_banks_4_wdata_valid) begin
          regs_4 <= io_banks_4_wdata_bits;
        end else begin
          regs_4 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_5 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (io_banks_5_wdata_valid) begin
          regs_5 <= io_banks_5_wdata_bits;
        end else begin
          regs_5 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_6 <= 1'h0;
    end else begin
      if (_T_744) begin
        if (io_banks_6_wdata_valid) begin
          regs_6 <= io_banks_6_wdata_bits;
        end else begin
          regs_6 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_7 <= 1'h0;
    end else begin
      if (_T_753) begin
        if (io_banks_7_wdata_valid) begin
          regs_7 <= io_banks_7_wdata_bits;
        end else begin
          regs_7 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_8 <= 1'h0;
    end else begin
      if (_T_762) begin
        if (io_banks_8_wdata_valid) begin
          regs_8 <= io_banks_8_wdata_bits;
        end else begin
          regs_8 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_9 <= 1'h0;
    end else begin
      if (_T_771) begin
        if (io_banks_9_wdata_valid) begin
          regs_9 <= io_banks_9_wdata_bits;
        end else begin
          regs_9 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_10 <= 1'h0;
    end else begin
      if (_T_780) begin
        if (io_banks_10_wdata_valid) begin
          regs_10 <= io_banks_10_wdata_bits;
        end else begin
          regs_10 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_11 <= 1'h0;
    end else begin
      if (_T_789) begin
        if (io_banks_11_wdata_valid) begin
          regs_11 <= io_banks_11_wdata_bits;
        end else begin
          regs_11 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_12 <= 1'h0;
    end else begin
      if (_T_798) begin
        if (io_banks_12_wdata_valid) begin
          regs_12 <= io_banks_12_wdata_bits;
        end else begin
          regs_12 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_13 <= 1'h0;
    end else begin
      if (_T_807) begin
        if (io_banks_13_wdata_valid) begin
          regs_13 <= io_banks_13_wdata_bits;
        end else begin
          regs_13 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_14 <= 1'h0;
    end else begin
      if (_T_816) begin
        if (io_banks_14_wdata_valid) begin
          regs_14 <= io_banks_14_wdata_bits;
        end else begin
          regs_14 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_15 <= 1'h0;
    end else begin
      if (_T_825) begin
        if (io_banks_15_wdata_valid) begin
          regs_15 <= io_banks_15_wdata_bits;
        end else begin
          regs_15 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_16 <= 1'h0;
    end else begin
      if (_T_834) begin
        if (io_banks_16_wdata_valid) begin
          regs_16 <= io_banks_16_wdata_bits;
        end else begin
          regs_16 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_17 <= 1'h0;
    end else begin
      if (_T_843) begin
        if (io_banks_17_wdata_valid) begin
          regs_17 <= io_banks_17_wdata_bits;
        end else begin
          regs_17 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_18 <= 1'h0;
    end else begin
      if (_T_852) begin
        if (io_banks_18_wdata_valid) begin
          regs_18 <= io_banks_18_wdata_bits;
        end else begin
          regs_18 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_19 <= 1'h0;
    end else begin
      if (_T_861) begin
        if (io_banks_19_wdata_valid) begin
          regs_19 <= io_banks_19_wdata_bits;
        end else begin
          regs_19 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_20 <= 1'h0;
    end else begin
      if (_T_870) begin
        if (io_banks_20_wdata_valid) begin
          regs_20 <= io_banks_20_wdata_bits;
        end else begin
          regs_20 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_21 <= 1'h0;
    end else begin
      if (_T_879) begin
        if (io_banks_21_wdata_valid) begin
          regs_21 <= io_banks_21_wdata_bits;
        end else begin
          regs_21 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_22 <= 1'h0;
    end else begin
      if (_T_888) begin
        if (io_banks_22_wdata_valid) begin
          regs_22 <= io_banks_22_wdata_bits;
        end else begin
          regs_22 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_23 <= 1'h0;
    end else begin
      if (_T_897) begin
        if (io_banks_23_wdata_valid) begin
          regs_23 <= io_banks_23_wdata_bits;
        end else begin
          regs_23 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_24 <= 1'h0;
    end else begin
      if (_T_906) begin
        if (io_banks_24_wdata_valid) begin
          regs_24 <= io_banks_24_wdata_bits;
        end else begin
          regs_24 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_25 <= 1'h0;
    end else begin
      if (_T_915) begin
        if (io_banks_25_wdata_valid) begin
          regs_25 <= io_banks_25_wdata_bits;
        end else begin
          regs_25 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_26 <= 1'h0;
    end else begin
      if (_T_924) begin
        if (io_banks_26_wdata_valid) begin
          regs_26 <= io_banks_26_wdata_bits;
        end else begin
          regs_26 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_27 <= 1'h0;
    end else begin
      if (_T_933) begin
        if (io_banks_27_wdata_valid) begin
          regs_27 <= io_banks_27_wdata_bits;
        end else begin
          regs_27 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_28 <= 1'h0;
    end else begin
      if (_T_942) begin
        if (io_banks_28_wdata_valid) begin
          regs_28 <= io_banks_28_wdata_bits;
        end else begin
          regs_28 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_29 <= 1'h0;
    end else begin
      if (_T_951) begin
        if (io_banks_29_wdata_valid) begin
          regs_29 <= io_banks_29_wdata_bits;
        end else begin
          regs_29 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_30 <= 1'h0;
    end else begin
      if (_T_960) begin
        if (io_banks_30_wdata_valid) begin
          regs_30 <= io_banks_30_wdata_bits;
        end else begin
          regs_30 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_31 <= 1'h0;
    end else begin
      if (_T_969) begin
        if (io_banks_31_wdata_valid) begin
          regs_31 <= io_banks_31_wdata_bits;
        end else begin
          regs_31 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_32 <= 1'h0;
    end else begin
      if (_T_978) begin
        if (io_banks_32_wdata_valid) begin
          regs_32 <= io_banks_32_wdata_bits;
        end else begin
          regs_32 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_33 <= 1'h0;
    end else begin
      if (_T_987) begin
        if (io_banks_33_wdata_valid) begin
          regs_33 <= io_banks_33_wdata_bits;
        end else begin
          regs_33 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_34 <= 1'h0;
    end else begin
      if (_T_996) begin
        if (io_banks_34_wdata_valid) begin
          regs_34 <= io_banks_34_wdata_bits;
        end else begin
          regs_34 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_35 <= 1'h0;
    end else begin
      if (_T_1005) begin
        if (io_banks_35_wdata_valid) begin
          regs_35 <= io_banks_35_wdata_bits;
        end else begin
          regs_35 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_36 <= 1'h0;
    end else begin
      if (_T_1014) begin
        if (io_banks_36_wdata_valid) begin
          regs_36 <= io_banks_36_wdata_bits;
        end else begin
          regs_36 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_37 <= 1'h0;
    end else begin
      if (_T_1023) begin
        if (io_banks_37_wdata_valid) begin
          regs_37 <= io_banks_37_wdata_bits;
        end else begin
          regs_37 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_38 <= 1'h0;
    end else begin
      if (_T_1032) begin
        if (io_banks_38_wdata_valid) begin
          regs_38 <= io_banks_38_wdata_bits;
        end else begin
          regs_38 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_39 <= 1'h0;
    end else begin
      if (_T_1041) begin
        if (io_banks_39_wdata_valid) begin
          regs_39 <= io_banks_39_wdata_bits;
        end else begin
          regs_39 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_40 <= 1'h0;
    end else begin
      if (_T_1050) begin
        if (io_banks_40_wdata_valid) begin
          regs_40 <= io_banks_40_wdata_bits;
        end else begin
          regs_40 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_41 <= 1'h0;
    end else begin
      if (_T_1059) begin
        if (io_banks_41_wdata_valid) begin
          regs_41 <= io_banks_41_wdata_bits;
        end else begin
          regs_41 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_42 <= 1'h0;
    end else begin
      if (_T_1068) begin
        if (io_banks_42_wdata_valid) begin
          regs_42 <= io_banks_42_wdata_bits;
        end else begin
          regs_42 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_43 <= 1'h0;
    end else begin
      if (_T_1077) begin
        if (io_banks_43_wdata_valid) begin
          regs_43 <= io_banks_43_wdata_bits;
        end else begin
          regs_43 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_44 <= 1'h0;
    end else begin
      if (_T_1086) begin
        if (io_banks_44_wdata_valid) begin
          regs_44 <= io_banks_44_wdata_bits;
        end else begin
          regs_44 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_45 <= 1'h0;
    end else begin
      if (_T_1095) begin
        if (io_banks_45_wdata_valid) begin
          regs_45 <= io_banks_45_wdata_bits;
        end else begin
          regs_45 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_46 <= 1'h0;
    end else begin
      if (_T_1104) begin
        if (io_banks_46_wdata_valid) begin
          regs_46 <= io_banks_46_wdata_bits;
        end else begin
          regs_46 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_47 <= 1'h0;
    end else begin
      if (_T_1113) begin
        if (io_banks_47_wdata_valid) begin
          regs_47 <= io_banks_47_wdata_bits;
        end else begin
          regs_47 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_48 <= 1'h0;
    end else begin
      if (_T_1122) begin
        if (io_banks_48_wdata_valid) begin
          regs_48 <= io_banks_48_wdata_bits;
        end else begin
          regs_48 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_49 <= 1'h0;
    end else begin
      if (_T_1131) begin
        if (io_banks_49_wdata_valid) begin
          regs_49 <= io_banks_49_wdata_bits;
        end else begin
          regs_49 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_50 <= 1'h0;
    end else begin
      if (_T_1140) begin
        if (io_banks_50_wdata_valid) begin
          regs_50 <= io_banks_50_wdata_bits;
        end else begin
          regs_50 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_51 <= 1'h0;
    end else begin
      if (_T_1149) begin
        if (io_banks_51_wdata_valid) begin
          regs_51 <= io_banks_51_wdata_bits;
        end else begin
          regs_51 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_52 <= 1'h0;
    end else begin
      if (_T_1158) begin
        if (io_banks_52_wdata_valid) begin
          regs_52 <= io_banks_52_wdata_bits;
        end else begin
          regs_52 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_53 <= 1'h0;
    end else begin
      if (_T_1167) begin
        if (io_banks_53_wdata_valid) begin
          regs_53 <= io_banks_53_wdata_bits;
        end else begin
          regs_53 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_54 <= 1'h0;
    end else begin
      if (_T_1176) begin
        if (io_banks_54_wdata_valid) begin
          regs_54 <= io_banks_54_wdata_bits;
        end else begin
          regs_54 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_55 <= 1'h0;
    end else begin
      if (_T_1185) begin
        if (io_banks_55_wdata_valid) begin
          regs_55 <= io_banks_55_wdata_bits;
        end else begin
          regs_55 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_56 <= 1'h0;
    end else begin
      if (_T_1194) begin
        if (io_banks_56_wdata_valid) begin
          regs_56 <= io_banks_56_wdata_bits;
        end else begin
          regs_56 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_57 <= 1'h0;
    end else begin
      if (_T_1203) begin
        if (io_banks_57_wdata_valid) begin
          regs_57 <= io_banks_57_wdata_bits;
        end else begin
          regs_57 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_58 <= 1'h0;
    end else begin
      if (_T_1212) begin
        if (io_banks_58_wdata_valid) begin
          regs_58 <= io_banks_58_wdata_bits;
        end else begin
          regs_58 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_59 <= 1'h0;
    end else begin
      if (_T_1221) begin
        if (io_banks_59_wdata_valid) begin
          regs_59 <= io_banks_59_wdata_bits;
        end else begin
          regs_59 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_60 <= 1'h0;
    end else begin
      if (_T_1230) begin
        if (io_banks_60_wdata_valid) begin
          regs_60 <= io_banks_60_wdata_bits;
        end else begin
          regs_60 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_61 <= 1'h0;
    end else begin
      if (_T_1239) begin
        if (io_banks_61_wdata_valid) begin
          regs_61 <= io_banks_61_wdata_bits;
        end else begin
          regs_61 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_62 <= 1'h0;
    end else begin
      if (_T_1248) begin
        if (io_banks_62_wdata_valid) begin
          regs_62 <= io_banks_62_wdata_bits;
        end else begin
          regs_62 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_63 <= 1'h0;
    end else begin
      if (_T_1257) begin
        if (io_banks_63_wdata_valid) begin
          regs_63 <= io_banks_63_wdata_bits;
        end else begin
          regs_63 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_33( // @[:@50533.2]
  input   clock, // @[:@50534.4]
  input   reset, // @[:@50535.4]
  output  io_in_ready, // @[:@50536.4]
  input   io_in_valid, // @[:@50536.4]
  input   io_in_bits, // @[:@50536.4]
  input   io_out_ready, // @[:@50536.4]
  output  io_out_valid, // @[:@50536.4]
  output  io_out_bits, // @[:@50536.4]
  input   io_banks_0_wdata_valid, // @[:@50536.4]
  input   io_banks_0_wdata_bits, // @[:@50536.4]
  input   io_banks_1_wdata_valid, // @[:@50536.4]
  input   io_banks_1_wdata_bits, // @[:@50536.4]
  input   io_banks_2_wdata_valid, // @[:@50536.4]
  input   io_banks_2_wdata_bits, // @[:@50536.4]
  input   io_banks_3_wdata_valid, // @[:@50536.4]
  input   io_banks_3_wdata_bits, // @[:@50536.4]
  input   io_banks_4_wdata_valid, // @[:@50536.4]
  input   io_banks_4_wdata_bits, // @[:@50536.4]
  input   io_banks_5_wdata_valid, // @[:@50536.4]
  input   io_banks_5_wdata_bits, // @[:@50536.4]
  input   io_banks_6_wdata_valid, // @[:@50536.4]
  input   io_banks_6_wdata_bits, // @[:@50536.4]
  input   io_banks_7_wdata_valid, // @[:@50536.4]
  input   io_banks_7_wdata_bits, // @[:@50536.4]
  input   io_banks_8_wdata_valid, // @[:@50536.4]
  input   io_banks_8_wdata_bits, // @[:@50536.4]
  input   io_banks_9_wdata_valid, // @[:@50536.4]
  input   io_banks_9_wdata_bits, // @[:@50536.4]
  input   io_banks_10_wdata_valid, // @[:@50536.4]
  input   io_banks_10_wdata_bits, // @[:@50536.4]
  input   io_banks_11_wdata_valid, // @[:@50536.4]
  input   io_banks_11_wdata_bits, // @[:@50536.4]
  input   io_banks_12_wdata_valid, // @[:@50536.4]
  input   io_banks_12_wdata_bits, // @[:@50536.4]
  input   io_banks_13_wdata_valid, // @[:@50536.4]
  input   io_banks_13_wdata_bits, // @[:@50536.4]
  input   io_banks_14_wdata_valid, // @[:@50536.4]
  input   io_banks_14_wdata_bits, // @[:@50536.4]
  input   io_banks_15_wdata_valid, // @[:@50536.4]
  input   io_banks_15_wdata_bits, // @[:@50536.4]
  input   io_banks_16_wdata_valid, // @[:@50536.4]
  input   io_banks_16_wdata_bits, // @[:@50536.4]
  input   io_banks_17_wdata_valid, // @[:@50536.4]
  input   io_banks_17_wdata_bits, // @[:@50536.4]
  input   io_banks_18_wdata_valid, // @[:@50536.4]
  input   io_banks_18_wdata_bits, // @[:@50536.4]
  input   io_banks_19_wdata_valid, // @[:@50536.4]
  input   io_banks_19_wdata_bits, // @[:@50536.4]
  input   io_banks_20_wdata_valid, // @[:@50536.4]
  input   io_banks_20_wdata_bits, // @[:@50536.4]
  input   io_banks_21_wdata_valid, // @[:@50536.4]
  input   io_banks_21_wdata_bits, // @[:@50536.4]
  input   io_banks_22_wdata_valid, // @[:@50536.4]
  input   io_banks_22_wdata_bits, // @[:@50536.4]
  input   io_banks_23_wdata_valid, // @[:@50536.4]
  input   io_banks_23_wdata_bits, // @[:@50536.4]
  input   io_banks_24_wdata_valid, // @[:@50536.4]
  input   io_banks_24_wdata_bits, // @[:@50536.4]
  input   io_banks_25_wdata_valid, // @[:@50536.4]
  input   io_banks_25_wdata_bits, // @[:@50536.4]
  input   io_banks_26_wdata_valid, // @[:@50536.4]
  input   io_banks_26_wdata_bits, // @[:@50536.4]
  input   io_banks_27_wdata_valid, // @[:@50536.4]
  input   io_banks_27_wdata_bits, // @[:@50536.4]
  input   io_banks_28_wdata_valid, // @[:@50536.4]
  input   io_banks_28_wdata_bits, // @[:@50536.4]
  input   io_banks_29_wdata_valid, // @[:@50536.4]
  input   io_banks_29_wdata_bits, // @[:@50536.4]
  input   io_banks_30_wdata_valid, // @[:@50536.4]
  input   io_banks_30_wdata_bits, // @[:@50536.4]
  input   io_banks_31_wdata_valid, // @[:@50536.4]
  input   io_banks_31_wdata_bits, // @[:@50536.4]
  input   io_banks_32_wdata_valid, // @[:@50536.4]
  input   io_banks_32_wdata_bits, // @[:@50536.4]
  input   io_banks_33_wdata_valid, // @[:@50536.4]
  input   io_banks_33_wdata_bits, // @[:@50536.4]
  input   io_banks_34_wdata_valid, // @[:@50536.4]
  input   io_banks_34_wdata_bits, // @[:@50536.4]
  input   io_banks_35_wdata_valid, // @[:@50536.4]
  input   io_banks_35_wdata_bits, // @[:@50536.4]
  input   io_banks_36_wdata_valid, // @[:@50536.4]
  input   io_banks_36_wdata_bits, // @[:@50536.4]
  input   io_banks_37_wdata_valid, // @[:@50536.4]
  input   io_banks_37_wdata_bits, // @[:@50536.4]
  input   io_banks_38_wdata_valid, // @[:@50536.4]
  input   io_banks_38_wdata_bits, // @[:@50536.4]
  input   io_banks_39_wdata_valid, // @[:@50536.4]
  input   io_banks_39_wdata_bits, // @[:@50536.4]
  input   io_banks_40_wdata_valid, // @[:@50536.4]
  input   io_banks_40_wdata_bits, // @[:@50536.4]
  input   io_banks_41_wdata_valid, // @[:@50536.4]
  input   io_banks_41_wdata_bits, // @[:@50536.4]
  input   io_banks_42_wdata_valid, // @[:@50536.4]
  input   io_banks_42_wdata_bits, // @[:@50536.4]
  input   io_banks_43_wdata_valid, // @[:@50536.4]
  input   io_banks_43_wdata_bits, // @[:@50536.4]
  input   io_banks_44_wdata_valid, // @[:@50536.4]
  input   io_banks_44_wdata_bits, // @[:@50536.4]
  input   io_banks_45_wdata_valid, // @[:@50536.4]
  input   io_banks_45_wdata_bits, // @[:@50536.4]
  input   io_banks_46_wdata_valid, // @[:@50536.4]
  input   io_banks_46_wdata_bits, // @[:@50536.4]
  input   io_banks_47_wdata_valid, // @[:@50536.4]
  input   io_banks_47_wdata_bits, // @[:@50536.4]
  input   io_banks_48_wdata_valid, // @[:@50536.4]
  input   io_banks_48_wdata_bits, // @[:@50536.4]
  input   io_banks_49_wdata_valid, // @[:@50536.4]
  input   io_banks_49_wdata_bits, // @[:@50536.4]
  input   io_banks_50_wdata_valid, // @[:@50536.4]
  input   io_banks_50_wdata_bits, // @[:@50536.4]
  input   io_banks_51_wdata_valid, // @[:@50536.4]
  input   io_banks_51_wdata_bits, // @[:@50536.4]
  input   io_banks_52_wdata_valid, // @[:@50536.4]
  input   io_banks_52_wdata_bits, // @[:@50536.4]
  input   io_banks_53_wdata_valid, // @[:@50536.4]
  input   io_banks_53_wdata_bits, // @[:@50536.4]
  input   io_banks_54_wdata_valid, // @[:@50536.4]
  input   io_banks_54_wdata_bits, // @[:@50536.4]
  input   io_banks_55_wdata_valid, // @[:@50536.4]
  input   io_banks_55_wdata_bits, // @[:@50536.4]
  input   io_banks_56_wdata_valid, // @[:@50536.4]
  input   io_banks_56_wdata_bits, // @[:@50536.4]
  input   io_banks_57_wdata_valid, // @[:@50536.4]
  input   io_banks_57_wdata_bits, // @[:@50536.4]
  input   io_banks_58_wdata_valid, // @[:@50536.4]
  input   io_banks_58_wdata_bits, // @[:@50536.4]
  input   io_banks_59_wdata_valid, // @[:@50536.4]
  input   io_banks_59_wdata_bits, // @[:@50536.4]
  input   io_banks_60_wdata_valid, // @[:@50536.4]
  input   io_banks_60_wdata_bits, // @[:@50536.4]
  input   io_banks_61_wdata_valid, // @[:@50536.4]
  input   io_banks_61_wdata_bits, // @[:@50536.4]
  input   io_banks_62_wdata_valid, // @[:@50536.4]
  input   io_banks_62_wdata_bits, // @[:@50536.4]
  input   io_banks_63_wdata_valid, // @[:@50536.4]
  input   io_banks_63_wdata_bits // @[:@50536.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@50802.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@50802.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@50802.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@50802.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@50802.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@50812.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@50812.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@50812.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@50812.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@50812.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@50827.4]
  wire [5:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@50827.4]
  wire [5:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_4_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_4_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_5_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_5_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_6_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_6_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_7_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_7_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_8_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_8_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_9_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_9_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_10_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_10_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_11_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_11_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_12_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_12_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_13_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_13_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_14_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_14_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_15_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_15_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_16_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_16_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_17_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_17_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_18_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_18_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_19_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_19_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_20_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_20_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_21_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_21_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_22_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_22_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_23_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_23_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_24_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_24_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_25_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_25_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_26_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_26_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_27_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_27_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_28_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_28_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_29_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_29_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_30_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_30_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_31_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_31_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_32_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_32_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_33_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_33_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_34_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_34_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_35_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_35_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_36_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_36_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_37_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_37_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_38_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_38_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_39_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_39_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_40_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_40_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_41_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_41_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_42_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_42_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_43_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_43_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_44_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_44_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_45_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_45_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_46_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_46_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_47_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_47_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_48_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_48_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_49_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_49_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_50_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_50_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_51_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_51_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_52_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_52_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_53_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_53_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_54_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_54_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_55_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_55_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_56_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_56_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_57_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_57_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_58_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_58_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_59_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_59_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_60_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_60_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_61_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_61_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_62_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_62_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_63_wdata_valid; // @[FIFO.scala 49:19:@50827.4]
  wire  FFRAM_io_banks_63_wdata_bits; // @[FIFO.scala 49:19:@50827.4]
  wire  writeEn; // @[FIFO.scala 30:29:@50800.4]
  wire  readEn; // @[FIFO.scala 31:29:@50801.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@50822.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@50823.4]
  wire  _T_824; // @[FIFO.scala 45:27:@50824.4]
  wire  empty; // @[FIFO.scala 45:24:@50825.4]
  wire  full; // @[FIFO.scala 46:23:@50826.4]
  wire  _T_1657; // @[FIFO.scala 83:17:@51993.4]
  wire  _GEN_64; // @[FIFO.scala 83:29:@51994.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@50802.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@50812.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM_16 FFRAM ( // @[FIFO.scala 49:19:@50827.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(FFRAM_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(FFRAM_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(FFRAM_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(FFRAM_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(FFRAM_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(FFRAM_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(FFRAM_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(FFRAM_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(FFRAM_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(FFRAM_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(FFRAM_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(FFRAM_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(FFRAM_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(FFRAM_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(FFRAM_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(FFRAM_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(FFRAM_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(FFRAM_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(FFRAM_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(FFRAM_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(FFRAM_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(FFRAM_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(FFRAM_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(FFRAM_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(FFRAM_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(FFRAM_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(FFRAM_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(FFRAM_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(FFRAM_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(FFRAM_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(FFRAM_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(FFRAM_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(FFRAM_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(FFRAM_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(FFRAM_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(FFRAM_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(FFRAM_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(FFRAM_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(FFRAM_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(FFRAM_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(FFRAM_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(FFRAM_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(FFRAM_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(FFRAM_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(FFRAM_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(FFRAM_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(FFRAM_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(FFRAM_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(FFRAM_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(FFRAM_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(FFRAM_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(FFRAM_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(FFRAM_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(FFRAM_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(FFRAM_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(FFRAM_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(FFRAM_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(FFRAM_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(FFRAM_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(FFRAM_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(FFRAM_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(FFRAM_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(FFRAM_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(FFRAM_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(FFRAM_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(FFRAM_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(FFRAM_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(FFRAM_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(FFRAM_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(FFRAM_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(FFRAM_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(FFRAM_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(FFRAM_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(FFRAM_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(FFRAM_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(FFRAM_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(FFRAM_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(FFRAM_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(FFRAM_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(FFRAM_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(FFRAM_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(FFRAM_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(FFRAM_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(FFRAM_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(FFRAM_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(FFRAM_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(FFRAM_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(FFRAM_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(FFRAM_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(FFRAM_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(FFRAM_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(FFRAM_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(FFRAM_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(FFRAM_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(FFRAM_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(FFRAM_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(FFRAM_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(FFRAM_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(FFRAM_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(FFRAM_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(FFRAM_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(FFRAM_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(FFRAM_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(FFRAM_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(FFRAM_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(FFRAM_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(FFRAM_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(FFRAM_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(FFRAM_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(FFRAM_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(FFRAM_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(FFRAM_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(FFRAM_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(FFRAM_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(FFRAM_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(FFRAM_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(FFRAM_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(FFRAM_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(FFRAM_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(FFRAM_io_banks_63_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@50800.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@50801.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@50823.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@50824.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@50825.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@50826.4]
  assign _T_1657 = writeEn != readEn; // @[FIFO.scala 83:17:@51993.4]
  assign _GEN_64 = _T_1657 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@51994.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@52000.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@51998.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@51032.4]
  assign enqCounter_clock = clock; // @[:@50803.4]
  assign enqCounter_reset = reset; // @[:@50804.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@50810.4]
  assign deqCounter_clock = clock; // @[:@50813.4]
  assign deqCounter_reset = reset; // @[:@50814.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@50820.4]
  assign FFRAM_clock = clock; // @[:@50828.4]
  assign FFRAM_reset = reset; // @[:@50829.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@51028.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@51029.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@51030.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@51031.4]
  assign FFRAM_io_banks_0_wdata_valid = io_banks_0_wdata_valid; // @[FIFO.scala 59:15:@51034.4]
  assign FFRAM_io_banks_0_wdata_bits = io_banks_0_wdata_bits; // @[FIFO.scala 59:15:@51033.4]
  assign FFRAM_io_banks_1_wdata_valid = io_banks_1_wdata_valid; // @[FIFO.scala 59:15:@51037.4]
  assign FFRAM_io_banks_1_wdata_bits = io_banks_1_wdata_bits; // @[FIFO.scala 59:15:@51036.4]
  assign FFRAM_io_banks_2_wdata_valid = io_banks_2_wdata_valid; // @[FIFO.scala 59:15:@51040.4]
  assign FFRAM_io_banks_2_wdata_bits = io_banks_2_wdata_bits; // @[FIFO.scala 59:15:@51039.4]
  assign FFRAM_io_banks_3_wdata_valid = io_banks_3_wdata_valid; // @[FIFO.scala 59:15:@51043.4]
  assign FFRAM_io_banks_3_wdata_bits = io_banks_3_wdata_bits; // @[FIFO.scala 59:15:@51042.4]
  assign FFRAM_io_banks_4_wdata_valid = io_banks_4_wdata_valid; // @[FIFO.scala 59:15:@51046.4]
  assign FFRAM_io_banks_4_wdata_bits = io_banks_4_wdata_bits; // @[FIFO.scala 59:15:@51045.4]
  assign FFRAM_io_banks_5_wdata_valid = io_banks_5_wdata_valid; // @[FIFO.scala 59:15:@51049.4]
  assign FFRAM_io_banks_5_wdata_bits = io_banks_5_wdata_bits; // @[FIFO.scala 59:15:@51048.4]
  assign FFRAM_io_banks_6_wdata_valid = io_banks_6_wdata_valid; // @[FIFO.scala 59:15:@51052.4]
  assign FFRAM_io_banks_6_wdata_bits = io_banks_6_wdata_bits; // @[FIFO.scala 59:15:@51051.4]
  assign FFRAM_io_banks_7_wdata_valid = io_banks_7_wdata_valid; // @[FIFO.scala 59:15:@51055.4]
  assign FFRAM_io_banks_7_wdata_bits = io_banks_7_wdata_bits; // @[FIFO.scala 59:15:@51054.4]
  assign FFRAM_io_banks_8_wdata_valid = io_banks_8_wdata_valid; // @[FIFO.scala 59:15:@51058.4]
  assign FFRAM_io_banks_8_wdata_bits = io_banks_8_wdata_bits; // @[FIFO.scala 59:15:@51057.4]
  assign FFRAM_io_banks_9_wdata_valid = io_banks_9_wdata_valid; // @[FIFO.scala 59:15:@51061.4]
  assign FFRAM_io_banks_9_wdata_bits = io_banks_9_wdata_bits; // @[FIFO.scala 59:15:@51060.4]
  assign FFRAM_io_banks_10_wdata_valid = io_banks_10_wdata_valid; // @[FIFO.scala 59:15:@51064.4]
  assign FFRAM_io_banks_10_wdata_bits = io_banks_10_wdata_bits; // @[FIFO.scala 59:15:@51063.4]
  assign FFRAM_io_banks_11_wdata_valid = io_banks_11_wdata_valid; // @[FIFO.scala 59:15:@51067.4]
  assign FFRAM_io_banks_11_wdata_bits = io_banks_11_wdata_bits; // @[FIFO.scala 59:15:@51066.4]
  assign FFRAM_io_banks_12_wdata_valid = io_banks_12_wdata_valid; // @[FIFO.scala 59:15:@51070.4]
  assign FFRAM_io_banks_12_wdata_bits = io_banks_12_wdata_bits; // @[FIFO.scala 59:15:@51069.4]
  assign FFRAM_io_banks_13_wdata_valid = io_banks_13_wdata_valid; // @[FIFO.scala 59:15:@51073.4]
  assign FFRAM_io_banks_13_wdata_bits = io_banks_13_wdata_bits; // @[FIFO.scala 59:15:@51072.4]
  assign FFRAM_io_banks_14_wdata_valid = io_banks_14_wdata_valid; // @[FIFO.scala 59:15:@51076.4]
  assign FFRAM_io_banks_14_wdata_bits = io_banks_14_wdata_bits; // @[FIFO.scala 59:15:@51075.4]
  assign FFRAM_io_banks_15_wdata_valid = io_banks_15_wdata_valid; // @[FIFO.scala 59:15:@51079.4]
  assign FFRAM_io_banks_15_wdata_bits = io_banks_15_wdata_bits; // @[FIFO.scala 59:15:@51078.4]
  assign FFRAM_io_banks_16_wdata_valid = io_banks_16_wdata_valid; // @[FIFO.scala 59:15:@51082.4]
  assign FFRAM_io_banks_16_wdata_bits = io_banks_16_wdata_bits; // @[FIFO.scala 59:15:@51081.4]
  assign FFRAM_io_banks_17_wdata_valid = io_banks_17_wdata_valid; // @[FIFO.scala 59:15:@51085.4]
  assign FFRAM_io_banks_17_wdata_bits = io_banks_17_wdata_bits; // @[FIFO.scala 59:15:@51084.4]
  assign FFRAM_io_banks_18_wdata_valid = io_banks_18_wdata_valid; // @[FIFO.scala 59:15:@51088.4]
  assign FFRAM_io_banks_18_wdata_bits = io_banks_18_wdata_bits; // @[FIFO.scala 59:15:@51087.4]
  assign FFRAM_io_banks_19_wdata_valid = io_banks_19_wdata_valid; // @[FIFO.scala 59:15:@51091.4]
  assign FFRAM_io_banks_19_wdata_bits = io_banks_19_wdata_bits; // @[FIFO.scala 59:15:@51090.4]
  assign FFRAM_io_banks_20_wdata_valid = io_banks_20_wdata_valid; // @[FIFO.scala 59:15:@51094.4]
  assign FFRAM_io_banks_20_wdata_bits = io_banks_20_wdata_bits; // @[FIFO.scala 59:15:@51093.4]
  assign FFRAM_io_banks_21_wdata_valid = io_banks_21_wdata_valid; // @[FIFO.scala 59:15:@51097.4]
  assign FFRAM_io_banks_21_wdata_bits = io_banks_21_wdata_bits; // @[FIFO.scala 59:15:@51096.4]
  assign FFRAM_io_banks_22_wdata_valid = io_banks_22_wdata_valid; // @[FIFO.scala 59:15:@51100.4]
  assign FFRAM_io_banks_22_wdata_bits = io_banks_22_wdata_bits; // @[FIFO.scala 59:15:@51099.4]
  assign FFRAM_io_banks_23_wdata_valid = io_banks_23_wdata_valid; // @[FIFO.scala 59:15:@51103.4]
  assign FFRAM_io_banks_23_wdata_bits = io_banks_23_wdata_bits; // @[FIFO.scala 59:15:@51102.4]
  assign FFRAM_io_banks_24_wdata_valid = io_banks_24_wdata_valid; // @[FIFO.scala 59:15:@51106.4]
  assign FFRAM_io_banks_24_wdata_bits = io_banks_24_wdata_bits; // @[FIFO.scala 59:15:@51105.4]
  assign FFRAM_io_banks_25_wdata_valid = io_banks_25_wdata_valid; // @[FIFO.scala 59:15:@51109.4]
  assign FFRAM_io_banks_25_wdata_bits = io_banks_25_wdata_bits; // @[FIFO.scala 59:15:@51108.4]
  assign FFRAM_io_banks_26_wdata_valid = io_banks_26_wdata_valid; // @[FIFO.scala 59:15:@51112.4]
  assign FFRAM_io_banks_26_wdata_bits = io_banks_26_wdata_bits; // @[FIFO.scala 59:15:@51111.4]
  assign FFRAM_io_banks_27_wdata_valid = io_banks_27_wdata_valid; // @[FIFO.scala 59:15:@51115.4]
  assign FFRAM_io_banks_27_wdata_bits = io_banks_27_wdata_bits; // @[FIFO.scala 59:15:@51114.4]
  assign FFRAM_io_banks_28_wdata_valid = io_banks_28_wdata_valid; // @[FIFO.scala 59:15:@51118.4]
  assign FFRAM_io_banks_28_wdata_bits = io_banks_28_wdata_bits; // @[FIFO.scala 59:15:@51117.4]
  assign FFRAM_io_banks_29_wdata_valid = io_banks_29_wdata_valid; // @[FIFO.scala 59:15:@51121.4]
  assign FFRAM_io_banks_29_wdata_bits = io_banks_29_wdata_bits; // @[FIFO.scala 59:15:@51120.4]
  assign FFRAM_io_banks_30_wdata_valid = io_banks_30_wdata_valid; // @[FIFO.scala 59:15:@51124.4]
  assign FFRAM_io_banks_30_wdata_bits = io_banks_30_wdata_bits; // @[FIFO.scala 59:15:@51123.4]
  assign FFRAM_io_banks_31_wdata_valid = io_banks_31_wdata_valid; // @[FIFO.scala 59:15:@51127.4]
  assign FFRAM_io_banks_31_wdata_bits = io_banks_31_wdata_bits; // @[FIFO.scala 59:15:@51126.4]
  assign FFRAM_io_banks_32_wdata_valid = io_banks_32_wdata_valid; // @[FIFO.scala 59:15:@51130.4]
  assign FFRAM_io_banks_32_wdata_bits = io_banks_32_wdata_bits; // @[FIFO.scala 59:15:@51129.4]
  assign FFRAM_io_banks_33_wdata_valid = io_banks_33_wdata_valid; // @[FIFO.scala 59:15:@51133.4]
  assign FFRAM_io_banks_33_wdata_bits = io_banks_33_wdata_bits; // @[FIFO.scala 59:15:@51132.4]
  assign FFRAM_io_banks_34_wdata_valid = io_banks_34_wdata_valid; // @[FIFO.scala 59:15:@51136.4]
  assign FFRAM_io_banks_34_wdata_bits = io_banks_34_wdata_bits; // @[FIFO.scala 59:15:@51135.4]
  assign FFRAM_io_banks_35_wdata_valid = io_banks_35_wdata_valid; // @[FIFO.scala 59:15:@51139.4]
  assign FFRAM_io_banks_35_wdata_bits = io_banks_35_wdata_bits; // @[FIFO.scala 59:15:@51138.4]
  assign FFRAM_io_banks_36_wdata_valid = io_banks_36_wdata_valid; // @[FIFO.scala 59:15:@51142.4]
  assign FFRAM_io_banks_36_wdata_bits = io_banks_36_wdata_bits; // @[FIFO.scala 59:15:@51141.4]
  assign FFRAM_io_banks_37_wdata_valid = io_banks_37_wdata_valid; // @[FIFO.scala 59:15:@51145.4]
  assign FFRAM_io_banks_37_wdata_bits = io_banks_37_wdata_bits; // @[FIFO.scala 59:15:@51144.4]
  assign FFRAM_io_banks_38_wdata_valid = io_banks_38_wdata_valid; // @[FIFO.scala 59:15:@51148.4]
  assign FFRAM_io_banks_38_wdata_bits = io_banks_38_wdata_bits; // @[FIFO.scala 59:15:@51147.4]
  assign FFRAM_io_banks_39_wdata_valid = io_banks_39_wdata_valid; // @[FIFO.scala 59:15:@51151.4]
  assign FFRAM_io_banks_39_wdata_bits = io_banks_39_wdata_bits; // @[FIFO.scala 59:15:@51150.4]
  assign FFRAM_io_banks_40_wdata_valid = io_banks_40_wdata_valid; // @[FIFO.scala 59:15:@51154.4]
  assign FFRAM_io_banks_40_wdata_bits = io_banks_40_wdata_bits; // @[FIFO.scala 59:15:@51153.4]
  assign FFRAM_io_banks_41_wdata_valid = io_banks_41_wdata_valid; // @[FIFO.scala 59:15:@51157.4]
  assign FFRAM_io_banks_41_wdata_bits = io_banks_41_wdata_bits; // @[FIFO.scala 59:15:@51156.4]
  assign FFRAM_io_banks_42_wdata_valid = io_banks_42_wdata_valid; // @[FIFO.scala 59:15:@51160.4]
  assign FFRAM_io_banks_42_wdata_bits = io_banks_42_wdata_bits; // @[FIFO.scala 59:15:@51159.4]
  assign FFRAM_io_banks_43_wdata_valid = io_banks_43_wdata_valid; // @[FIFO.scala 59:15:@51163.4]
  assign FFRAM_io_banks_43_wdata_bits = io_banks_43_wdata_bits; // @[FIFO.scala 59:15:@51162.4]
  assign FFRAM_io_banks_44_wdata_valid = io_banks_44_wdata_valid; // @[FIFO.scala 59:15:@51166.4]
  assign FFRAM_io_banks_44_wdata_bits = io_banks_44_wdata_bits; // @[FIFO.scala 59:15:@51165.4]
  assign FFRAM_io_banks_45_wdata_valid = io_banks_45_wdata_valid; // @[FIFO.scala 59:15:@51169.4]
  assign FFRAM_io_banks_45_wdata_bits = io_banks_45_wdata_bits; // @[FIFO.scala 59:15:@51168.4]
  assign FFRAM_io_banks_46_wdata_valid = io_banks_46_wdata_valid; // @[FIFO.scala 59:15:@51172.4]
  assign FFRAM_io_banks_46_wdata_bits = io_banks_46_wdata_bits; // @[FIFO.scala 59:15:@51171.4]
  assign FFRAM_io_banks_47_wdata_valid = io_banks_47_wdata_valid; // @[FIFO.scala 59:15:@51175.4]
  assign FFRAM_io_banks_47_wdata_bits = io_banks_47_wdata_bits; // @[FIFO.scala 59:15:@51174.4]
  assign FFRAM_io_banks_48_wdata_valid = io_banks_48_wdata_valid; // @[FIFO.scala 59:15:@51178.4]
  assign FFRAM_io_banks_48_wdata_bits = io_banks_48_wdata_bits; // @[FIFO.scala 59:15:@51177.4]
  assign FFRAM_io_banks_49_wdata_valid = io_banks_49_wdata_valid; // @[FIFO.scala 59:15:@51181.4]
  assign FFRAM_io_banks_49_wdata_bits = io_banks_49_wdata_bits; // @[FIFO.scala 59:15:@51180.4]
  assign FFRAM_io_banks_50_wdata_valid = io_banks_50_wdata_valid; // @[FIFO.scala 59:15:@51184.4]
  assign FFRAM_io_banks_50_wdata_bits = io_banks_50_wdata_bits; // @[FIFO.scala 59:15:@51183.4]
  assign FFRAM_io_banks_51_wdata_valid = io_banks_51_wdata_valid; // @[FIFO.scala 59:15:@51187.4]
  assign FFRAM_io_banks_51_wdata_bits = io_banks_51_wdata_bits; // @[FIFO.scala 59:15:@51186.4]
  assign FFRAM_io_banks_52_wdata_valid = io_banks_52_wdata_valid; // @[FIFO.scala 59:15:@51190.4]
  assign FFRAM_io_banks_52_wdata_bits = io_banks_52_wdata_bits; // @[FIFO.scala 59:15:@51189.4]
  assign FFRAM_io_banks_53_wdata_valid = io_banks_53_wdata_valid; // @[FIFO.scala 59:15:@51193.4]
  assign FFRAM_io_banks_53_wdata_bits = io_banks_53_wdata_bits; // @[FIFO.scala 59:15:@51192.4]
  assign FFRAM_io_banks_54_wdata_valid = io_banks_54_wdata_valid; // @[FIFO.scala 59:15:@51196.4]
  assign FFRAM_io_banks_54_wdata_bits = io_banks_54_wdata_bits; // @[FIFO.scala 59:15:@51195.4]
  assign FFRAM_io_banks_55_wdata_valid = io_banks_55_wdata_valid; // @[FIFO.scala 59:15:@51199.4]
  assign FFRAM_io_banks_55_wdata_bits = io_banks_55_wdata_bits; // @[FIFO.scala 59:15:@51198.4]
  assign FFRAM_io_banks_56_wdata_valid = io_banks_56_wdata_valid; // @[FIFO.scala 59:15:@51202.4]
  assign FFRAM_io_banks_56_wdata_bits = io_banks_56_wdata_bits; // @[FIFO.scala 59:15:@51201.4]
  assign FFRAM_io_banks_57_wdata_valid = io_banks_57_wdata_valid; // @[FIFO.scala 59:15:@51205.4]
  assign FFRAM_io_banks_57_wdata_bits = io_banks_57_wdata_bits; // @[FIFO.scala 59:15:@51204.4]
  assign FFRAM_io_banks_58_wdata_valid = io_banks_58_wdata_valid; // @[FIFO.scala 59:15:@51208.4]
  assign FFRAM_io_banks_58_wdata_bits = io_banks_58_wdata_bits; // @[FIFO.scala 59:15:@51207.4]
  assign FFRAM_io_banks_59_wdata_valid = io_banks_59_wdata_valid; // @[FIFO.scala 59:15:@51211.4]
  assign FFRAM_io_banks_59_wdata_bits = io_banks_59_wdata_bits; // @[FIFO.scala 59:15:@51210.4]
  assign FFRAM_io_banks_60_wdata_valid = io_banks_60_wdata_valid; // @[FIFO.scala 59:15:@51214.4]
  assign FFRAM_io_banks_60_wdata_bits = io_banks_60_wdata_bits; // @[FIFO.scala 59:15:@51213.4]
  assign FFRAM_io_banks_61_wdata_valid = io_banks_61_wdata_valid; // @[FIFO.scala 59:15:@51217.4]
  assign FFRAM_io_banks_61_wdata_bits = io_banks_61_wdata_bits; // @[FIFO.scala 59:15:@51216.4]
  assign FFRAM_io_banks_62_wdata_valid = io_banks_62_wdata_valid; // @[FIFO.scala 59:15:@51220.4]
  assign FFRAM_io_banks_62_wdata_bits = io_banks_62_wdata_bits; // @[FIFO.scala 59:15:@51219.4]
  assign FFRAM_io_banks_63_wdata_valid = io_banks_63_wdata_valid; // @[FIFO.scala 59:15:@51223.4]
  assign FFRAM_io_banks_63_wdata_bits = io_banks_63_wdata_bits; // @[FIFO.scala 59:15:@51222.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_1657) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module StreamControllerStore( // @[:@52002.2]
  input         clock, // @[:@52003.4]
  input         reset, // @[:@52004.4]
  input         io_dram_cmd_ready, // @[:@52005.4]
  output        io_dram_cmd_valid, // @[:@52005.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@52005.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@52005.4]
  input         io_dram_wdata_ready, // @[:@52005.4]
  output        io_dram_wdata_valid, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@52005.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@52005.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@52005.4]
  output        io_dram_wresp_ready, // @[:@52005.4]
  input         io_dram_wresp_valid, // @[:@52005.4]
  output        io_store_cmd_ready, // @[:@52005.4]
  input         io_store_cmd_valid, // @[:@52005.4]
  input  [63:0] io_store_cmd_bits_addr, // @[:@52005.4]
  input  [31:0] io_store_cmd_bits_size, // @[:@52005.4]
  output        io_store_data_ready, // @[:@52005.4]
  input         io_store_data_valid, // @[:@52005.4]
  input  [31:0] io_store_data_bits_wdata_0, // @[:@52005.4]
  input         io_store_data_bits_wstrb, // @[:@52005.4]
  input         io_store_wresp_ready, // @[:@52005.4]
  output        io_store_wresp_valid, // @[:@52005.4]
  output        io_store_wresp_bits // @[:@52005.4]
);
  wire  cmd_clock; // @[StreamController.scala 75:19:@52130.4]
  wire  cmd_reset; // @[StreamController.scala 75:19:@52130.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 75:19:@52130.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 75:19:@52130.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 75:19:@52130.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 75:19:@52130.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 75:19:@52130.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 75:19:@52130.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 75:19:@52130.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 75:19:@52130.4]
  wire  wdata_clock; // @[StreamController.scala 88:21:@52536.4]
  wire  wdata_reset; // @[StreamController.scala 88:21:@52536.4]
  wire  wdata_io_in_ready; // @[StreamController.scala 88:21:@52536.4]
  wire  wdata_io_in_valid; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_in_bits_data_0; // @[StreamController.scala 88:21:@52536.4]
  wire  wdata_io_in_bits_strobe; // @[StreamController.scala 88:21:@52536.4]
  wire  wdata_io_out_ready; // @[StreamController.scala 88:21:@52536.4]
  wire  wdata_io_out_valid; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_0; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_1; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_2; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_3; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_4; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_5; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_6; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_7; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_8; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_9; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_10; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_11; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_12; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_13; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_14; // @[StreamController.scala 88:21:@52536.4]
  wire [31:0] wdata_io_out_bits_data_15; // @[StreamController.scala 88:21:@52536.4]
  wire [63:0] wdata_io_out_bits_strobe; // @[StreamController.scala 88:21:@52536.4]
  wire  wresp_clock; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_reset; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_in_ready; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_in_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_in_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_out_ready; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_out_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_out_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_0_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_0_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_1_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_1_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_2_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_2_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_3_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_3_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_4_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_4_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_5_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_5_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_6_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_6_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_7_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_7_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_8_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_8_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_9_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_9_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_10_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_10_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_11_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_11_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_12_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_12_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_13_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_13_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_14_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_14_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_15_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_15_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_16_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_16_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_17_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_17_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_18_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_18_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_19_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_19_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_20_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_20_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_21_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_21_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_22_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_22_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_23_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_23_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_24_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_24_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_25_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_25_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_26_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_26_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_27_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_27_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_28_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_28_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_29_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_29_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_30_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_30_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_31_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_31_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_32_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_32_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_33_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_33_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_34_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_34_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_35_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_35_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_36_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_36_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_37_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_37_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_38_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_38_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_39_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_39_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_40_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_40_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_41_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_41_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_42_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_42_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_43_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_43_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_44_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_44_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_45_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_45_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_46_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_46_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_47_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_47_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_48_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_48_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_49_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_49_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_50_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_50_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_51_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_51_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_52_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_52_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_53_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_53_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_54_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_54_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_55_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_55_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_56_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_56_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_57_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_57_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_58_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_58_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_59_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_59_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_60_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_60_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_61_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_61_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_62_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_62_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_63_wdata_valid; // @[StreamController.scala 100:21:@52777.4]
  wire  wresp_io_banks_63_wdata_bits; // @[StreamController.scala 100:21:@52777.4]
  wire [25:0] _T_111; // @[StreamController.scala 21:10:@52533.4]
  FIFO cmd ( // @[StreamController.scala 75:19:@52130.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert wdata ( // @[StreamController.scala 88:21:@52536.4]
    .clock(wdata_clock),
    .reset(wdata_reset),
    .io_in_ready(wdata_io_in_ready),
    .io_in_valid(wdata_io_in_valid),
    .io_in_bits_data_0(wdata_io_in_bits_data_0),
    .io_in_bits_strobe(wdata_io_in_bits_strobe),
    .io_out_ready(wdata_io_out_ready),
    .io_out_valid(wdata_io_out_valid),
    .io_out_bits_data_0(wdata_io_out_bits_data_0),
    .io_out_bits_data_1(wdata_io_out_bits_data_1),
    .io_out_bits_data_2(wdata_io_out_bits_data_2),
    .io_out_bits_data_3(wdata_io_out_bits_data_3),
    .io_out_bits_data_4(wdata_io_out_bits_data_4),
    .io_out_bits_data_5(wdata_io_out_bits_data_5),
    .io_out_bits_data_6(wdata_io_out_bits_data_6),
    .io_out_bits_data_7(wdata_io_out_bits_data_7),
    .io_out_bits_data_8(wdata_io_out_bits_data_8),
    .io_out_bits_data_9(wdata_io_out_bits_data_9),
    .io_out_bits_data_10(wdata_io_out_bits_data_10),
    .io_out_bits_data_11(wdata_io_out_bits_data_11),
    .io_out_bits_data_12(wdata_io_out_bits_data_12),
    .io_out_bits_data_13(wdata_io_out_bits_data_13),
    .io_out_bits_data_14(wdata_io_out_bits_data_14),
    .io_out_bits_data_15(wdata_io_out_bits_data_15),
    .io_out_bits_strobe(wdata_io_out_bits_strobe)
  );
  FIFO_33 wresp ( // @[StreamController.scala 100:21:@52777.4]
    .clock(wresp_clock),
    .reset(wresp_reset),
    .io_in_ready(wresp_io_in_ready),
    .io_in_valid(wresp_io_in_valid),
    .io_in_bits(wresp_io_in_bits),
    .io_out_ready(wresp_io_out_ready),
    .io_out_valid(wresp_io_out_valid),
    .io_out_bits(wresp_io_out_bits),
    .io_banks_0_wdata_valid(wresp_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(wresp_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(wresp_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(wresp_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(wresp_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(wresp_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(wresp_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(wresp_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(wresp_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(wresp_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(wresp_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(wresp_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(wresp_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(wresp_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(wresp_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(wresp_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(wresp_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(wresp_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(wresp_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(wresp_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(wresp_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(wresp_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(wresp_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(wresp_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(wresp_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(wresp_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(wresp_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(wresp_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(wresp_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(wresp_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(wresp_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(wresp_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(wresp_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(wresp_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(wresp_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(wresp_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(wresp_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(wresp_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(wresp_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(wresp_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(wresp_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(wresp_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(wresp_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(wresp_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(wresp_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(wresp_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(wresp_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(wresp_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(wresp_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(wresp_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(wresp_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(wresp_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(wresp_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(wresp_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(wresp_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(wresp_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(wresp_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(wresp_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(wresp_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(wresp_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(wresp_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(wresp_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(wresp_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(wresp_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(wresp_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(wresp_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(wresp_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(wresp_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(wresp_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(wresp_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(wresp_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(wresp_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(wresp_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(wresp_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(wresp_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(wresp_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(wresp_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(wresp_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(wresp_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(wresp_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(wresp_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(wresp_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(wresp_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(wresp_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(wresp_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(wresp_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(wresp_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(wresp_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(wresp_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(wresp_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(wresp_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(wresp_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(wresp_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(wresp_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(wresp_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(wresp_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(wresp_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(wresp_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(wresp_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(wresp_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(wresp_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(wresp_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(wresp_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(wresp_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(wresp_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(wresp_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(wresp_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(wresp_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(wresp_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(wresp_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(wresp_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(wresp_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(wresp_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(wresp_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(wresp_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(wresp_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(wresp_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(wresp_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(wresp_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(wresp_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(wresp_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(wresp_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(wresp_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(wresp_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(wresp_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(wresp_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(wresp_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(wresp_io_banks_63_wdata_bits)
  );
  assign _T_111 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@52533.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 81:21:@52530.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 83:25:@52531.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_111}; // @[StreamController.scala 85:25:@52534.4]
  assign io_dram_wdata_valid = wdata_io_out_valid; // @[StreamController.scala 95:23:@52566.4]
  assign io_dram_wdata_bits_wdata_0 = wdata_io_out_bits_data_0; // @[StreamController.scala 96:28:@52567.4]
  assign io_dram_wdata_bits_wdata_1 = wdata_io_out_bits_data_1; // @[StreamController.scala 96:28:@52568.4]
  assign io_dram_wdata_bits_wdata_2 = wdata_io_out_bits_data_2; // @[StreamController.scala 96:28:@52569.4]
  assign io_dram_wdata_bits_wdata_3 = wdata_io_out_bits_data_3; // @[StreamController.scala 96:28:@52570.4]
  assign io_dram_wdata_bits_wdata_4 = wdata_io_out_bits_data_4; // @[StreamController.scala 96:28:@52571.4]
  assign io_dram_wdata_bits_wdata_5 = wdata_io_out_bits_data_5; // @[StreamController.scala 96:28:@52572.4]
  assign io_dram_wdata_bits_wdata_6 = wdata_io_out_bits_data_6; // @[StreamController.scala 96:28:@52573.4]
  assign io_dram_wdata_bits_wdata_7 = wdata_io_out_bits_data_7; // @[StreamController.scala 96:28:@52574.4]
  assign io_dram_wdata_bits_wdata_8 = wdata_io_out_bits_data_8; // @[StreamController.scala 96:28:@52575.4]
  assign io_dram_wdata_bits_wdata_9 = wdata_io_out_bits_data_9; // @[StreamController.scala 96:28:@52576.4]
  assign io_dram_wdata_bits_wdata_10 = wdata_io_out_bits_data_10; // @[StreamController.scala 96:28:@52577.4]
  assign io_dram_wdata_bits_wdata_11 = wdata_io_out_bits_data_11; // @[StreamController.scala 96:28:@52578.4]
  assign io_dram_wdata_bits_wdata_12 = wdata_io_out_bits_data_12; // @[StreamController.scala 96:28:@52579.4]
  assign io_dram_wdata_bits_wdata_13 = wdata_io_out_bits_data_13; // @[StreamController.scala 96:28:@52580.4]
  assign io_dram_wdata_bits_wdata_14 = wdata_io_out_bits_data_14; // @[StreamController.scala 96:28:@52581.4]
  assign io_dram_wdata_bits_wdata_15 = wdata_io_out_bits_data_15; // @[StreamController.scala 96:28:@52582.4]
  assign io_dram_wdata_bits_wstrb_0 = wdata_io_out_bits_strobe[63]; // @[StreamController.scala 97:28:@52712.4]
  assign io_dram_wdata_bits_wstrb_1 = wdata_io_out_bits_strobe[62]; // @[StreamController.scala 97:28:@52713.4]
  assign io_dram_wdata_bits_wstrb_2 = wdata_io_out_bits_strobe[61]; // @[StreamController.scala 97:28:@52714.4]
  assign io_dram_wdata_bits_wstrb_3 = wdata_io_out_bits_strobe[60]; // @[StreamController.scala 97:28:@52715.4]
  assign io_dram_wdata_bits_wstrb_4 = wdata_io_out_bits_strobe[59]; // @[StreamController.scala 97:28:@52716.4]
  assign io_dram_wdata_bits_wstrb_5 = wdata_io_out_bits_strobe[58]; // @[StreamController.scala 97:28:@52717.4]
  assign io_dram_wdata_bits_wstrb_6 = wdata_io_out_bits_strobe[57]; // @[StreamController.scala 97:28:@52718.4]
  assign io_dram_wdata_bits_wstrb_7 = wdata_io_out_bits_strobe[56]; // @[StreamController.scala 97:28:@52719.4]
  assign io_dram_wdata_bits_wstrb_8 = wdata_io_out_bits_strobe[55]; // @[StreamController.scala 97:28:@52720.4]
  assign io_dram_wdata_bits_wstrb_9 = wdata_io_out_bits_strobe[54]; // @[StreamController.scala 97:28:@52721.4]
  assign io_dram_wdata_bits_wstrb_10 = wdata_io_out_bits_strobe[53]; // @[StreamController.scala 97:28:@52722.4]
  assign io_dram_wdata_bits_wstrb_11 = wdata_io_out_bits_strobe[52]; // @[StreamController.scala 97:28:@52723.4]
  assign io_dram_wdata_bits_wstrb_12 = wdata_io_out_bits_strobe[51]; // @[StreamController.scala 97:28:@52724.4]
  assign io_dram_wdata_bits_wstrb_13 = wdata_io_out_bits_strobe[50]; // @[StreamController.scala 97:28:@52725.4]
  assign io_dram_wdata_bits_wstrb_14 = wdata_io_out_bits_strobe[49]; // @[StreamController.scala 97:28:@52726.4]
  assign io_dram_wdata_bits_wstrb_15 = wdata_io_out_bits_strobe[48]; // @[StreamController.scala 97:28:@52727.4]
  assign io_dram_wdata_bits_wstrb_16 = wdata_io_out_bits_strobe[47]; // @[StreamController.scala 97:28:@52728.4]
  assign io_dram_wdata_bits_wstrb_17 = wdata_io_out_bits_strobe[46]; // @[StreamController.scala 97:28:@52729.4]
  assign io_dram_wdata_bits_wstrb_18 = wdata_io_out_bits_strobe[45]; // @[StreamController.scala 97:28:@52730.4]
  assign io_dram_wdata_bits_wstrb_19 = wdata_io_out_bits_strobe[44]; // @[StreamController.scala 97:28:@52731.4]
  assign io_dram_wdata_bits_wstrb_20 = wdata_io_out_bits_strobe[43]; // @[StreamController.scala 97:28:@52732.4]
  assign io_dram_wdata_bits_wstrb_21 = wdata_io_out_bits_strobe[42]; // @[StreamController.scala 97:28:@52733.4]
  assign io_dram_wdata_bits_wstrb_22 = wdata_io_out_bits_strobe[41]; // @[StreamController.scala 97:28:@52734.4]
  assign io_dram_wdata_bits_wstrb_23 = wdata_io_out_bits_strobe[40]; // @[StreamController.scala 97:28:@52735.4]
  assign io_dram_wdata_bits_wstrb_24 = wdata_io_out_bits_strobe[39]; // @[StreamController.scala 97:28:@52736.4]
  assign io_dram_wdata_bits_wstrb_25 = wdata_io_out_bits_strobe[38]; // @[StreamController.scala 97:28:@52737.4]
  assign io_dram_wdata_bits_wstrb_26 = wdata_io_out_bits_strobe[37]; // @[StreamController.scala 97:28:@52738.4]
  assign io_dram_wdata_bits_wstrb_27 = wdata_io_out_bits_strobe[36]; // @[StreamController.scala 97:28:@52739.4]
  assign io_dram_wdata_bits_wstrb_28 = wdata_io_out_bits_strobe[35]; // @[StreamController.scala 97:28:@52740.4]
  assign io_dram_wdata_bits_wstrb_29 = wdata_io_out_bits_strobe[34]; // @[StreamController.scala 97:28:@52741.4]
  assign io_dram_wdata_bits_wstrb_30 = wdata_io_out_bits_strobe[33]; // @[StreamController.scala 97:28:@52742.4]
  assign io_dram_wdata_bits_wstrb_31 = wdata_io_out_bits_strobe[32]; // @[StreamController.scala 97:28:@52743.4]
  assign io_dram_wdata_bits_wstrb_32 = wdata_io_out_bits_strobe[31]; // @[StreamController.scala 97:28:@52744.4]
  assign io_dram_wdata_bits_wstrb_33 = wdata_io_out_bits_strobe[30]; // @[StreamController.scala 97:28:@52745.4]
  assign io_dram_wdata_bits_wstrb_34 = wdata_io_out_bits_strobe[29]; // @[StreamController.scala 97:28:@52746.4]
  assign io_dram_wdata_bits_wstrb_35 = wdata_io_out_bits_strobe[28]; // @[StreamController.scala 97:28:@52747.4]
  assign io_dram_wdata_bits_wstrb_36 = wdata_io_out_bits_strobe[27]; // @[StreamController.scala 97:28:@52748.4]
  assign io_dram_wdata_bits_wstrb_37 = wdata_io_out_bits_strobe[26]; // @[StreamController.scala 97:28:@52749.4]
  assign io_dram_wdata_bits_wstrb_38 = wdata_io_out_bits_strobe[25]; // @[StreamController.scala 97:28:@52750.4]
  assign io_dram_wdata_bits_wstrb_39 = wdata_io_out_bits_strobe[24]; // @[StreamController.scala 97:28:@52751.4]
  assign io_dram_wdata_bits_wstrb_40 = wdata_io_out_bits_strobe[23]; // @[StreamController.scala 97:28:@52752.4]
  assign io_dram_wdata_bits_wstrb_41 = wdata_io_out_bits_strobe[22]; // @[StreamController.scala 97:28:@52753.4]
  assign io_dram_wdata_bits_wstrb_42 = wdata_io_out_bits_strobe[21]; // @[StreamController.scala 97:28:@52754.4]
  assign io_dram_wdata_bits_wstrb_43 = wdata_io_out_bits_strobe[20]; // @[StreamController.scala 97:28:@52755.4]
  assign io_dram_wdata_bits_wstrb_44 = wdata_io_out_bits_strobe[19]; // @[StreamController.scala 97:28:@52756.4]
  assign io_dram_wdata_bits_wstrb_45 = wdata_io_out_bits_strobe[18]; // @[StreamController.scala 97:28:@52757.4]
  assign io_dram_wdata_bits_wstrb_46 = wdata_io_out_bits_strobe[17]; // @[StreamController.scala 97:28:@52758.4]
  assign io_dram_wdata_bits_wstrb_47 = wdata_io_out_bits_strobe[16]; // @[StreamController.scala 97:28:@52759.4]
  assign io_dram_wdata_bits_wstrb_48 = wdata_io_out_bits_strobe[15]; // @[StreamController.scala 97:28:@52760.4]
  assign io_dram_wdata_bits_wstrb_49 = wdata_io_out_bits_strobe[14]; // @[StreamController.scala 97:28:@52761.4]
  assign io_dram_wdata_bits_wstrb_50 = wdata_io_out_bits_strobe[13]; // @[StreamController.scala 97:28:@52762.4]
  assign io_dram_wdata_bits_wstrb_51 = wdata_io_out_bits_strobe[12]; // @[StreamController.scala 97:28:@52763.4]
  assign io_dram_wdata_bits_wstrb_52 = wdata_io_out_bits_strobe[11]; // @[StreamController.scala 97:28:@52764.4]
  assign io_dram_wdata_bits_wstrb_53 = wdata_io_out_bits_strobe[10]; // @[StreamController.scala 97:28:@52765.4]
  assign io_dram_wdata_bits_wstrb_54 = wdata_io_out_bits_strobe[9]; // @[StreamController.scala 97:28:@52766.4]
  assign io_dram_wdata_bits_wstrb_55 = wdata_io_out_bits_strobe[8]; // @[StreamController.scala 97:28:@52767.4]
  assign io_dram_wdata_bits_wstrb_56 = wdata_io_out_bits_strobe[7]; // @[StreamController.scala 97:28:@52768.4]
  assign io_dram_wdata_bits_wstrb_57 = wdata_io_out_bits_strobe[6]; // @[StreamController.scala 97:28:@52769.4]
  assign io_dram_wdata_bits_wstrb_58 = wdata_io_out_bits_strobe[5]; // @[StreamController.scala 97:28:@52770.4]
  assign io_dram_wdata_bits_wstrb_59 = wdata_io_out_bits_strobe[4]; // @[StreamController.scala 97:28:@52771.4]
  assign io_dram_wdata_bits_wstrb_60 = wdata_io_out_bits_strobe[3]; // @[StreamController.scala 97:28:@52772.4]
  assign io_dram_wdata_bits_wstrb_61 = wdata_io_out_bits_strobe[2]; // @[StreamController.scala 97:28:@52773.4]
  assign io_dram_wdata_bits_wstrb_62 = wdata_io_out_bits_strobe[1]; // @[StreamController.scala 97:28:@52774.4]
  assign io_dram_wdata_bits_wstrb_63 = wdata_io_out_bits_strobe[0]; // @[StreamController.scala 97:28:@52775.4]
  assign io_dram_wresp_ready = wresp_io_in_ready; // @[StreamController.scala 104:23:@53044.4]
  assign io_store_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 79:22:@52528.4]
  assign io_store_data_ready = wdata_io_in_ready; // @[StreamController.scala 93:23:@52565.4]
  assign io_store_wresp_valid = wresp_io_out_valid; // @[StreamController.scala 106:24:@53045.4]
  assign io_store_wresp_bits = wresp_io_out_bits; // @[StreamController.scala 107:23:@53046.4]
  assign cmd_clock = clock; // @[:@52131.4]
  assign cmd_reset = reset; // @[:@52132.4]
  assign cmd_io_in_valid = io_store_cmd_valid; // @[StreamController.scala 77:19:@52525.4]
  assign cmd_io_in_bits_addr = io_store_cmd_bits_addr; // @[StreamController.scala 78:18:@52527.4]
  assign cmd_io_in_bits_size = io_store_cmd_bits_size; // @[StreamController.scala 78:18:@52526.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 80:20:@52529.4]
  assign wdata_clock = clock; // @[:@52537.4]
  assign wdata_reset = reset; // @[:@52538.4]
  assign wdata_io_in_valid = io_store_data_valid; // @[StreamController.scala 90:21:@52562.4]
  assign wdata_io_in_bits_data_0 = io_store_data_bits_wdata_0; // @[StreamController.scala 91:25:@52563.4]
  assign wdata_io_in_bits_strobe = io_store_data_bits_wstrb; // @[StreamController.scala 92:27:@52564.4]
  assign wdata_io_out_ready = io_dram_wdata_ready; // @[StreamController.scala 98:22:@52776.4]
  assign wresp_clock = clock; // @[:@52778.4]
  assign wresp_reset = reset; // @[:@52779.4]
  assign wresp_io_in_valid = io_dram_wresp_valid; // @[StreamController.scala 102:21:@53042.4]
  assign wresp_io_in_bits = 1'h1; // @[StreamController.scala 103:20:@53043.4]
  assign wresp_io_out_ready = io_store_wresp_ready; // @[StreamController.scala 108:22:@53047.4]
  assign wresp_io_banks_0_wdata_valid = 1'h0;
  assign wresp_io_banks_0_wdata_bits = 1'h0;
  assign wresp_io_banks_1_wdata_valid = 1'h0;
  assign wresp_io_banks_1_wdata_bits = 1'h0;
  assign wresp_io_banks_2_wdata_valid = 1'h0;
  assign wresp_io_banks_2_wdata_bits = 1'h0;
  assign wresp_io_banks_3_wdata_valid = 1'h0;
  assign wresp_io_banks_3_wdata_bits = 1'h0;
  assign wresp_io_banks_4_wdata_valid = 1'h0;
  assign wresp_io_banks_4_wdata_bits = 1'h0;
  assign wresp_io_banks_5_wdata_valid = 1'h0;
  assign wresp_io_banks_5_wdata_bits = 1'h0;
  assign wresp_io_banks_6_wdata_valid = 1'h0;
  assign wresp_io_banks_6_wdata_bits = 1'h0;
  assign wresp_io_banks_7_wdata_valid = 1'h0;
  assign wresp_io_banks_7_wdata_bits = 1'h0;
  assign wresp_io_banks_8_wdata_valid = 1'h0;
  assign wresp_io_banks_8_wdata_bits = 1'h0;
  assign wresp_io_banks_9_wdata_valid = 1'h0;
  assign wresp_io_banks_9_wdata_bits = 1'h0;
  assign wresp_io_banks_10_wdata_valid = 1'h0;
  assign wresp_io_banks_10_wdata_bits = 1'h0;
  assign wresp_io_banks_11_wdata_valid = 1'h0;
  assign wresp_io_banks_11_wdata_bits = 1'h0;
  assign wresp_io_banks_12_wdata_valid = 1'h0;
  assign wresp_io_banks_12_wdata_bits = 1'h0;
  assign wresp_io_banks_13_wdata_valid = 1'h0;
  assign wresp_io_banks_13_wdata_bits = 1'h0;
  assign wresp_io_banks_14_wdata_valid = 1'h0;
  assign wresp_io_banks_14_wdata_bits = 1'h0;
  assign wresp_io_banks_15_wdata_valid = 1'h0;
  assign wresp_io_banks_15_wdata_bits = 1'h0;
  assign wresp_io_banks_16_wdata_valid = 1'h0;
  assign wresp_io_banks_16_wdata_bits = 1'h0;
  assign wresp_io_banks_17_wdata_valid = 1'h0;
  assign wresp_io_banks_17_wdata_bits = 1'h0;
  assign wresp_io_banks_18_wdata_valid = 1'h0;
  assign wresp_io_banks_18_wdata_bits = 1'h0;
  assign wresp_io_banks_19_wdata_valid = 1'h0;
  assign wresp_io_banks_19_wdata_bits = 1'h0;
  assign wresp_io_banks_20_wdata_valid = 1'h0;
  assign wresp_io_banks_20_wdata_bits = 1'h0;
  assign wresp_io_banks_21_wdata_valid = 1'h0;
  assign wresp_io_banks_21_wdata_bits = 1'h0;
  assign wresp_io_banks_22_wdata_valid = 1'h0;
  assign wresp_io_banks_22_wdata_bits = 1'h0;
  assign wresp_io_banks_23_wdata_valid = 1'h0;
  assign wresp_io_banks_23_wdata_bits = 1'h0;
  assign wresp_io_banks_24_wdata_valid = 1'h0;
  assign wresp_io_banks_24_wdata_bits = 1'h0;
  assign wresp_io_banks_25_wdata_valid = 1'h0;
  assign wresp_io_banks_25_wdata_bits = 1'h0;
  assign wresp_io_banks_26_wdata_valid = 1'h0;
  assign wresp_io_banks_26_wdata_bits = 1'h0;
  assign wresp_io_banks_27_wdata_valid = 1'h0;
  assign wresp_io_banks_27_wdata_bits = 1'h0;
  assign wresp_io_banks_28_wdata_valid = 1'h0;
  assign wresp_io_banks_28_wdata_bits = 1'h0;
  assign wresp_io_banks_29_wdata_valid = 1'h0;
  assign wresp_io_banks_29_wdata_bits = 1'h0;
  assign wresp_io_banks_30_wdata_valid = 1'h0;
  assign wresp_io_banks_30_wdata_bits = 1'h0;
  assign wresp_io_banks_31_wdata_valid = 1'h0;
  assign wresp_io_banks_31_wdata_bits = 1'h0;
  assign wresp_io_banks_32_wdata_valid = 1'h0;
  assign wresp_io_banks_32_wdata_bits = 1'h0;
  assign wresp_io_banks_33_wdata_valid = 1'h0;
  assign wresp_io_banks_33_wdata_bits = 1'h0;
  assign wresp_io_banks_34_wdata_valid = 1'h0;
  assign wresp_io_banks_34_wdata_bits = 1'h0;
  assign wresp_io_banks_35_wdata_valid = 1'h0;
  assign wresp_io_banks_35_wdata_bits = 1'h0;
  assign wresp_io_banks_36_wdata_valid = 1'h0;
  assign wresp_io_banks_36_wdata_bits = 1'h0;
  assign wresp_io_banks_37_wdata_valid = 1'h0;
  assign wresp_io_banks_37_wdata_bits = 1'h0;
  assign wresp_io_banks_38_wdata_valid = 1'h0;
  assign wresp_io_banks_38_wdata_bits = 1'h0;
  assign wresp_io_banks_39_wdata_valid = 1'h0;
  assign wresp_io_banks_39_wdata_bits = 1'h0;
  assign wresp_io_banks_40_wdata_valid = 1'h0;
  assign wresp_io_banks_40_wdata_bits = 1'h0;
  assign wresp_io_banks_41_wdata_valid = 1'h0;
  assign wresp_io_banks_41_wdata_bits = 1'h0;
  assign wresp_io_banks_42_wdata_valid = 1'h0;
  assign wresp_io_banks_42_wdata_bits = 1'h0;
  assign wresp_io_banks_43_wdata_valid = 1'h0;
  assign wresp_io_banks_43_wdata_bits = 1'h0;
  assign wresp_io_banks_44_wdata_valid = 1'h0;
  assign wresp_io_banks_44_wdata_bits = 1'h0;
  assign wresp_io_banks_45_wdata_valid = 1'h0;
  assign wresp_io_banks_45_wdata_bits = 1'h0;
  assign wresp_io_banks_46_wdata_valid = 1'h0;
  assign wresp_io_banks_46_wdata_bits = 1'h0;
  assign wresp_io_banks_47_wdata_valid = 1'h0;
  assign wresp_io_banks_47_wdata_bits = 1'h0;
  assign wresp_io_banks_48_wdata_valid = 1'h0;
  assign wresp_io_banks_48_wdata_bits = 1'h0;
  assign wresp_io_banks_49_wdata_valid = 1'h0;
  assign wresp_io_banks_49_wdata_bits = 1'h0;
  assign wresp_io_banks_50_wdata_valid = 1'h0;
  assign wresp_io_banks_50_wdata_bits = 1'h0;
  assign wresp_io_banks_51_wdata_valid = 1'h0;
  assign wresp_io_banks_51_wdata_bits = 1'h0;
  assign wresp_io_banks_52_wdata_valid = 1'h0;
  assign wresp_io_banks_52_wdata_bits = 1'h0;
  assign wresp_io_banks_53_wdata_valid = 1'h0;
  assign wresp_io_banks_53_wdata_bits = 1'h0;
  assign wresp_io_banks_54_wdata_valid = 1'h0;
  assign wresp_io_banks_54_wdata_bits = 1'h0;
  assign wresp_io_banks_55_wdata_valid = 1'h0;
  assign wresp_io_banks_55_wdata_bits = 1'h0;
  assign wresp_io_banks_56_wdata_valid = 1'h0;
  assign wresp_io_banks_56_wdata_bits = 1'h0;
  assign wresp_io_banks_57_wdata_valid = 1'h0;
  assign wresp_io_banks_57_wdata_bits = 1'h0;
  assign wresp_io_banks_58_wdata_valid = 1'h0;
  assign wresp_io_banks_58_wdata_bits = 1'h0;
  assign wresp_io_banks_59_wdata_valid = 1'h0;
  assign wresp_io_banks_59_wdata_bits = 1'h0;
  assign wresp_io_banks_60_wdata_valid = 1'h0;
  assign wresp_io_banks_60_wdata_bits = 1'h0;
  assign wresp_io_banks_61_wdata_valid = 1'h0;
  assign wresp_io_banks_61_wdata_bits = 1'h0;
  assign wresp_io_banks_62_wdata_valid = 1'h0;
  assign wresp_io_banks_62_wdata_bits = 1'h0;
  assign wresp_io_banks_63_wdata_valid = 1'h0;
  assign wresp_io_banks_63_wdata_bits = 1'h0;
endmodule
module MuxPipe( // @[:@53113.2]
  output        io_in_ready, // @[:@53116.4]
  input         io_in_valid, // @[:@53116.4]
  input  [63:0] io_in_bits_0_addr, // @[:@53116.4]
  input  [31:0] io_in_bits_0_size, // @[:@53116.4]
  input         io_in_bits_0_isWr, // @[:@53116.4]
  input  [31:0] io_in_bits_0_tag, // @[:@53116.4]
  input         io_out_ready, // @[:@53116.4]
  output        io_out_valid, // @[:@53116.4]
  output [63:0] io_out_bits_addr, // @[:@53116.4]
  output [31:0] io_out_bits_size, // @[:@53116.4]
  output        io_out_bits_isWr, // @[:@53116.4]
  output [31:0] io_out_bits_tag // @[:@53116.4]
);
  wire  _T_42; // @[MuxN.scala 28:31:@53118.4]
  assign _T_42 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@53118.4]
  assign io_in_ready = io_out_ready | _T_42; // @[MuxN.scala 71:15:@53127.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@53126.4]
  assign io_out_bits_addr = io_in_bits_0_addr; // @[MuxN.scala 72:15:@53132.4]
  assign io_out_bits_size = io_in_bits_0_size; // @[MuxN.scala 72:15:@53131.4]
  assign io_out_bits_isWr = io_in_bits_0_isWr; // @[MuxN.scala 72:15:@53129.4]
  assign io_out_bits_tag = io_in_bits_0_tag; // @[MuxN.scala 72:15:@53128.4]
endmodule
module MuxPipe_1( // @[:@53134.2]
  output        io_in_ready, // @[:@53137.4]
  input         io_in_valid, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_0, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_1, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_2, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_3, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_4, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_5, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_6, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_7, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_8, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_9, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_10, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_11, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_12, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_13, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_14, // @[:@53137.4]
  input  [31:0] io_in_bits_0_wdata_15, // @[:@53137.4]
  input         io_in_bits_0_wstrb_0, // @[:@53137.4]
  input         io_in_bits_0_wstrb_1, // @[:@53137.4]
  input         io_in_bits_0_wstrb_2, // @[:@53137.4]
  input         io_in_bits_0_wstrb_3, // @[:@53137.4]
  input         io_in_bits_0_wstrb_4, // @[:@53137.4]
  input         io_in_bits_0_wstrb_5, // @[:@53137.4]
  input         io_in_bits_0_wstrb_6, // @[:@53137.4]
  input         io_in_bits_0_wstrb_7, // @[:@53137.4]
  input         io_in_bits_0_wstrb_8, // @[:@53137.4]
  input         io_in_bits_0_wstrb_9, // @[:@53137.4]
  input         io_in_bits_0_wstrb_10, // @[:@53137.4]
  input         io_in_bits_0_wstrb_11, // @[:@53137.4]
  input         io_in_bits_0_wstrb_12, // @[:@53137.4]
  input         io_in_bits_0_wstrb_13, // @[:@53137.4]
  input         io_in_bits_0_wstrb_14, // @[:@53137.4]
  input         io_in_bits_0_wstrb_15, // @[:@53137.4]
  input         io_in_bits_0_wstrb_16, // @[:@53137.4]
  input         io_in_bits_0_wstrb_17, // @[:@53137.4]
  input         io_in_bits_0_wstrb_18, // @[:@53137.4]
  input         io_in_bits_0_wstrb_19, // @[:@53137.4]
  input         io_in_bits_0_wstrb_20, // @[:@53137.4]
  input         io_in_bits_0_wstrb_21, // @[:@53137.4]
  input         io_in_bits_0_wstrb_22, // @[:@53137.4]
  input         io_in_bits_0_wstrb_23, // @[:@53137.4]
  input         io_in_bits_0_wstrb_24, // @[:@53137.4]
  input         io_in_bits_0_wstrb_25, // @[:@53137.4]
  input         io_in_bits_0_wstrb_26, // @[:@53137.4]
  input         io_in_bits_0_wstrb_27, // @[:@53137.4]
  input         io_in_bits_0_wstrb_28, // @[:@53137.4]
  input         io_in_bits_0_wstrb_29, // @[:@53137.4]
  input         io_in_bits_0_wstrb_30, // @[:@53137.4]
  input         io_in_bits_0_wstrb_31, // @[:@53137.4]
  input         io_in_bits_0_wstrb_32, // @[:@53137.4]
  input         io_in_bits_0_wstrb_33, // @[:@53137.4]
  input         io_in_bits_0_wstrb_34, // @[:@53137.4]
  input         io_in_bits_0_wstrb_35, // @[:@53137.4]
  input         io_in_bits_0_wstrb_36, // @[:@53137.4]
  input         io_in_bits_0_wstrb_37, // @[:@53137.4]
  input         io_in_bits_0_wstrb_38, // @[:@53137.4]
  input         io_in_bits_0_wstrb_39, // @[:@53137.4]
  input         io_in_bits_0_wstrb_40, // @[:@53137.4]
  input         io_in_bits_0_wstrb_41, // @[:@53137.4]
  input         io_in_bits_0_wstrb_42, // @[:@53137.4]
  input         io_in_bits_0_wstrb_43, // @[:@53137.4]
  input         io_in_bits_0_wstrb_44, // @[:@53137.4]
  input         io_in_bits_0_wstrb_45, // @[:@53137.4]
  input         io_in_bits_0_wstrb_46, // @[:@53137.4]
  input         io_in_bits_0_wstrb_47, // @[:@53137.4]
  input         io_in_bits_0_wstrb_48, // @[:@53137.4]
  input         io_in_bits_0_wstrb_49, // @[:@53137.4]
  input         io_in_bits_0_wstrb_50, // @[:@53137.4]
  input         io_in_bits_0_wstrb_51, // @[:@53137.4]
  input         io_in_bits_0_wstrb_52, // @[:@53137.4]
  input         io_in_bits_0_wstrb_53, // @[:@53137.4]
  input         io_in_bits_0_wstrb_54, // @[:@53137.4]
  input         io_in_bits_0_wstrb_55, // @[:@53137.4]
  input         io_in_bits_0_wstrb_56, // @[:@53137.4]
  input         io_in_bits_0_wstrb_57, // @[:@53137.4]
  input         io_in_bits_0_wstrb_58, // @[:@53137.4]
  input         io_in_bits_0_wstrb_59, // @[:@53137.4]
  input         io_in_bits_0_wstrb_60, // @[:@53137.4]
  input         io_in_bits_0_wstrb_61, // @[:@53137.4]
  input         io_in_bits_0_wstrb_62, // @[:@53137.4]
  input         io_in_bits_0_wstrb_63, // @[:@53137.4]
  input         io_out_ready, // @[:@53137.4]
  output        io_out_valid, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_0, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_1, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_2, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_3, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_4, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_5, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_6, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_7, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_8, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_9, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_10, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_11, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_12, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_13, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_14, // @[:@53137.4]
  output [31:0] io_out_bits_wdata_15, // @[:@53137.4]
  output        io_out_bits_wstrb_0, // @[:@53137.4]
  output        io_out_bits_wstrb_1, // @[:@53137.4]
  output        io_out_bits_wstrb_2, // @[:@53137.4]
  output        io_out_bits_wstrb_3, // @[:@53137.4]
  output        io_out_bits_wstrb_4, // @[:@53137.4]
  output        io_out_bits_wstrb_5, // @[:@53137.4]
  output        io_out_bits_wstrb_6, // @[:@53137.4]
  output        io_out_bits_wstrb_7, // @[:@53137.4]
  output        io_out_bits_wstrb_8, // @[:@53137.4]
  output        io_out_bits_wstrb_9, // @[:@53137.4]
  output        io_out_bits_wstrb_10, // @[:@53137.4]
  output        io_out_bits_wstrb_11, // @[:@53137.4]
  output        io_out_bits_wstrb_12, // @[:@53137.4]
  output        io_out_bits_wstrb_13, // @[:@53137.4]
  output        io_out_bits_wstrb_14, // @[:@53137.4]
  output        io_out_bits_wstrb_15, // @[:@53137.4]
  output        io_out_bits_wstrb_16, // @[:@53137.4]
  output        io_out_bits_wstrb_17, // @[:@53137.4]
  output        io_out_bits_wstrb_18, // @[:@53137.4]
  output        io_out_bits_wstrb_19, // @[:@53137.4]
  output        io_out_bits_wstrb_20, // @[:@53137.4]
  output        io_out_bits_wstrb_21, // @[:@53137.4]
  output        io_out_bits_wstrb_22, // @[:@53137.4]
  output        io_out_bits_wstrb_23, // @[:@53137.4]
  output        io_out_bits_wstrb_24, // @[:@53137.4]
  output        io_out_bits_wstrb_25, // @[:@53137.4]
  output        io_out_bits_wstrb_26, // @[:@53137.4]
  output        io_out_bits_wstrb_27, // @[:@53137.4]
  output        io_out_bits_wstrb_28, // @[:@53137.4]
  output        io_out_bits_wstrb_29, // @[:@53137.4]
  output        io_out_bits_wstrb_30, // @[:@53137.4]
  output        io_out_bits_wstrb_31, // @[:@53137.4]
  output        io_out_bits_wstrb_32, // @[:@53137.4]
  output        io_out_bits_wstrb_33, // @[:@53137.4]
  output        io_out_bits_wstrb_34, // @[:@53137.4]
  output        io_out_bits_wstrb_35, // @[:@53137.4]
  output        io_out_bits_wstrb_36, // @[:@53137.4]
  output        io_out_bits_wstrb_37, // @[:@53137.4]
  output        io_out_bits_wstrb_38, // @[:@53137.4]
  output        io_out_bits_wstrb_39, // @[:@53137.4]
  output        io_out_bits_wstrb_40, // @[:@53137.4]
  output        io_out_bits_wstrb_41, // @[:@53137.4]
  output        io_out_bits_wstrb_42, // @[:@53137.4]
  output        io_out_bits_wstrb_43, // @[:@53137.4]
  output        io_out_bits_wstrb_44, // @[:@53137.4]
  output        io_out_bits_wstrb_45, // @[:@53137.4]
  output        io_out_bits_wstrb_46, // @[:@53137.4]
  output        io_out_bits_wstrb_47, // @[:@53137.4]
  output        io_out_bits_wstrb_48, // @[:@53137.4]
  output        io_out_bits_wstrb_49, // @[:@53137.4]
  output        io_out_bits_wstrb_50, // @[:@53137.4]
  output        io_out_bits_wstrb_51, // @[:@53137.4]
  output        io_out_bits_wstrb_52, // @[:@53137.4]
  output        io_out_bits_wstrb_53, // @[:@53137.4]
  output        io_out_bits_wstrb_54, // @[:@53137.4]
  output        io_out_bits_wstrb_55, // @[:@53137.4]
  output        io_out_bits_wstrb_56, // @[:@53137.4]
  output        io_out_bits_wstrb_57, // @[:@53137.4]
  output        io_out_bits_wstrb_58, // @[:@53137.4]
  output        io_out_bits_wstrb_59, // @[:@53137.4]
  output        io_out_bits_wstrb_60, // @[:@53137.4]
  output        io_out_bits_wstrb_61, // @[:@53137.4]
  output        io_out_bits_wstrb_62, // @[:@53137.4]
  output        io_out_bits_wstrb_63 // @[:@53137.4]
);
  wire  _T_146; // @[MuxN.scala 28:31:@53139.4]
  assign _T_146 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@53139.4]
  assign io_in_ready = io_out_ready | _T_146; // @[MuxN.scala 71:15:@53224.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@53223.4]
  assign io_out_bits_wdata_0 = io_in_bits_0_wdata_0; // @[MuxN.scala 72:15:@53290.4]
  assign io_out_bits_wdata_1 = io_in_bits_0_wdata_1; // @[MuxN.scala 72:15:@53291.4]
  assign io_out_bits_wdata_2 = io_in_bits_0_wdata_2; // @[MuxN.scala 72:15:@53292.4]
  assign io_out_bits_wdata_3 = io_in_bits_0_wdata_3; // @[MuxN.scala 72:15:@53293.4]
  assign io_out_bits_wdata_4 = io_in_bits_0_wdata_4; // @[MuxN.scala 72:15:@53294.4]
  assign io_out_bits_wdata_5 = io_in_bits_0_wdata_5; // @[MuxN.scala 72:15:@53295.4]
  assign io_out_bits_wdata_6 = io_in_bits_0_wdata_6; // @[MuxN.scala 72:15:@53296.4]
  assign io_out_bits_wdata_7 = io_in_bits_0_wdata_7; // @[MuxN.scala 72:15:@53297.4]
  assign io_out_bits_wdata_8 = io_in_bits_0_wdata_8; // @[MuxN.scala 72:15:@53298.4]
  assign io_out_bits_wdata_9 = io_in_bits_0_wdata_9; // @[MuxN.scala 72:15:@53299.4]
  assign io_out_bits_wdata_10 = io_in_bits_0_wdata_10; // @[MuxN.scala 72:15:@53300.4]
  assign io_out_bits_wdata_11 = io_in_bits_0_wdata_11; // @[MuxN.scala 72:15:@53301.4]
  assign io_out_bits_wdata_12 = io_in_bits_0_wdata_12; // @[MuxN.scala 72:15:@53302.4]
  assign io_out_bits_wdata_13 = io_in_bits_0_wdata_13; // @[MuxN.scala 72:15:@53303.4]
  assign io_out_bits_wdata_14 = io_in_bits_0_wdata_14; // @[MuxN.scala 72:15:@53304.4]
  assign io_out_bits_wdata_15 = io_in_bits_0_wdata_15; // @[MuxN.scala 72:15:@53305.4]
  assign io_out_bits_wstrb_0 = io_in_bits_0_wstrb_0; // @[MuxN.scala 72:15:@53226.4]
  assign io_out_bits_wstrb_1 = io_in_bits_0_wstrb_1; // @[MuxN.scala 72:15:@53227.4]
  assign io_out_bits_wstrb_2 = io_in_bits_0_wstrb_2; // @[MuxN.scala 72:15:@53228.4]
  assign io_out_bits_wstrb_3 = io_in_bits_0_wstrb_3; // @[MuxN.scala 72:15:@53229.4]
  assign io_out_bits_wstrb_4 = io_in_bits_0_wstrb_4; // @[MuxN.scala 72:15:@53230.4]
  assign io_out_bits_wstrb_5 = io_in_bits_0_wstrb_5; // @[MuxN.scala 72:15:@53231.4]
  assign io_out_bits_wstrb_6 = io_in_bits_0_wstrb_6; // @[MuxN.scala 72:15:@53232.4]
  assign io_out_bits_wstrb_7 = io_in_bits_0_wstrb_7; // @[MuxN.scala 72:15:@53233.4]
  assign io_out_bits_wstrb_8 = io_in_bits_0_wstrb_8; // @[MuxN.scala 72:15:@53234.4]
  assign io_out_bits_wstrb_9 = io_in_bits_0_wstrb_9; // @[MuxN.scala 72:15:@53235.4]
  assign io_out_bits_wstrb_10 = io_in_bits_0_wstrb_10; // @[MuxN.scala 72:15:@53236.4]
  assign io_out_bits_wstrb_11 = io_in_bits_0_wstrb_11; // @[MuxN.scala 72:15:@53237.4]
  assign io_out_bits_wstrb_12 = io_in_bits_0_wstrb_12; // @[MuxN.scala 72:15:@53238.4]
  assign io_out_bits_wstrb_13 = io_in_bits_0_wstrb_13; // @[MuxN.scala 72:15:@53239.4]
  assign io_out_bits_wstrb_14 = io_in_bits_0_wstrb_14; // @[MuxN.scala 72:15:@53240.4]
  assign io_out_bits_wstrb_15 = io_in_bits_0_wstrb_15; // @[MuxN.scala 72:15:@53241.4]
  assign io_out_bits_wstrb_16 = io_in_bits_0_wstrb_16; // @[MuxN.scala 72:15:@53242.4]
  assign io_out_bits_wstrb_17 = io_in_bits_0_wstrb_17; // @[MuxN.scala 72:15:@53243.4]
  assign io_out_bits_wstrb_18 = io_in_bits_0_wstrb_18; // @[MuxN.scala 72:15:@53244.4]
  assign io_out_bits_wstrb_19 = io_in_bits_0_wstrb_19; // @[MuxN.scala 72:15:@53245.4]
  assign io_out_bits_wstrb_20 = io_in_bits_0_wstrb_20; // @[MuxN.scala 72:15:@53246.4]
  assign io_out_bits_wstrb_21 = io_in_bits_0_wstrb_21; // @[MuxN.scala 72:15:@53247.4]
  assign io_out_bits_wstrb_22 = io_in_bits_0_wstrb_22; // @[MuxN.scala 72:15:@53248.4]
  assign io_out_bits_wstrb_23 = io_in_bits_0_wstrb_23; // @[MuxN.scala 72:15:@53249.4]
  assign io_out_bits_wstrb_24 = io_in_bits_0_wstrb_24; // @[MuxN.scala 72:15:@53250.4]
  assign io_out_bits_wstrb_25 = io_in_bits_0_wstrb_25; // @[MuxN.scala 72:15:@53251.4]
  assign io_out_bits_wstrb_26 = io_in_bits_0_wstrb_26; // @[MuxN.scala 72:15:@53252.4]
  assign io_out_bits_wstrb_27 = io_in_bits_0_wstrb_27; // @[MuxN.scala 72:15:@53253.4]
  assign io_out_bits_wstrb_28 = io_in_bits_0_wstrb_28; // @[MuxN.scala 72:15:@53254.4]
  assign io_out_bits_wstrb_29 = io_in_bits_0_wstrb_29; // @[MuxN.scala 72:15:@53255.4]
  assign io_out_bits_wstrb_30 = io_in_bits_0_wstrb_30; // @[MuxN.scala 72:15:@53256.4]
  assign io_out_bits_wstrb_31 = io_in_bits_0_wstrb_31; // @[MuxN.scala 72:15:@53257.4]
  assign io_out_bits_wstrb_32 = io_in_bits_0_wstrb_32; // @[MuxN.scala 72:15:@53258.4]
  assign io_out_bits_wstrb_33 = io_in_bits_0_wstrb_33; // @[MuxN.scala 72:15:@53259.4]
  assign io_out_bits_wstrb_34 = io_in_bits_0_wstrb_34; // @[MuxN.scala 72:15:@53260.4]
  assign io_out_bits_wstrb_35 = io_in_bits_0_wstrb_35; // @[MuxN.scala 72:15:@53261.4]
  assign io_out_bits_wstrb_36 = io_in_bits_0_wstrb_36; // @[MuxN.scala 72:15:@53262.4]
  assign io_out_bits_wstrb_37 = io_in_bits_0_wstrb_37; // @[MuxN.scala 72:15:@53263.4]
  assign io_out_bits_wstrb_38 = io_in_bits_0_wstrb_38; // @[MuxN.scala 72:15:@53264.4]
  assign io_out_bits_wstrb_39 = io_in_bits_0_wstrb_39; // @[MuxN.scala 72:15:@53265.4]
  assign io_out_bits_wstrb_40 = io_in_bits_0_wstrb_40; // @[MuxN.scala 72:15:@53266.4]
  assign io_out_bits_wstrb_41 = io_in_bits_0_wstrb_41; // @[MuxN.scala 72:15:@53267.4]
  assign io_out_bits_wstrb_42 = io_in_bits_0_wstrb_42; // @[MuxN.scala 72:15:@53268.4]
  assign io_out_bits_wstrb_43 = io_in_bits_0_wstrb_43; // @[MuxN.scala 72:15:@53269.4]
  assign io_out_bits_wstrb_44 = io_in_bits_0_wstrb_44; // @[MuxN.scala 72:15:@53270.4]
  assign io_out_bits_wstrb_45 = io_in_bits_0_wstrb_45; // @[MuxN.scala 72:15:@53271.4]
  assign io_out_bits_wstrb_46 = io_in_bits_0_wstrb_46; // @[MuxN.scala 72:15:@53272.4]
  assign io_out_bits_wstrb_47 = io_in_bits_0_wstrb_47; // @[MuxN.scala 72:15:@53273.4]
  assign io_out_bits_wstrb_48 = io_in_bits_0_wstrb_48; // @[MuxN.scala 72:15:@53274.4]
  assign io_out_bits_wstrb_49 = io_in_bits_0_wstrb_49; // @[MuxN.scala 72:15:@53275.4]
  assign io_out_bits_wstrb_50 = io_in_bits_0_wstrb_50; // @[MuxN.scala 72:15:@53276.4]
  assign io_out_bits_wstrb_51 = io_in_bits_0_wstrb_51; // @[MuxN.scala 72:15:@53277.4]
  assign io_out_bits_wstrb_52 = io_in_bits_0_wstrb_52; // @[MuxN.scala 72:15:@53278.4]
  assign io_out_bits_wstrb_53 = io_in_bits_0_wstrb_53; // @[MuxN.scala 72:15:@53279.4]
  assign io_out_bits_wstrb_54 = io_in_bits_0_wstrb_54; // @[MuxN.scala 72:15:@53280.4]
  assign io_out_bits_wstrb_55 = io_in_bits_0_wstrb_55; // @[MuxN.scala 72:15:@53281.4]
  assign io_out_bits_wstrb_56 = io_in_bits_0_wstrb_56; // @[MuxN.scala 72:15:@53282.4]
  assign io_out_bits_wstrb_57 = io_in_bits_0_wstrb_57; // @[MuxN.scala 72:15:@53283.4]
  assign io_out_bits_wstrb_58 = io_in_bits_0_wstrb_58; // @[MuxN.scala 72:15:@53284.4]
  assign io_out_bits_wstrb_59 = io_in_bits_0_wstrb_59; // @[MuxN.scala 72:15:@53285.4]
  assign io_out_bits_wstrb_60 = io_in_bits_0_wstrb_60; // @[MuxN.scala 72:15:@53286.4]
  assign io_out_bits_wstrb_61 = io_in_bits_0_wstrb_61; // @[MuxN.scala 72:15:@53287.4]
  assign io_out_bits_wstrb_62 = io_in_bits_0_wstrb_62; // @[MuxN.scala 72:15:@53288.4]
  assign io_out_bits_wstrb_63 = io_in_bits_0_wstrb_63; // @[MuxN.scala 72:15:@53289.4]
endmodule
module ElementCounter( // @[:@53307.2]
  input         clock, // @[:@53308.4]
  input         reset, // @[:@53309.4]
  input         io_reset, // @[:@53310.4]
  input         io_enable, // @[:@53310.4]
  output [31:0] io_out // @[:@53310.4]
);
  reg [31:0] count; // @[Counter.scala 37:22:@53312.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_14; // @[Counter.scala 39:24:@53313.4]
  wire [31:0] newCount; // @[Counter.scala 39:24:@53314.4]
  wire [31:0] _GEN_0; // @[Counter.scala 43:26:@53319.6]
  wire [31:0] _GEN_1; // @[Counter.scala 41:18:@53315.4]
  assign _T_14 = count + 32'h1; // @[Counter.scala 39:24:@53313.4]
  assign newCount = count + 32'h1; // @[Counter.scala 39:24:@53314.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 43:26:@53319.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 41:18:@53315.4]
  assign io_out = count; // @[Counter.scala 47:10:@53322.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module StreamArbiter( // @[:@53324.2]
  input         clock, // @[:@53325.4]
  input         reset, // @[:@53326.4]
  output        io_app_0_cmd_ready, // @[:@53327.4]
  input         io_app_0_cmd_valid, // @[:@53327.4]
  input  [63:0] io_app_0_cmd_bits_addr, // @[:@53327.4]
  input  [31:0] io_app_0_cmd_bits_size, // @[:@53327.4]
  input         io_app_0_cmd_bits_isWr, // @[:@53327.4]
  input  [31:0] io_app_0_cmd_bits_tag, // @[:@53327.4]
  output        io_app_0_wdata_ready, // @[:@53327.4]
  input         io_app_0_wdata_valid, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_0, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_1, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_2, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_3, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_4, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_5, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_6, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_7, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_8, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_9, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_10, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_11, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_12, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_13, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_14, // @[:@53327.4]
  input  [31:0] io_app_0_wdata_bits_wdata_15, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_0, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_1, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_2, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_3, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_4, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_5, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_6, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_7, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_8, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_9, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_10, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_11, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_12, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_13, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_14, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_15, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_16, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_17, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_18, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_19, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_20, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_21, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_22, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_23, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_24, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_25, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_26, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_27, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_28, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_29, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_30, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_31, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_32, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_33, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_34, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_35, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_36, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_37, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_38, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_39, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_40, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_41, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_42, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_43, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_44, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_45, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_46, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_47, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_48, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_49, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_50, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_51, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_52, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_53, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_54, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_55, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_56, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_57, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_58, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_59, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_60, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_61, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_62, // @[:@53327.4]
  input         io_app_0_wdata_bits_wstrb_63, // @[:@53327.4]
  input         io_app_0_rresp_ready, // @[:@53327.4]
  input         io_app_0_wresp_ready, // @[:@53327.4]
  output        io_app_0_wresp_valid, // @[:@53327.4]
  input         io_dram_cmd_ready, // @[:@53327.4]
  output        io_dram_cmd_valid, // @[:@53327.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@53327.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@53327.4]
  output        io_dram_cmd_bits_isWr, // @[:@53327.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@53327.4]
  input         io_dram_wdata_ready, // @[:@53327.4]
  output        io_dram_wdata_valid, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@53327.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@53327.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@53327.4]
  output        io_dram_rresp_ready, // @[:@53327.4]
  output        io_dram_wresp_ready, // @[:@53327.4]
  input         io_dram_wresp_valid, // @[:@53327.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@53327.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@53556.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@53556.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@53556.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@53556.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@53556.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@53563.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@53563.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@53563.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@53563.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@53563.4]
  wire  cmdMux_io_in_ready; // @[StreamArbiter.scala 25:22:@53573.4]
  wire  cmdMux_io_in_valid; // @[StreamArbiter.scala 25:22:@53573.4]
  wire [63:0] cmdMux_io_in_bits_0_addr; // @[StreamArbiter.scala 25:22:@53573.4]
  wire [31:0] cmdMux_io_in_bits_0_size; // @[StreamArbiter.scala 25:22:@53573.4]
  wire  cmdMux_io_in_bits_0_isWr; // @[StreamArbiter.scala 25:22:@53573.4]
  wire [31:0] cmdMux_io_in_bits_0_tag; // @[StreamArbiter.scala 25:22:@53573.4]
  wire  cmdMux_io_out_ready; // @[StreamArbiter.scala 25:22:@53573.4]
  wire  cmdMux_io_out_valid; // @[StreamArbiter.scala 25:22:@53573.4]
  wire [63:0] cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 25:22:@53573.4]
  wire [31:0] cmdMux_io_out_bits_size; // @[StreamArbiter.scala 25:22:@53573.4]
  wire  cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 25:22:@53573.4]
  wire [31:0] cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 25:22:@53573.4]
  wire  wdataMux_io_in_ready; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_valid; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_0; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_1; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_2; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_3; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_4; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_5; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_6; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_7; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_8; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_9; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_10; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_11; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_12; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_13; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_14; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_15; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_0; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_1; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_2; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_3; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_4; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_5; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_6; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_7; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_8; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_9; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_10; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_11; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_12; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_13; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_14; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_15; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_16; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_17; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_18; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_19; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_20; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_21; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_22; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_23; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_24; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_25; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_26; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_27; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_28; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_29; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_30; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_31; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_32; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_33; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_34; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_35; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_36; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_37; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_38; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_39; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_40; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_41; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_42; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_43; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_44; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_45; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_46; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_47; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_48; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_49; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_50; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_51; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_52; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_53; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_54; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_55; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_56; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_57; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_58; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_59; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_60; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_61; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_62; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_in_bits_0_wstrb_63; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_ready; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_valid; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 35:24:@53596.4]
  wire [31:0] wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 35:24:@53596.4]
  wire  elementCtr_clock; // @[StreamArbiter.scala 36:26:@53599.4]
  wire  elementCtr_reset; // @[StreamArbiter.scala 36:26:@53599.4]
  wire  elementCtr_io_reset; // @[StreamArbiter.scala 36:26:@53599.4]
  wire  elementCtr_io_enable; // @[StreamArbiter.scala 36:26:@53599.4]
  wire [31:0] elementCtr_io_out; // @[StreamArbiter.scala 36:26:@53599.4]
  wire  _T_346; // @[package.scala 96:25:@53568.4 package.scala 96:25:@53569.4]
  wire  cmdIdx; // @[StreamArbiter.scala 21:16:@53570.4]
  wire [1:0] cmdInDecoder; // @[OneHot.scala 45:35:@53572.4]
  wire  _T_355; // @[FringeBundles.scala 114:28:@53588.4]
  wire [22:0] _T_356; // @[FringeBundles.scala 114:28:@53590.4]
  wire [23:0] _T_358; // @[FringeBundles.scala 115:37:@53593.4]
  wire  _T_360; // @[StreamArbiter.scala 37:49:@53602.4]
  wire [31:0] _T_365; // @[:@53606.4 :@53607.4]
  wire [7:0] _T_366; // @[FringeBundles.scala 114:28:@53608.4]
  wire [255:0] cmdOutDecoder; // @[OneHot.scala 45:35:@53614.4]
  wire  _T_379; // @[StreamArbiter.scala 42:78:@53617.4]
  wire  _T_380; // @[StreamArbiter.scala 42:121:@53618.4]
  wire [7:0] _T_395; // @[FringeBundles.scala 140:28:@53805.4]
  wire [255:0] wrespDecoder; // @[OneHot.scala 45:35:@53812.4]
  wire  _T_400; // @[StreamArbiter.scala 61:55:@53817.4]
  wire  _T_403; // @[StreamArbiter.scala 62:85:@53821.4]
  wire  _T_404; // @[StreamArbiter.scala 62:70:@53822.4]
  wire  _T_409; // @[StreamArbiter.scala 67:58:@53846.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@53556.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@53563.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  MuxPipe cmdMux ( // @[StreamArbiter.scala 25:22:@53573.4]
    .io_in_ready(cmdMux_io_in_ready),
    .io_in_valid(cmdMux_io_in_valid),
    .io_in_bits_0_addr(cmdMux_io_in_bits_0_addr),
    .io_in_bits_0_size(cmdMux_io_in_bits_0_size),
    .io_in_bits_0_isWr(cmdMux_io_in_bits_0_isWr),
    .io_in_bits_0_tag(cmdMux_io_in_bits_0_tag),
    .io_out_ready(cmdMux_io_out_ready),
    .io_out_valid(cmdMux_io_out_valid),
    .io_out_bits_addr(cmdMux_io_out_bits_addr),
    .io_out_bits_size(cmdMux_io_out_bits_size),
    .io_out_bits_isWr(cmdMux_io_out_bits_isWr),
    .io_out_bits_tag(cmdMux_io_out_bits_tag)
  );
  MuxPipe_1 wdataMux ( // @[StreamArbiter.scala 35:24:@53596.4]
    .io_in_ready(wdataMux_io_in_ready),
    .io_in_valid(wdataMux_io_in_valid),
    .io_in_bits_0_wdata_0(wdataMux_io_in_bits_0_wdata_0),
    .io_in_bits_0_wdata_1(wdataMux_io_in_bits_0_wdata_1),
    .io_in_bits_0_wdata_2(wdataMux_io_in_bits_0_wdata_2),
    .io_in_bits_0_wdata_3(wdataMux_io_in_bits_0_wdata_3),
    .io_in_bits_0_wdata_4(wdataMux_io_in_bits_0_wdata_4),
    .io_in_bits_0_wdata_5(wdataMux_io_in_bits_0_wdata_5),
    .io_in_bits_0_wdata_6(wdataMux_io_in_bits_0_wdata_6),
    .io_in_bits_0_wdata_7(wdataMux_io_in_bits_0_wdata_7),
    .io_in_bits_0_wdata_8(wdataMux_io_in_bits_0_wdata_8),
    .io_in_bits_0_wdata_9(wdataMux_io_in_bits_0_wdata_9),
    .io_in_bits_0_wdata_10(wdataMux_io_in_bits_0_wdata_10),
    .io_in_bits_0_wdata_11(wdataMux_io_in_bits_0_wdata_11),
    .io_in_bits_0_wdata_12(wdataMux_io_in_bits_0_wdata_12),
    .io_in_bits_0_wdata_13(wdataMux_io_in_bits_0_wdata_13),
    .io_in_bits_0_wdata_14(wdataMux_io_in_bits_0_wdata_14),
    .io_in_bits_0_wdata_15(wdataMux_io_in_bits_0_wdata_15),
    .io_in_bits_0_wstrb_0(wdataMux_io_in_bits_0_wstrb_0),
    .io_in_bits_0_wstrb_1(wdataMux_io_in_bits_0_wstrb_1),
    .io_in_bits_0_wstrb_2(wdataMux_io_in_bits_0_wstrb_2),
    .io_in_bits_0_wstrb_3(wdataMux_io_in_bits_0_wstrb_3),
    .io_in_bits_0_wstrb_4(wdataMux_io_in_bits_0_wstrb_4),
    .io_in_bits_0_wstrb_5(wdataMux_io_in_bits_0_wstrb_5),
    .io_in_bits_0_wstrb_6(wdataMux_io_in_bits_0_wstrb_6),
    .io_in_bits_0_wstrb_7(wdataMux_io_in_bits_0_wstrb_7),
    .io_in_bits_0_wstrb_8(wdataMux_io_in_bits_0_wstrb_8),
    .io_in_bits_0_wstrb_9(wdataMux_io_in_bits_0_wstrb_9),
    .io_in_bits_0_wstrb_10(wdataMux_io_in_bits_0_wstrb_10),
    .io_in_bits_0_wstrb_11(wdataMux_io_in_bits_0_wstrb_11),
    .io_in_bits_0_wstrb_12(wdataMux_io_in_bits_0_wstrb_12),
    .io_in_bits_0_wstrb_13(wdataMux_io_in_bits_0_wstrb_13),
    .io_in_bits_0_wstrb_14(wdataMux_io_in_bits_0_wstrb_14),
    .io_in_bits_0_wstrb_15(wdataMux_io_in_bits_0_wstrb_15),
    .io_in_bits_0_wstrb_16(wdataMux_io_in_bits_0_wstrb_16),
    .io_in_bits_0_wstrb_17(wdataMux_io_in_bits_0_wstrb_17),
    .io_in_bits_0_wstrb_18(wdataMux_io_in_bits_0_wstrb_18),
    .io_in_bits_0_wstrb_19(wdataMux_io_in_bits_0_wstrb_19),
    .io_in_bits_0_wstrb_20(wdataMux_io_in_bits_0_wstrb_20),
    .io_in_bits_0_wstrb_21(wdataMux_io_in_bits_0_wstrb_21),
    .io_in_bits_0_wstrb_22(wdataMux_io_in_bits_0_wstrb_22),
    .io_in_bits_0_wstrb_23(wdataMux_io_in_bits_0_wstrb_23),
    .io_in_bits_0_wstrb_24(wdataMux_io_in_bits_0_wstrb_24),
    .io_in_bits_0_wstrb_25(wdataMux_io_in_bits_0_wstrb_25),
    .io_in_bits_0_wstrb_26(wdataMux_io_in_bits_0_wstrb_26),
    .io_in_bits_0_wstrb_27(wdataMux_io_in_bits_0_wstrb_27),
    .io_in_bits_0_wstrb_28(wdataMux_io_in_bits_0_wstrb_28),
    .io_in_bits_0_wstrb_29(wdataMux_io_in_bits_0_wstrb_29),
    .io_in_bits_0_wstrb_30(wdataMux_io_in_bits_0_wstrb_30),
    .io_in_bits_0_wstrb_31(wdataMux_io_in_bits_0_wstrb_31),
    .io_in_bits_0_wstrb_32(wdataMux_io_in_bits_0_wstrb_32),
    .io_in_bits_0_wstrb_33(wdataMux_io_in_bits_0_wstrb_33),
    .io_in_bits_0_wstrb_34(wdataMux_io_in_bits_0_wstrb_34),
    .io_in_bits_0_wstrb_35(wdataMux_io_in_bits_0_wstrb_35),
    .io_in_bits_0_wstrb_36(wdataMux_io_in_bits_0_wstrb_36),
    .io_in_bits_0_wstrb_37(wdataMux_io_in_bits_0_wstrb_37),
    .io_in_bits_0_wstrb_38(wdataMux_io_in_bits_0_wstrb_38),
    .io_in_bits_0_wstrb_39(wdataMux_io_in_bits_0_wstrb_39),
    .io_in_bits_0_wstrb_40(wdataMux_io_in_bits_0_wstrb_40),
    .io_in_bits_0_wstrb_41(wdataMux_io_in_bits_0_wstrb_41),
    .io_in_bits_0_wstrb_42(wdataMux_io_in_bits_0_wstrb_42),
    .io_in_bits_0_wstrb_43(wdataMux_io_in_bits_0_wstrb_43),
    .io_in_bits_0_wstrb_44(wdataMux_io_in_bits_0_wstrb_44),
    .io_in_bits_0_wstrb_45(wdataMux_io_in_bits_0_wstrb_45),
    .io_in_bits_0_wstrb_46(wdataMux_io_in_bits_0_wstrb_46),
    .io_in_bits_0_wstrb_47(wdataMux_io_in_bits_0_wstrb_47),
    .io_in_bits_0_wstrb_48(wdataMux_io_in_bits_0_wstrb_48),
    .io_in_bits_0_wstrb_49(wdataMux_io_in_bits_0_wstrb_49),
    .io_in_bits_0_wstrb_50(wdataMux_io_in_bits_0_wstrb_50),
    .io_in_bits_0_wstrb_51(wdataMux_io_in_bits_0_wstrb_51),
    .io_in_bits_0_wstrb_52(wdataMux_io_in_bits_0_wstrb_52),
    .io_in_bits_0_wstrb_53(wdataMux_io_in_bits_0_wstrb_53),
    .io_in_bits_0_wstrb_54(wdataMux_io_in_bits_0_wstrb_54),
    .io_in_bits_0_wstrb_55(wdataMux_io_in_bits_0_wstrb_55),
    .io_in_bits_0_wstrb_56(wdataMux_io_in_bits_0_wstrb_56),
    .io_in_bits_0_wstrb_57(wdataMux_io_in_bits_0_wstrb_57),
    .io_in_bits_0_wstrb_58(wdataMux_io_in_bits_0_wstrb_58),
    .io_in_bits_0_wstrb_59(wdataMux_io_in_bits_0_wstrb_59),
    .io_in_bits_0_wstrb_60(wdataMux_io_in_bits_0_wstrb_60),
    .io_in_bits_0_wstrb_61(wdataMux_io_in_bits_0_wstrb_61),
    .io_in_bits_0_wstrb_62(wdataMux_io_in_bits_0_wstrb_62),
    .io_in_bits_0_wstrb_63(wdataMux_io_in_bits_0_wstrb_63),
    .io_out_ready(wdataMux_io_out_ready),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  ElementCounter elementCtr ( // @[StreamArbiter.scala 36:26:@53599.4]
    .clock(elementCtr_clock),
    .reset(elementCtr_reset),
    .io_reset(elementCtr_io_reset),
    .io_enable(elementCtr_io_enable),
    .io_out(elementCtr_io_out)
  );
  assign _T_346 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@53568.4 package.scala 96:25:@53569.4]
  assign cmdIdx = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[StreamArbiter.scala 21:16:@53570.4]
  assign cmdInDecoder = 2'h1 << cmdIdx; // @[OneHot.scala 45:35:@53572.4]
  assign _T_355 = io_app_0_cmd_bits_tag[8]; // @[FringeBundles.scala 114:28:@53588.4]
  assign _T_356 = io_app_0_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@53590.4]
  assign _T_358 = {_T_356,_T_355}; // @[FringeBundles.scala 115:37:@53593.4]
  assign _T_360 = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:49:@53602.4]
  assign _T_365 = cmdMux_io_out_bits_tag; // @[:@53606.4 :@53607.4]
  assign _T_366 = _T_365[7:0]; // @[FringeBundles.scala 114:28:@53608.4]
  assign cmdOutDecoder = 256'h1 << _T_366; // @[OneHot.scala 45:35:@53614.4]
  assign _T_379 = io_app_0_wdata_valid & cmdMux_io_out_valid; // @[StreamArbiter.scala 42:78:@53617.4]
  assign _T_380 = elementCtr_io_out < cmdMux_io_out_bits_size; // @[StreamArbiter.scala 42:121:@53618.4]
  assign _T_395 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@53805.4]
  assign wrespDecoder = 256'h1 << _T_395; // @[OneHot.scala 45:35:@53812.4]
  assign _T_400 = cmdInDecoder[0]; // @[StreamArbiter.scala 61:55:@53817.4]
  assign _T_403 = cmdOutDecoder[0]; // @[StreamArbiter.scala 62:85:@53821.4]
  assign _T_404 = _T_360 & _T_403; // @[StreamArbiter.scala 62:70:@53822.4]
  assign _T_409 = wrespDecoder[0]; // @[StreamArbiter.scala 67:58:@53846.4]
  assign io_app_0_cmd_ready = cmdMux_io_in_ready & _T_400; // @[StreamArbiter.scala 61:19:@53819.4]
  assign io_app_0_wdata_ready = _T_404 & _T_380; // @[StreamArbiter.scala 62:21:@53825.4]
  assign io_app_0_wresp_valid = io_dram_wresp_valid & _T_409; // @[StreamArbiter.scala 67:21:@53848.4]
  assign io_dram_cmd_valid = cmdMux_io_out_valid; // @[StreamArbiter.scala 46:15:@53708.4]
  assign io_dram_cmd_bits_addr = cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 46:15:@53707.4]
  assign io_dram_cmd_bits_size = cmdMux_io_out_bits_size; // @[StreamArbiter.scala 46:15:@53706.4]
  assign io_dram_cmd_bits_isWr = cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 46:15:@53704.4]
  assign io_dram_cmd_bits_tag = cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 46:15:@53703.4]
  assign io_dram_wdata_valid = wdataMux_io_out_valid; // @[StreamArbiter.scala 47:17:@53791.4]
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 47:17:@53775.4]
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 47:17:@53776.4]
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 47:17:@53777.4]
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 47:17:@53778.4]
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 47:17:@53779.4]
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 47:17:@53780.4]
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 47:17:@53781.4]
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 47:17:@53782.4]
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 47:17:@53783.4]
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 47:17:@53784.4]
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 47:17:@53785.4]
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 47:17:@53786.4]
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 47:17:@53787.4]
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 47:17:@53788.4]
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 47:17:@53789.4]
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 47:17:@53790.4]
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 47:17:@53711.4]
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 47:17:@53712.4]
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 47:17:@53713.4]
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 47:17:@53714.4]
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 47:17:@53715.4]
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 47:17:@53716.4]
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 47:17:@53717.4]
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 47:17:@53718.4]
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 47:17:@53719.4]
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 47:17:@53720.4]
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 47:17:@53721.4]
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 47:17:@53722.4]
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 47:17:@53723.4]
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 47:17:@53724.4]
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 47:17:@53725.4]
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 47:17:@53726.4]
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 47:17:@53727.4]
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 47:17:@53728.4]
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 47:17:@53729.4]
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 47:17:@53730.4]
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 47:17:@53731.4]
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 47:17:@53732.4]
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 47:17:@53733.4]
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 47:17:@53734.4]
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 47:17:@53735.4]
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 47:17:@53736.4]
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 47:17:@53737.4]
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 47:17:@53738.4]
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 47:17:@53739.4]
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 47:17:@53740.4]
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 47:17:@53741.4]
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 47:17:@53742.4]
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 47:17:@53743.4]
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 47:17:@53744.4]
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 47:17:@53745.4]
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 47:17:@53746.4]
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 47:17:@53747.4]
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 47:17:@53748.4]
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 47:17:@53749.4]
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 47:17:@53750.4]
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 47:17:@53751.4]
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 47:17:@53752.4]
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 47:17:@53753.4]
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 47:17:@53754.4]
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 47:17:@53755.4]
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 47:17:@53756.4]
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 47:17:@53757.4]
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 47:17:@53758.4]
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 47:17:@53759.4]
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 47:17:@53760.4]
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 47:17:@53761.4]
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 47:17:@53762.4]
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 47:17:@53763.4]
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 47:17:@53764.4]
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 47:17:@53765.4]
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 47:17:@53766.4]
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 47:17:@53767.4]
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 47:17:@53768.4]
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 47:17:@53769.4]
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 47:17:@53770.4]
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 47:17:@53771.4]
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 47:17:@53772.4]
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 47:17:@53773.4]
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 47:17:@53774.4]
  assign io_dram_rresp_ready = io_app_0_rresp_ready; // @[StreamArbiter.scala 72:23:@53852.4]
  assign io_dram_wresp_ready = io_app_0_wresp_ready; // @[StreamArbiter.scala 73:23:@53855.4]
  assign RetimeWrapper_clock = clock; // @[:@53557.4]
  assign RetimeWrapper_reset = reset; // @[:@53558.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@53560.4]
  assign RetimeWrapper_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@53559.4]
  assign RetimeWrapper_1_clock = clock; // @[:@53564.4]
  assign RetimeWrapper_1_reset = reset; // @[:@53565.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@53567.4]
  assign RetimeWrapper_1_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@53566.4]
  assign cmdMux_io_in_valid = io_app_0_cmd_valid; // @[StreamArbiter.scala 26:22:@53576.4]
  assign cmdMux_io_in_bits_0_addr = io_app_0_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@53582.4]
  assign cmdMux_io_in_bits_0_size = io_app_0_cmd_bits_size; // @[StreamArbiter.scala 29:9:@53581.4]
  assign cmdMux_io_in_bits_0_isWr = io_app_0_cmd_bits_isWr; // @[StreamArbiter.scala 29:9:@53579.4]
  assign cmdMux_io_in_bits_0_tag = {_T_358,8'h0}; // @[StreamArbiter.scala 29:9:@53578.4 FringeBundles.scala 115:32:@53595.4]
  assign cmdMux_io_out_ready = io_dram_cmd_valid & io_dram_cmd_ready; // @[StreamArbiter.scala 46:15:@53709.4 StreamArbiter.scala 57:23:@53815.4]
  assign wdataMux_io_in_valid = _T_379 & _T_380; // @[StreamArbiter.scala 42:24:@53620.4]
  assign wdataMux_io_in_bits_0_wdata_0 = io_app_0_wdata_bits_wdata_0; // @[StreamArbiter.scala 44:23:@53687.4]
  assign wdataMux_io_in_bits_0_wdata_1 = io_app_0_wdata_bits_wdata_1; // @[StreamArbiter.scala 44:23:@53688.4]
  assign wdataMux_io_in_bits_0_wdata_2 = io_app_0_wdata_bits_wdata_2; // @[StreamArbiter.scala 44:23:@53689.4]
  assign wdataMux_io_in_bits_0_wdata_3 = io_app_0_wdata_bits_wdata_3; // @[StreamArbiter.scala 44:23:@53690.4]
  assign wdataMux_io_in_bits_0_wdata_4 = io_app_0_wdata_bits_wdata_4; // @[StreamArbiter.scala 44:23:@53691.4]
  assign wdataMux_io_in_bits_0_wdata_5 = io_app_0_wdata_bits_wdata_5; // @[StreamArbiter.scala 44:23:@53692.4]
  assign wdataMux_io_in_bits_0_wdata_6 = io_app_0_wdata_bits_wdata_6; // @[StreamArbiter.scala 44:23:@53693.4]
  assign wdataMux_io_in_bits_0_wdata_7 = io_app_0_wdata_bits_wdata_7; // @[StreamArbiter.scala 44:23:@53694.4]
  assign wdataMux_io_in_bits_0_wdata_8 = io_app_0_wdata_bits_wdata_8; // @[StreamArbiter.scala 44:23:@53695.4]
  assign wdataMux_io_in_bits_0_wdata_9 = io_app_0_wdata_bits_wdata_9; // @[StreamArbiter.scala 44:23:@53696.4]
  assign wdataMux_io_in_bits_0_wdata_10 = io_app_0_wdata_bits_wdata_10; // @[StreamArbiter.scala 44:23:@53697.4]
  assign wdataMux_io_in_bits_0_wdata_11 = io_app_0_wdata_bits_wdata_11; // @[StreamArbiter.scala 44:23:@53698.4]
  assign wdataMux_io_in_bits_0_wdata_12 = io_app_0_wdata_bits_wdata_12; // @[StreamArbiter.scala 44:23:@53699.4]
  assign wdataMux_io_in_bits_0_wdata_13 = io_app_0_wdata_bits_wdata_13; // @[StreamArbiter.scala 44:23:@53700.4]
  assign wdataMux_io_in_bits_0_wdata_14 = io_app_0_wdata_bits_wdata_14; // @[StreamArbiter.scala 44:23:@53701.4]
  assign wdataMux_io_in_bits_0_wdata_15 = io_app_0_wdata_bits_wdata_15; // @[StreamArbiter.scala 44:23:@53702.4]
  assign wdataMux_io_in_bits_0_wstrb_0 = io_app_0_wdata_bits_wstrb_0; // @[StreamArbiter.scala 44:23:@53623.4]
  assign wdataMux_io_in_bits_0_wstrb_1 = io_app_0_wdata_bits_wstrb_1; // @[StreamArbiter.scala 44:23:@53624.4]
  assign wdataMux_io_in_bits_0_wstrb_2 = io_app_0_wdata_bits_wstrb_2; // @[StreamArbiter.scala 44:23:@53625.4]
  assign wdataMux_io_in_bits_0_wstrb_3 = io_app_0_wdata_bits_wstrb_3; // @[StreamArbiter.scala 44:23:@53626.4]
  assign wdataMux_io_in_bits_0_wstrb_4 = io_app_0_wdata_bits_wstrb_4; // @[StreamArbiter.scala 44:23:@53627.4]
  assign wdataMux_io_in_bits_0_wstrb_5 = io_app_0_wdata_bits_wstrb_5; // @[StreamArbiter.scala 44:23:@53628.4]
  assign wdataMux_io_in_bits_0_wstrb_6 = io_app_0_wdata_bits_wstrb_6; // @[StreamArbiter.scala 44:23:@53629.4]
  assign wdataMux_io_in_bits_0_wstrb_7 = io_app_0_wdata_bits_wstrb_7; // @[StreamArbiter.scala 44:23:@53630.4]
  assign wdataMux_io_in_bits_0_wstrb_8 = io_app_0_wdata_bits_wstrb_8; // @[StreamArbiter.scala 44:23:@53631.4]
  assign wdataMux_io_in_bits_0_wstrb_9 = io_app_0_wdata_bits_wstrb_9; // @[StreamArbiter.scala 44:23:@53632.4]
  assign wdataMux_io_in_bits_0_wstrb_10 = io_app_0_wdata_bits_wstrb_10; // @[StreamArbiter.scala 44:23:@53633.4]
  assign wdataMux_io_in_bits_0_wstrb_11 = io_app_0_wdata_bits_wstrb_11; // @[StreamArbiter.scala 44:23:@53634.4]
  assign wdataMux_io_in_bits_0_wstrb_12 = io_app_0_wdata_bits_wstrb_12; // @[StreamArbiter.scala 44:23:@53635.4]
  assign wdataMux_io_in_bits_0_wstrb_13 = io_app_0_wdata_bits_wstrb_13; // @[StreamArbiter.scala 44:23:@53636.4]
  assign wdataMux_io_in_bits_0_wstrb_14 = io_app_0_wdata_bits_wstrb_14; // @[StreamArbiter.scala 44:23:@53637.4]
  assign wdataMux_io_in_bits_0_wstrb_15 = io_app_0_wdata_bits_wstrb_15; // @[StreamArbiter.scala 44:23:@53638.4]
  assign wdataMux_io_in_bits_0_wstrb_16 = io_app_0_wdata_bits_wstrb_16; // @[StreamArbiter.scala 44:23:@53639.4]
  assign wdataMux_io_in_bits_0_wstrb_17 = io_app_0_wdata_bits_wstrb_17; // @[StreamArbiter.scala 44:23:@53640.4]
  assign wdataMux_io_in_bits_0_wstrb_18 = io_app_0_wdata_bits_wstrb_18; // @[StreamArbiter.scala 44:23:@53641.4]
  assign wdataMux_io_in_bits_0_wstrb_19 = io_app_0_wdata_bits_wstrb_19; // @[StreamArbiter.scala 44:23:@53642.4]
  assign wdataMux_io_in_bits_0_wstrb_20 = io_app_0_wdata_bits_wstrb_20; // @[StreamArbiter.scala 44:23:@53643.4]
  assign wdataMux_io_in_bits_0_wstrb_21 = io_app_0_wdata_bits_wstrb_21; // @[StreamArbiter.scala 44:23:@53644.4]
  assign wdataMux_io_in_bits_0_wstrb_22 = io_app_0_wdata_bits_wstrb_22; // @[StreamArbiter.scala 44:23:@53645.4]
  assign wdataMux_io_in_bits_0_wstrb_23 = io_app_0_wdata_bits_wstrb_23; // @[StreamArbiter.scala 44:23:@53646.4]
  assign wdataMux_io_in_bits_0_wstrb_24 = io_app_0_wdata_bits_wstrb_24; // @[StreamArbiter.scala 44:23:@53647.4]
  assign wdataMux_io_in_bits_0_wstrb_25 = io_app_0_wdata_bits_wstrb_25; // @[StreamArbiter.scala 44:23:@53648.4]
  assign wdataMux_io_in_bits_0_wstrb_26 = io_app_0_wdata_bits_wstrb_26; // @[StreamArbiter.scala 44:23:@53649.4]
  assign wdataMux_io_in_bits_0_wstrb_27 = io_app_0_wdata_bits_wstrb_27; // @[StreamArbiter.scala 44:23:@53650.4]
  assign wdataMux_io_in_bits_0_wstrb_28 = io_app_0_wdata_bits_wstrb_28; // @[StreamArbiter.scala 44:23:@53651.4]
  assign wdataMux_io_in_bits_0_wstrb_29 = io_app_0_wdata_bits_wstrb_29; // @[StreamArbiter.scala 44:23:@53652.4]
  assign wdataMux_io_in_bits_0_wstrb_30 = io_app_0_wdata_bits_wstrb_30; // @[StreamArbiter.scala 44:23:@53653.4]
  assign wdataMux_io_in_bits_0_wstrb_31 = io_app_0_wdata_bits_wstrb_31; // @[StreamArbiter.scala 44:23:@53654.4]
  assign wdataMux_io_in_bits_0_wstrb_32 = io_app_0_wdata_bits_wstrb_32; // @[StreamArbiter.scala 44:23:@53655.4]
  assign wdataMux_io_in_bits_0_wstrb_33 = io_app_0_wdata_bits_wstrb_33; // @[StreamArbiter.scala 44:23:@53656.4]
  assign wdataMux_io_in_bits_0_wstrb_34 = io_app_0_wdata_bits_wstrb_34; // @[StreamArbiter.scala 44:23:@53657.4]
  assign wdataMux_io_in_bits_0_wstrb_35 = io_app_0_wdata_bits_wstrb_35; // @[StreamArbiter.scala 44:23:@53658.4]
  assign wdataMux_io_in_bits_0_wstrb_36 = io_app_0_wdata_bits_wstrb_36; // @[StreamArbiter.scala 44:23:@53659.4]
  assign wdataMux_io_in_bits_0_wstrb_37 = io_app_0_wdata_bits_wstrb_37; // @[StreamArbiter.scala 44:23:@53660.4]
  assign wdataMux_io_in_bits_0_wstrb_38 = io_app_0_wdata_bits_wstrb_38; // @[StreamArbiter.scala 44:23:@53661.4]
  assign wdataMux_io_in_bits_0_wstrb_39 = io_app_0_wdata_bits_wstrb_39; // @[StreamArbiter.scala 44:23:@53662.4]
  assign wdataMux_io_in_bits_0_wstrb_40 = io_app_0_wdata_bits_wstrb_40; // @[StreamArbiter.scala 44:23:@53663.4]
  assign wdataMux_io_in_bits_0_wstrb_41 = io_app_0_wdata_bits_wstrb_41; // @[StreamArbiter.scala 44:23:@53664.4]
  assign wdataMux_io_in_bits_0_wstrb_42 = io_app_0_wdata_bits_wstrb_42; // @[StreamArbiter.scala 44:23:@53665.4]
  assign wdataMux_io_in_bits_0_wstrb_43 = io_app_0_wdata_bits_wstrb_43; // @[StreamArbiter.scala 44:23:@53666.4]
  assign wdataMux_io_in_bits_0_wstrb_44 = io_app_0_wdata_bits_wstrb_44; // @[StreamArbiter.scala 44:23:@53667.4]
  assign wdataMux_io_in_bits_0_wstrb_45 = io_app_0_wdata_bits_wstrb_45; // @[StreamArbiter.scala 44:23:@53668.4]
  assign wdataMux_io_in_bits_0_wstrb_46 = io_app_0_wdata_bits_wstrb_46; // @[StreamArbiter.scala 44:23:@53669.4]
  assign wdataMux_io_in_bits_0_wstrb_47 = io_app_0_wdata_bits_wstrb_47; // @[StreamArbiter.scala 44:23:@53670.4]
  assign wdataMux_io_in_bits_0_wstrb_48 = io_app_0_wdata_bits_wstrb_48; // @[StreamArbiter.scala 44:23:@53671.4]
  assign wdataMux_io_in_bits_0_wstrb_49 = io_app_0_wdata_bits_wstrb_49; // @[StreamArbiter.scala 44:23:@53672.4]
  assign wdataMux_io_in_bits_0_wstrb_50 = io_app_0_wdata_bits_wstrb_50; // @[StreamArbiter.scala 44:23:@53673.4]
  assign wdataMux_io_in_bits_0_wstrb_51 = io_app_0_wdata_bits_wstrb_51; // @[StreamArbiter.scala 44:23:@53674.4]
  assign wdataMux_io_in_bits_0_wstrb_52 = io_app_0_wdata_bits_wstrb_52; // @[StreamArbiter.scala 44:23:@53675.4]
  assign wdataMux_io_in_bits_0_wstrb_53 = io_app_0_wdata_bits_wstrb_53; // @[StreamArbiter.scala 44:23:@53676.4]
  assign wdataMux_io_in_bits_0_wstrb_54 = io_app_0_wdata_bits_wstrb_54; // @[StreamArbiter.scala 44:23:@53677.4]
  assign wdataMux_io_in_bits_0_wstrb_55 = io_app_0_wdata_bits_wstrb_55; // @[StreamArbiter.scala 44:23:@53678.4]
  assign wdataMux_io_in_bits_0_wstrb_56 = io_app_0_wdata_bits_wstrb_56; // @[StreamArbiter.scala 44:23:@53679.4]
  assign wdataMux_io_in_bits_0_wstrb_57 = io_app_0_wdata_bits_wstrb_57; // @[StreamArbiter.scala 44:23:@53680.4]
  assign wdataMux_io_in_bits_0_wstrb_58 = io_app_0_wdata_bits_wstrb_58; // @[StreamArbiter.scala 44:23:@53681.4]
  assign wdataMux_io_in_bits_0_wstrb_59 = io_app_0_wdata_bits_wstrb_59; // @[StreamArbiter.scala 44:23:@53682.4]
  assign wdataMux_io_in_bits_0_wstrb_60 = io_app_0_wdata_bits_wstrb_60; // @[StreamArbiter.scala 44:23:@53683.4]
  assign wdataMux_io_in_bits_0_wstrb_61 = io_app_0_wdata_bits_wstrb_61; // @[StreamArbiter.scala 44:23:@53684.4]
  assign wdataMux_io_in_bits_0_wstrb_62 = io_app_0_wdata_bits_wstrb_62; // @[StreamArbiter.scala 44:23:@53685.4]
  assign wdataMux_io_in_bits_0_wstrb_63 = io_app_0_wdata_bits_wstrb_63; // @[StreamArbiter.scala 44:23:@53686.4]
  assign wdataMux_io_out_ready = io_dram_wdata_valid & io_dram_wdata_ready; // @[StreamArbiter.scala 47:17:@53792.4 StreamArbiter.scala 58:25:@53816.4]
  assign elementCtr_clock = clock; // @[:@53600.4]
  assign elementCtr_reset = reset; // @[:@53601.4]
  assign elementCtr_io_reset = cmdMux_io_out_ready; // @[StreamArbiter.scala 38:23:@53604.4]
  assign elementCtr_io_enable = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:24:@53603.4]
endmodule
module Counter_72( // @[:@53857.2]
  input         clock, // @[:@53858.4]
  input         reset, // @[:@53859.4]
  input         io_reset, // @[:@53860.4]
  input         io_enable, // @[:@53860.4]
  input  [31:0] io_stride, // @[:@53860.4]
  output [31:0] io_out, // @[:@53860.4]
  output [31:0] io_next // @[:@53860.4]
);
  reg [31:0] count; // @[Counter.scala 15:22:@53862.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_17; // @[Counter.scala 17:24:@53863.4]
  wire [31:0] newCount; // @[Counter.scala 17:24:@53864.4]
  wire [31:0] _GEN_0; // @[Counter.scala 21:26:@53869.6]
  wire [31:0] _GEN_1; // @[Counter.scala 19:18:@53865.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@53863.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@53864.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@53869.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 19:18:@53865.4]
  assign io_out = count; // @[Counter.scala 25:10:@53872.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@53873.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module AXICmdSplit( // @[:@53875.2]
  input         clock, // @[:@53876.4]
  input         reset, // @[:@53877.4]
  output        io_in_cmd_ready, // @[:@53878.4]
  input         io_in_cmd_valid, // @[:@53878.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@53878.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@53878.4]
  input         io_in_cmd_bits_isWr, // @[:@53878.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@53878.4]
  output        io_in_wdata_ready, // @[:@53878.4]
  input         io_in_wdata_valid, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@53878.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@53878.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@53878.4]
  input         io_in_rresp_ready, // @[:@53878.4]
  input         io_in_wresp_ready, // @[:@53878.4]
  output        io_in_wresp_valid, // @[:@53878.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@53878.4]
  input         io_out_cmd_ready, // @[:@53878.4]
  output        io_out_cmd_valid, // @[:@53878.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@53878.4]
  output [31:0] io_out_cmd_bits_size, // @[:@53878.4]
  output        io_out_cmd_bits_isWr, // @[:@53878.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@53878.4]
  input         io_out_wdata_ready, // @[:@53878.4]
  output        io_out_wdata_valid, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@53878.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@53878.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@53878.4]
  output        io_out_rresp_ready, // @[:@53878.4]
  output        io_out_wresp_ready, // @[:@53878.4]
  input         io_out_wresp_valid, // @[:@53878.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@53878.4]
);
  wire  cmdSizeCounter_clock; // @[AXIProtocol.scala 18:30:@53992.4]
  wire  cmdSizeCounter_reset; // @[AXIProtocol.scala 18:30:@53992.4]
  wire  cmdSizeCounter_io_reset; // @[AXIProtocol.scala 18:30:@53992.4]
  wire  cmdSizeCounter_io_enable; // @[AXIProtocol.scala 18:30:@53992.4]
  wire [31:0] cmdSizeCounter_io_stride; // @[AXIProtocol.scala 18:30:@53992.4]
  wire [31:0] cmdSizeCounter_io_out; // @[AXIProtocol.scala 18:30:@53992.4]
  wire [31:0] cmdSizeCounter_io_next; // @[AXIProtocol.scala 18:30:@53992.4]
  wire [32:0] _T_199; // @[AXIProtocol.scala 20:46:@53995.4]
  wire [32:0] _T_200; // @[AXIProtocol.scala 20:46:@53996.4]
  wire [31:0] cmdSizeRemaining; // @[AXIProtocol.scala 20:46:@53997.4]
  wire  lastCmd; // @[AXIProtocol.scala 23:35:@53998.4]
  wire [37:0] _GEN_0; // @[AXIProtocol.scala 27:47:@54001.4]
  wire [37:0] addrOffsetBytes; // @[AXIProtocol.scala 27:47:@54001.4]
  wire [63:0] _GEN_1; // @[AXIProtocol.scala 28:49:@54002.4]
  wire [64:0] _T_201; // @[AXIProtocol.scala 28:49:@54002.4]
  wire [63:0] cmdAddr_bits; // @[AXIProtocol.scala 28:49:@54003.4]
  wire [57:0] _T_204; // @[FringeBundles.scala 158:22:@54006.4]
  wire [7:0] cmdTag_streamID; // @[FringeBundles.scala 114:28:@54013.4]
  wire [22:0] cmdTag_uid; // @[FringeBundles.scala 114:28:@54017.4]
  wire [23:0] _T_214; // @[FringeBundles.scala 115:37:@54020.4]
  wire  cmdIssue; // @[AXIProtocol.scala 36:35:@54023.4]
  wire  _T_223; // @[FringeBundles.scala 140:28:@54034.4]
  Counter_72 cmdSizeCounter ( // @[AXIProtocol.scala 18:30:@53992.4]
    .clock(cmdSizeCounter_clock),
    .reset(cmdSizeCounter_reset),
    .io_reset(cmdSizeCounter_io_reset),
    .io_enable(cmdSizeCounter_io_enable),
    .io_stride(cmdSizeCounter_io_stride),
    .io_out(cmdSizeCounter_io_out),
    .io_next(cmdSizeCounter_io_next)
  );
  assign _T_199 = io_in_cmd_bits_size - cmdSizeCounter_io_out; // @[AXIProtocol.scala 20:46:@53995.4]
  assign _T_200 = $unsigned(_T_199); // @[AXIProtocol.scala 20:46:@53996.4]
  assign cmdSizeRemaining = _T_200[31:0]; // @[AXIProtocol.scala 20:46:@53997.4]
  assign lastCmd = cmdSizeRemaining <= 32'h100; // @[AXIProtocol.scala 23:35:@53998.4]
  assign _GEN_0 = {{6'd0}, cmdSizeCounter_io_out}; // @[AXIProtocol.scala 27:47:@54001.4]
  assign addrOffsetBytes = _GEN_0 << 6; // @[AXIProtocol.scala 27:47:@54001.4]
  assign _GEN_1 = {{26'd0}, addrOffsetBytes}; // @[AXIProtocol.scala 28:49:@54002.4]
  assign _T_201 = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@54002.4]
  assign cmdAddr_bits = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@54003.4]
  assign _T_204 = cmdAddr_bits[63:6]; // @[FringeBundles.scala 158:22:@54006.4]
  assign cmdTag_streamID = io_in_cmd_bits_tag[7:0]; // @[FringeBundles.scala 114:28:@54013.4]
  assign cmdTag_uid = io_in_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@54017.4]
  assign _T_214 = {cmdTag_uid,lastCmd}; // @[FringeBundles.scala 115:37:@54020.4]
  assign cmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 36:35:@54023.4]
  assign _T_223 = io_out_wresp_bits_tag[8]; // @[FringeBundles.scala 140:28:@54034.4]
  assign io_in_cmd_ready = lastCmd & cmdIssue; // @[AXIProtocol.scala 15:10:@53991.4 AXIProtocol.scala 38:19:@54025.4]
  assign io_in_wdata_ready = io_out_wdata_ready; // @[AXIProtocol.scala 15:10:@53984.4]
  assign io_in_wresp_valid = io_out_wresp_valid & _T_223; // @[AXIProtocol.scala 15:10:@53881.4 AXIProtocol.scala 46:21:@54039.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 15:10:@53880.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 15:10:@53990.4]
  assign io_out_cmd_bits_addr = {_T_204,6'h0}; // @[AXIProtocol.scala 15:10:@53989.4 AXIProtocol.scala 29:24:@54008.4]
  assign io_out_cmd_bits_size = lastCmd ? cmdSizeRemaining : 32'h100; // @[AXIProtocol.scala 15:10:@53988.4 AXIProtocol.scala 25:24:@54000.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 15:10:@53986.4]
  assign io_out_cmd_bits_tag = {_T_214,cmdTag_streamID}; // @[AXIProtocol.scala 15:10:@53985.4 FringeBundles.scala 115:32:@54022.4]
  assign io_out_wdata_valid = io_in_wdata_valid; // @[AXIProtocol.scala 15:10:@53983.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 15:10:@53967.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 15:10:@53968.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 15:10:@53969.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 15:10:@53970.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 15:10:@53971.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 15:10:@53972.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 15:10:@53973.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 15:10:@53974.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 15:10:@53975.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 15:10:@53976.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 15:10:@53977.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 15:10:@53978.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 15:10:@53979.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 15:10:@53980.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 15:10:@53981.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 15:10:@53982.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 15:10:@53903.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 15:10:@53904.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 15:10:@53905.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 15:10:@53906.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 15:10:@53907.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 15:10:@53908.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 15:10:@53909.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 15:10:@53910.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 15:10:@53911.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 15:10:@53912.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 15:10:@53913.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 15:10:@53914.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 15:10:@53915.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 15:10:@53916.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 15:10:@53917.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 15:10:@53918.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 15:10:@53919.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 15:10:@53920.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 15:10:@53921.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 15:10:@53922.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 15:10:@53923.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 15:10:@53924.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 15:10:@53925.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 15:10:@53926.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 15:10:@53927.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 15:10:@53928.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 15:10:@53929.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 15:10:@53930.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 15:10:@53931.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 15:10:@53932.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 15:10:@53933.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 15:10:@53934.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 15:10:@53935.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 15:10:@53936.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 15:10:@53937.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 15:10:@53938.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 15:10:@53939.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 15:10:@53940.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 15:10:@53941.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 15:10:@53942.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 15:10:@53943.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 15:10:@53944.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 15:10:@53945.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 15:10:@53946.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 15:10:@53947.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 15:10:@53948.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 15:10:@53949.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 15:10:@53950.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 15:10:@53951.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 15:10:@53952.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 15:10:@53953.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 15:10:@53954.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 15:10:@53955.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 15:10:@53956.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 15:10:@53957.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 15:10:@53958.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 15:10:@53959.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 15:10:@53960.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 15:10:@53961.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 15:10:@53962.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 15:10:@53963.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 15:10:@53964.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 15:10:@53965.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 15:10:@53966.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 15:10:@53901.4]
  assign io_out_wresp_ready = _T_223 ? io_in_wresp_ready : 1'h1; // @[AXIProtocol.scala 15:10:@53882.4 AXIProtocol.scala 47:22:@54041.4]
  assign cmdSizeCounter_clock = clock; // @[:@53993.4]
  assign cmdSizeCounter_reset = reset; // @[:@53994.4]
  assign cmdSizeCounter_io_reset = lastCmd & cmdIssue; // @[AXIProtocol.scala 40:27:@54026.4]
  assign cmdSizeCounter_io_enable = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 41:28:@54027.4]
  assign cmdSizeCounter_io_stride = 32'h100; // @[AXIProtocol.scala 42:28:@54028.4]
endmodule
module AXICmdIssue( // @[:@54061.2]
  input         clock, // @[:@54062.4]
  input         reset, // @[:@54063.4]
  output        io_in_cmd_ready, // @[:@54064.4]
  input         io_in_cmd_valid, // @[:@54064.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@54064.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@54064.4]
  input         io_in_cmd_bits_isWr, // @[:@54064.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@54064.4]
  output        io_in_wdata_ready, // @[:@54064.4]
  input         io_in_wdata_valid, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@54064.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@54064.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@54064.4]
  input         io_in_rresp_ready, // @[:@54064.4]
  input         io_in_wresp_ready, // @[:@54064.4]
  output        io_in_wresp_valid, // @[:@54064.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@54064.4]
  input         io_out_cmd_ready, // @[:@54064.4]
  output        io_out_cmd_valid, // @[:@54064.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@54064.4]
  output [31:0] io_out_cmd_bits_size, // @[:@54064.4]
  output        io_out_cmd_bits_isWr, // @[:@54064.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@54064.4]
  input         io_out_wdata_ready, // @[:@54064.4]
  output        io_out_wdata_valid, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@54064.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@54064.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@54064.4]
  output        io_out_wdata_bits_wlast, // @[:@54064.4]
  output        io_out_rresp_ready, // @[:@54064.4]
  output        io_out_wresp_ready, // @[:@54064.4]
  input         io_out_wresp_valid, // @[:@54064.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@54064.4]
);
  wire  wdataCounter_clock; // @[AXIProtocol.scala 59:28:@54178.4]
  wire  wdataCounter_reset; // @[AXIProtocol.scala 59:28:@54178.4]
  wire  wdataCounter_io_reset; // @[AXIProtocol.scala 59:28:@54178.4]
  wire  wdataCounter_io_enable; // @[AXIProtocol.scala 59:28:@54178.4]
  wire [31:0] wdataCounter_io_stride; // @[AXIProtocol.scala 59:28:@54178.4]
  wire [31:0] wdataCounter_io_out; // @[AXIProtocol.scala 59:28:@54178.4]
  wire [31:0] wdataCounter_io_next; // @[AXIProtocol.scala 59:28:@54178.4]
  reg  writeIssued; // @[AXIProtocol.scala 61:28:@54181.4]
  reg [31:0] _RAND_0;
  wire  dramCmdIssue; // @[AXIProtocol.scala 63:39:@54182.4]
  wire  dramWriteIssue; // @[AXIProtocol.scala 64:43:@54183.4]
  wire  _T_201; // @[AXIProtocol.scala 68:54:@54184.4]
  wire  wlast; // @[AXIProtocol.scala 68:30:@54185.4]
  wire  _T_203; // @[AXIProtocol.scala 72:28:@54191.6]
  wire  _GEN_0; // @[AXIProtocol.scala 72:40:@54192.6]
  wire  _GEN_1; // @[AXIProtocol.scala 70:15:@54187.4]
  wire  _T_208; // @[AXIProtocol.scala 84:55:@54201.4]
  wire  _T_210; // @[AXIProtocol.scala 84:44:@54202.4]
  Counter_72 wdataCounter ( // @[AXIProtocol.scala 59:28:@54178.4]
    .clock(wdataCounter_clock),
    .reset(wdataCounter_reset),
    .io_reset(wdataCounter_io_reset),
    .io_enable(wdataCounter_io_enable),
    .io_stride(wdataCounter_io_stride),
    .io_out(wdataCounter_io_out),
    .io_next(wdataCounter_io_next)
  );
  assign dramCmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 63:39:@54182.4]
  assign dramWriteIssue = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 64:43:@54183.4]
  assign _T_201 = wdataCounter_io_next == io_in_cmd_bits_size; // @[AXIProtocol.scala 68:54:@54184.4]
  assign wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 68:30:@54185.4]
  assign _T_203 = dramCmdIssue & io_in_cmd_bits_isWr; // @[AXIProtocol.scala 72:28:@54191.6]
  assign _GEN_0 = _T_203 ? 1'h1 : writeIssued; // @[AXIProtocol.scala 72:40:@54192.6]
  assign _GEN_1 = wlast ? 1'h0 : _GEN_0; // @[AXIProtocol.scala 70:15:@54187.4]
  assign _T_208 = writeIssued == 1'h0; // @[AXIProtocol.scala 84:55:@54201.4]
  assign _T_210 = io_in_cmd_bits_isWr ? _T_208 : 1'h1; // @[AXIProtocol.scala 84:44:@54202.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? wlast : dramCmdIssue; // @[AXIProtocol.scala 56:10:@54177.4 AXIProtocol.scala 81:19:@54199.4]
  assign io_in_wdata_ready = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 56:10:@54170.4 AXIProtocol.scala 82:21:@54200.4]
  assign io_in_wresp_valid = io_out_wresp_valid; // @[AXIProtocol.scala 56:10:@54067.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 56:10:@54066.4]
  assign io_out_cmd_valid = io_in_cmd_valid & _T_210; // @[AXIProtocol.scala 56:10:@54176.4 AXIProtocol.scala 84:20:@54204.4]
  assign io_out_cmd_bits_addr = io_in_cmd_bits_addr; // @[AXIProtocol.scala 56:10:@54175.4]
  assign io_out_cmd_bits_size = io_in_cmd_bits_size; // @[AXIProtocol.scala 56:10:@54174.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 56:10:@54172.4]
  assign io_out_cmd_bits_tag = io_in_cmd_bits_tag; // @[AXIProtocol.scala 56:10:@54171.4]
  assign io_out_wdata_valid = io_in_wdata_valid & writeIssued; // @[AXIProtocol.scala 56:10:@54169.4 AXIProtocol.scala 86:22:@54206.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 56:10:@54153.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 56:10:@54154.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 56:10:@54155.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 56:10:@54156.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 56:10:@54157.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 56:10:@54158.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 56:10:@54159.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 56:10:@54160.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 56:10:@54161.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 56:10:@54162.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 56:10:@54163.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 56:10:@54164.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 56:10:@54165.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 56:10:@54166.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 56:10:@54167.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 56:10:@54168.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 56:10:@54089.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 56:10:@54090.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 56:10:@54091.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 56:10:@54092.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 56:10:@54093.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 56:10:@54094.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 56:10:@54095.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 56:10:@54096.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 56:10:@54097.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 56:10:@54098.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 56:10:@54099.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 56:10:@54100.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 56:10:@54101.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 56:10:@54102.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 56:10:@54103.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 56:10:@54104.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 56:10:@54105.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 56:10:@54106.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 56:10:@54107.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 56:10:@54108.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 56:10:@54109.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 56:10:@54110.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 56:10:@54111.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 56:10:@54112.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 56:10:@54113.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 56:10:@54114.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 56:10:@54115.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 56:10:@54116.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 56:10:@54117.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 56:10:@54118.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 56:10:@54119.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 56:10:@54120.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 56:10:@54121.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 56:10:@54122.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 56:10:@54123.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 56:10:@54124.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 56:10:@54125.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 56:10:@54126.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 56:10:@54127.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 56:10:@54128.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 56:10:@54129.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 56:10:@54130.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 56:10:@54131.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 56:10:@54132.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 56:10:@54133.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 56:10:@54134.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 56:10:@54135.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 56:10:@54136.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 56:10:@54137.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 56:10:@54138.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 56:10:@54139.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 56:10:@54140.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 56:10:@54141.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 56:10:@54142.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 56:10:@54143.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 56:10:@54144.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 56:10:@54145.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 56:10:@54146.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 56:10:@54147.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 56:10:@54148.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 56:10:@54149.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 56:10:@54150.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 56:10:@54151.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 56:10:@54152.4]
  assign io_out_wdata_bits_wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 56:10:@54088.4 AXIProtocol.scala 87:27:@54207.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 56:10:@54087.4]
  assign io_out_wresp_ready = io_in_wresp_ready; // @[AXIProtocol.scala 56:10:@54068.4]
  assign wdataCounter_clock = clock; // @[:@54179.4]
  assign wdataCounter_reset = reset; // @[:@54180.4]
  assign wdataCounter_io_reset = dramWriteIssue & _T_201; // @[AXIProtocol.scala 76:25:@54195.4]
  assign wdataCounter_io_enable = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 77:26:@54196.4]
  assign wdataCounter_io_stride = 32'h1; // @[AXIProtocol.scala 78:26:@54197.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeIssued = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      writeIssued <= 1'h0;
    end else begin
      if (wlast) begin
        writeIssued <= 1'h0;
      end else begin
        if (_T_203) begin
          writeIssued <= 1'h1;
        end
      end
    end
  end
endmodule
module DRAMArbiter( // @[:@54209.2]
  input         clock, // @[:@54210.4]
  input         reset, // @[:@54211.4]
  input         io_enable, // @[:@54212.4]
  output        io_app_stores_0_cmd_ready, // @[:@54212.4]
  input         io_app_stores_0_cmd_valid, // @[:@54212.4]
  input  [63:0] io_app_stores_0_cmd_bits_addr, // @[:@54212.4]
  input  [31:0] io_app_stores_0_cmd_bits_size, // @[:@54212.4]
  output        io_app_stores_0_data_ready, // @[:@54212.4]
  input         io_app_stores_0_data_valid, // @[:@54212.4]
  input  [31:0] io_app_stores_0_data_bits_wdata_0, // @[:@54212.4]
  input         io_app_stores_0_data_bits_wstrb, // @[:@54212.4]
  input         io_app_stores_0_wresp_ready, // @[:@54212.4]
  output        io_app_stores_0_wresp_valid, // @[:@54212.4]
  output        io_app_stores_0_wresp_bits, // @[:@54212.4]
  input         io_dram_cmd_ready, // @[:@54212.4]
  output        io_dram_cmd_valid, // @[:@54212.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@54212.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@54212.4]
  output        io_dram_cmd_bits_isWr, // @[:@54212.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@54212.4]
  input         io_dram_wdata_ready, // @[:@54212.4]
  output        io_dram_wdata_valid, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@54212.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@54212.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@54212.4]
  output        io_dram_wdata_bits_wlast, // @[:@54212.4]
  output        io_dram_rresp_ready, // @[:@54212.4]
  output        io_dram_wresp_ready, // @[:@54212.4]
  input         io_dram_wresp_valid, // @[:@54212.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@54212.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@55098.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@55112.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@55340.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@55455.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@55455.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@55098.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@55112.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@55340.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@55455.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_app_stores_0_cmd_ready = StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 68:18:@55111.4]
  assign io_app_stores_0_data_ready = StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 68:18:@55107.4]
  assign io_app_stores_0_wresp_valid = StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 68:18:@55102.4]
  assign io_app_stores_0_wresp_bits = StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 68:18:@55101.4]
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@55680.4 DRAMArbiter.scala 100:23:@55683.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@55679.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@55678.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@55676.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@55675.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@55673.4 DRAMArbiter.scala 101:25:@55685.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@55657.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@55658.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@55659.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@55660.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@55661.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@55662.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@55663.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@55664.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@55665.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@55666.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@55667.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@55668.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@55669.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@55670.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@55671.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@55672.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@55593.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@55594.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@55595.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@55596.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@55597.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@55598.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@55599.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@55600.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@55601.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@55602.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@55603.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@55604.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@55605.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@55606.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@55607.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@55608.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@55609.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@55610.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@55611.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@55612.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@55613.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@55614.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@55615.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@55616.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@55617.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@55618.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@55619.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@55620.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@55621.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@55622.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@55623.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@55624.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@55625.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@55626.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@55627.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@55628.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@55629.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@55630.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@55631.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@55632.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@55633.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@55634.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@55635.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@55636.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@55637.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@55638.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@55639.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@55640.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@55641.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@55642.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@55643.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@55644.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@55645.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@55646.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@55647.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@55648.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@55649.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@55650.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@55651.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@55652.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@55653.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@55654.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@55655.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@55656.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@55592.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@55591.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@55572.4]
  assign StreamControllerStore_clock = clock; // @[:@55099.4]
  assign StreamControllerStore_reset = reset; // @[:@55100.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@55227.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@55220.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@55117.4]
  assign StreamControllerStore_io_store_cmd_valid = io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 68:18:@55110.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = io_app_stores_0_cmd_bits_addr; // @[DRAMArbiter.scala 68:18:@55109.4]
  assign StreamControllerStore_io_store_cmd_bits_size = io_app_stores_0_cmd_bits_size; // @[DRAMArbiter.scala 68:18:@55108.4]
  assign StreamControllerStore_io_store_data_valid = io_app_stores_0_data_valid; // @[DRAMArbiter.scala 68:18:@55106.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = io_app_stores_0_data_bits_wdata_0; // @[DRAMArbiter.scala 68:18:@55105.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = io_app_stores_0_data_bits_wstrb; // @[DRAMArbiter.scala 68:18:@55104.4]
  assign StreamControllerStore_io_store_wresp_ready = io_app_stores_0_wresp_ready; // @[DRAMArbiter.scala 68:18:@55103.4]
  assign StreamArbiter_clock = clock; // @[:@55113.4]
  assign StreamArbiter_reset = reset; // @[:@55114.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@55338.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@55337.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@55336.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@55334.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@55333.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@55331.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@55315.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@55316.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@55317.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@55318.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@55319.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@55320.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@55321.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@55322.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@55323.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@55324.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@55325.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@55326.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@55327.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@55328.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@55329.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@55330.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@55251.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@55252.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@55253.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@55254.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@55255.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@55256.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@55257.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@55258.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@55259.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@55260.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@55261.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@55262.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@55263.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@55264.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@55265.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@55266.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@55267.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@55268.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@55269.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@55270.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@55271.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@55272.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@55273.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@55274.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@55275.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@55276.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@55277.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@55278.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@55279.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@55280.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@55281.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@55282.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@55283.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@55284.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@55285.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@55286.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@55287.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@55288.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@55289.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@55290.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@55291.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@55292.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@55293.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@55294.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@55295.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@55296.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@55297.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@55298.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@55299.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@55300.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@55301.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@55302.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@55303.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@55304.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@55305.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@55306.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@55307.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@55308.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@55309.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@55310.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@55311.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@55312.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@55313.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@55314.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@55249.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@55230.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@55454.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@55447.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@55344.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@55343.4]
  assign AXICmdSplit_clock = clock; // @[:@55341.4]
  assign AXICmdSplit_reset = reset; // @[:@55342.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@55453.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@55452.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@55451.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@55449.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@55448.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@55446.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@55430.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@55431.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@55432.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@55433.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@55434.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@55435.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@55436.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@55437.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@55438.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@55439.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@55440.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@55441.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@55442.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@55443.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@55444.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@55445.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@55366.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@55367.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@55368.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@55369.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@55370.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@55371.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@55372.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@55373.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@55374.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@55375.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@55376.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@55377.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@55378.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@55379.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@55380.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@55381.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@55382.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@55383.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@55384.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@55385.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@55386.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@55387.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@55388.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@55389.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@55390.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@55391.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@55392.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@55393.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@55394.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@55395.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@55396.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@55397.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@55398.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@55399.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@55400.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@55401.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@55402.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@55403.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@55404.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@55405.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@55406.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@55407.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@55408.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@55409.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@55410.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@55411.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@55412.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@55413.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@55414.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@55415.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@55416.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@55417.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@55418.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@55419.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@55420.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@55421.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@55422.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@55423.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@55424.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@55425.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@55426.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@55427.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@55428.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@55429.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@55364.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@55345.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@55569.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@55562.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@55459.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@55458.4]
  assign AXICmdIssue_clock = clock; // @[:@55456.4]
  assign AXICmdIssue_reset = reset; // @[:@55457.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@55568.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@55567.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@55566.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@55564.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@55563.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@55561.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@55545.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@55546.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@55547.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@55548.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@55549.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@55550.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@55551.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@55552.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@55553.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@55554.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@55555.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@55556.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@55557.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@55558.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@55559.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@55560.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@55481.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@55482.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@55483.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@55484.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@55485.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@55486.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@55487.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@55488.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@55489.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@55490.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@55491.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@55492.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@55493.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@55494.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@55495.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@55496.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@55497.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@55498.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@55499.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@55500.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@55501.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@55502.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@55503.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@55504.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@55505.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@55506.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@55507.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@55508.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@55509.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@55510.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@55511.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@55512.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@55513.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@55514.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@55515.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@55516.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@55517.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@55518.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@55519.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@55520.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@55521.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@55522.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@55523.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@55524.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@55525.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@55526.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@55527.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@55528.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@55529.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@55530.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@55531.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@55532.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@55533.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@55534.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@55535.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@55536.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@55537.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@55538.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@55539.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@55540.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@55541.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@55542.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@55543.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@55544.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@55479.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@55460.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@55681.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@55674.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@55571.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@55570.4]
endmodule
module DRAMArbiter_1( // @[:@69910.2]
  input         clock, // @[:@69911.4]
  input         reset, // @[:@69912.4]
  input         io_enable, // @[:@69913.4]
  input         io_dram_cmd_ready, // @[:@69913.4]
  output        io_dram_cmd_valid, // @[:@69913.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@69913.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@69913.4]
  output        io_dram_cmd_bits_isWr, // @[:@69913.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@69913.4]
  input         io_dram_wdata_ready, // @[:@69913.4]
  output        io_dram_wdata_valid, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@69913.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@69913.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@69913.4]
  output        io_dram_wdata_bits_wlast, // @[:@69913.4]
  output        io_dram_rresp_ready, // @[:@69913.4]
  output        io_dram_wresp_ready, // @[:@69913.4]
  input         io_dram_wresp_valid, // @[:@69913.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@69913.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@70799.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@70813.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@71041.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@71156.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@71156.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@70799.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@70813.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@71041.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@71156.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@71381.4 DRAMArbiter.scala 100:23:@71384.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@71380.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@71379.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@71377.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@71376.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@71374.4 DRAMArbiter.scala 101:25:@71386.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@71358.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@71359.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@71360.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@71361.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@71362.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@71363.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@71364.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@71365.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@71366.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@71367.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@71368.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@71369.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@71370.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@71371.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@71372.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@71373.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@71294.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@71295.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@71296.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@71297.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@71298.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@71299.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@71300.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@71301.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@71302.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@71303.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@71304.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@71305.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@71306.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@71307.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@71308.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@71309.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@71310.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@71311.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@71312.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@71313.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@71314.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@71315.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@71316.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@71317.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@71318.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@71319.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@71320.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@71321.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@71322.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@71323.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@71324.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@71325.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@71326.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@71327.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@71328.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@71329.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@71330.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@71331.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@71332.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@71333.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@71334.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@71335.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@71336.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@71337.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@71338.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@71339.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@71340.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@71341.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@71342.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@71343.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@71344.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@71345.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@71346.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@71347.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@71348.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@71349.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@71350.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@71351.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@71352.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@71353.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@71354.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@71355.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@71356.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@71357.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@71293.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@71292.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@71273.4]
  assign StreamControllerStore_clock = clock; // @[:@70800.4]
  assign StreamControllerStore_reset = reset; // @[:@70801.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@70928.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@70921.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@70818.4]
  assign StreamControllerStore_io_store_cmd_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@70811.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = 64'h0; // @[DRAMArbiter.scala 68:18:@70810.4]
  assign StreamControllerStore_io_store_cmd_bits_size = 32'h0; // @[DRAMArbiter.scala 68:18:@70809.4]
  assign StreamControllerStore_io_store_data_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@70807.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = 32'h0; // @[DRAMArbiter.scala 68:18:@70806.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = 1'h0; // @[DRAMArbiter.scala 68:18:@70805.4]
  assign StreamControllerStore_io_store_wresp_ready = 1'h0; // @[DRAMArbiter.scala 68:18:@70804.4]
  assign StreamArbiter_clock = clock; // @[:@70814.4]
  assign StreamArbiter_reset = reset; // @[:@70815.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@71039.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@71038.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@71037.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@71035.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@71034.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@71032.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@71016.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@71017.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@71018.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@71019.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@71020.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@71021.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@71022.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@71023.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@71024.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@71025.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@71026.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@71027.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@71028.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@71029.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@71030.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@71031.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@70952.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@70953.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@70954.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@70955.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@70956.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@70957.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@70958.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@70959.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@70960.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@70961.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@70962.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@70963.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@70964.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@70965.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@70966.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@70967.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@70968.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@70969.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@70970.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@70971.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@70972.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@70973.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@70974.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@70975.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@70976.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@70977.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@70978.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@70979.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@70980.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@70981.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@70982.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@70983.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@70984.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@70985.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@70986.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@70987.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@70988.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@70989.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@70990.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@70991.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@70992.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@70993.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@70994.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@70995.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@70996.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@70997.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@70998.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@70999.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@71000.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@71001.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@71002.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@71003.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@71004.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@71005.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@71006.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@71007.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@71008.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@71009.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@71010.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@71011.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@71012.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@71013.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@71014.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@71015.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@70950.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@70931.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@71155.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@71148.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@71045.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@71044.4]
  assign AXICmdSplit_clock = clock; // @[:@71042.4]
  assign AXICmdSplit_reset = reset; // @[:@71043.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@71154.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@71153.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@71152.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@71150.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@71149.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@71147.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@71131.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@71132.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@71133.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@71134.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@71135.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@71136.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@71137.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@71138.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@71139.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@71140.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@71141.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@71142.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@71143.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@71144.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@71145.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@71146.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@71067.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@71068.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@71069.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@71070.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@71071.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@71072.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@71073.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@71074.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@71075.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@71076.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@71077.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@71078.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@71079.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@71080.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@71081.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@71082.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@71083.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@71084.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@71085.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@71086.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@71087.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@71088.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@71089.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@71090.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@71091.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@71092.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@71093.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@71094.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@71095.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@71096.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@71097.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@71098.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@71099.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@71100.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@71101.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@71102.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@71103.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@71104.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@71105.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@71106.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@71107.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@71108.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@71109.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@71110.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@71111.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@71112.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@71113.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@71114.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@71115.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@71116.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@71117.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@71118.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@71119.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@71120.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@71121.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@71122.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@71123.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@71124.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@71125.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@71126.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@71127.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@71128.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@71129.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@71130.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@71065.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@71046.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@71270.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@71263.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@71160.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@71159.4]
  assign AXICmdIssue_clock = clock; // @[:@71157.4]
  assign AXICmdIssue_reset = reset; // @[:@71158.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@71269.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@71268.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@71267.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@71265.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@71264.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@71262.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@71246.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@71247.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@71248.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@71249.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@71250.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@71251.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@71252.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@71253.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@71254.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@71255.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@71256.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@71257.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@71258.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@71259.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@71260.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@71261.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@71182.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@71183.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@71184.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@71185.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@71186.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@71187.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@71188.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@71189.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@71190.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@71191.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@71192.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@71193.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@71194.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@71195.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@71196.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@71197.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@71198.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@71199.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@71200.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@71201.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@71202.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@71203.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@71204.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@71205.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@71206.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@71207.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@71208.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@71209.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@71210.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@71211.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@71212.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@71213.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@71214.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@71215.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@71216.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@71217.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@71218.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@71219.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@71220.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@71221.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@71222.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@71223.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@71224.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@71225.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@71226.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@71227.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@71228.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@71229.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@71230.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@71231.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@71232.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@71233.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@71234.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@71235.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@71236.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@71237.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@71238.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@71239.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@71240.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@71241.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@71242.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@71243.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@71244.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@71245.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@71180.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@71161.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@71382.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@71375.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@71272.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@71271.4]
endmodule
module DRAMHeap( // @[:@102018.2]
  input         io_accel_0_req_valid, // @[:@102021.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@102021.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@102021.4]
  output        io_accel_0_resp_valid, // @[:@102021.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@102021.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@102021.4]
  output        io_host_0_req_valid, // @[:@102021.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@102021.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@102021.4]
  input         io_host_0_resp_valid, // @[:@102021.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@102021.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@102021.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@102028.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@102030.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@102029.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@102025.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@102024.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@102023.4]
endmodule
module RetimeWrapper_424( // @[:@102044.2]
  input         clock, // @[:@102045.4]
  input         reset, // @[:@102046.4]
  input         io_flow, // @[:@102047.4]
  input  [63:0] io_in, // @[:@102047.4]
  output [63:0] io_out // @[:@102047.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@102049.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@102049.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@102049.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@102049.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@102049.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@102049.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@102049.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@102062.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@102061.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@102060.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@102059.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@102058.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@102056.4]
endmodule
module FringeFF( // @[:@102064.2]
  input         clock, // @[:@102065.4]
  input         reset, // @[:@102066.4]
  input  [63:0] io_in, // @[:@102067.4]
  input         io_reset, // @[:@102067.4]
  output [63:0] io_out, // @[:@102067.4]
  input         io_enable // @[:@102067.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@102070.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@102070.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@102070.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@102070.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@102070.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@102075.4 package.scala 96:25:@102076.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@102081.6]
  RetimeWrapper_424 RetimeWrapper ( // @[package.scala 93:22:@102070.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@102075.4 package.scala 96:25:@102076.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@102081.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@102087.4]
  assign RetimeWrapper_clock = clock; // @[:@102071.4]
  assign RetimeWrapper_reset = reset; // @[:@102072.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@102074.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@102073.4]
endmodule
module MuxN( // @[:@130703.2]
  input  [63:0] io_ins_0, // @[:@130706.4]
  input  [63:0] io_ins_1, // @[:@130706.4]
  input  [63:0] io_ins_2, // @[:@130706.4]
  input  [63:0] io_ins_3, // @[:@130706.4]
  input  [63:0] io_ins_4, // @[:@130706.4]
  input  [63:0] io_ins_5, // @[:@130706.4]
  input  [63:0] io_ins_6, // @[:@130706.4]
  input  [63:0] io_ins_7, // @[:@130706.4]
  input  [63:0] io_ins_8, // @[:@130706.4]
  input  [63:0] io_ins_9, // @[:@130706.4]
  input  [63:0] io_ins_10, // @[:@130706.4]
  input  [63:0] io_ins_11, // @[:@130706.4]
  input  [63:0] io_ins_12, // @[:@130706.4]
  input  [63:0] io_ins_13, // @[:@130706.4]
  input  [63:0] io_ins_14, // @[:@130706.4]
  input  [63:0] io_ins_15, // @[:@130706.4]
  input  [63:0] io_ins_16, // @[:@130706.4]
  input  [63:0] io_ins_17, // @[:@130706.4]
  input  [63:0] io_ins_18, // @[:@130706.4]
  input  [63:0] io_ins_19, // @[:@130706.4]
  input  [63:0] io_ins_20, // @[:@130706.4]
  input  [63:0] io_ins_21, // @[:@130706.4]
  input  [63:0] io_ins_22, // @[:@130706.4]
  input  [63:0] io_ins_23, // @[:@130706.4]
  input  [63:0] io_ins_24, // @[:@130706.4]
  input  [63:0] io_ins_25, // @[:@130706.4]
  input  [63:0] io_ins_26, // @[:@130706.4]
  input  [63:0] io_ins_27, // @[:@130706.4]
  input  [63:0] io_ins_28, // @[:@130706.4]
  input  [63:0] io_ins_29, // @[:@130706.4]
  input  [63:0] io_ins_30, // @[:@130706.4]
  input  [63:0] io_ins_31, // @[:@130706.4]
  input  [63:0] io_ins_32, // @[:@130706.4]
  input  [63:0] io_ins_33, // @[:@130706.4]
  input  [63:0] io_ins_34, // @[:@130706.4]
  input  [63:0] io_ins_35, // @[:@130706.4]
  input  [63:0] io_ins_36, // @[:@130706.4]
  input  [63:0] io_ins_37, // @[:@130706.4]
  input  [63:0] io_ins_38, // @[:@130706.4]
  input  [63:0] io_ins_39, // @[:@130706.4]
  input  [63:0] io_ins_40, // @[:@130706.4]
  input  [63:0] io_ins_41, // @[:@130706.4]
  input  [63:0] io_ins_42, // @[:@130706.4]
  input  [63:0] io_ins_43, // @[:@130706.4]
  input  [63:0] io_ins_44, // @[:@130706.4]
  input  [63:0] io_ins_45, // @[:@130706.4]
  input  [63:0] io_ins_46, // @[:@130706.4]
  input  [63:0] io_ins_47, // @[:@130706.4]
  input  [63:0] io_ins_48, // @[:@130706.4]
  input  [63:0] io_ins_49, // @[:@130706.4]
  input  [63:0] io_ins_50, // @[:@130706.4]
  input  [63:0] io_ins_51, // @[:@130706.4]
  input  [63:0] io_ins_52, // @[:@130706.4]
  input  [63:0] io_ins_53, // @[:@130706.4]
  input  [63:0] io_ins_54, // @[:@130706.4]
  input  [63:0] io_ins_55, // @[:@130706.4]
  input  [63:0] io_ins_56, // @[:@130706.4]
  input  [63:0] io_ins_57, // @[:@130706.4]
  input  [63:0] io_ins_58, // @[:@130706.4]
  input  [63:0] io_ins_59, // @[:@130706.4]
  input  [63:0] io_ins_60, // @[:@130706.4]
  input  [63:0] io_ins_61, // @[:@130706.4]
  input  [63:0] io_ins_62, // @[:@130706.4]
  input  [63:0] io_ins_63, // @[:@130706.4]
  input  [63:0] io_ins_64, // @[:@130706.4]
  input  [63:0] io_ins_65, // @[:@130706.4]
  input  [63:0] io_ins_66, // @[:@130706.4]
  input  [63:0] io_ins_67, // @[:@130706.4]
  input  [63:0] io_ins_68, // @[:@130706.4]
  input  [63:0] io_ins_69, // @[:@130706.4]
  input  [63:0] io_ins_70, // @[:@130706.4]
  input  [63:0] io_ins_71, // @[:@130706.4]
  input  [63:0] io_ins_72, // @[:@130706.4]
  input  [63:0] io_ins_73, // @[:@130706.4]
  input  [63:0] io_ins_74, // @[:@130706.4]
  input  [63:0] io_ins_75, // @[:@130706.4]
  input  [63:0] io_ins_76, // @[:@130706.4]
  input  [63:0] io_ins_77, // @[:@130706.4]
  input  [63:0] io_ins_78, // @[:@130706.4]
  input  [63:0] io_ins_79, // @[:@130706.4]
  input  [63:0] io_ins_80, // @[:@130706.4]
  input  [63:0] io_ins_81, // @[:@130706.4]
  input  [63:0] io_ins_82, // @[:@130706.4]
  input  [63:0] io_ins_83, // @[:@130706.4]
  input  [63:0] io_ins_84, // @[:@130706.4]
  input  [63:0] io_ins_85, // @[:@130706.4]
  input  [63:0] io_ins_86, // @[:@130706.4]
  input  [63:0] io_ins_87, // @[:@130706.4]
  input  [63:0] io_ins_88, // @[:@130706.4]
  input  [63:0] io_ins_89, // @[:@130706.4]
  input  [63:0] io_ins_90, // @[:@130706.4]
  input  [63:0] io_ins_91, // @[:@130706.4]
  input  [63:0] io_ins_92, // @[:@130706.4]
  input  [63:0] io_ins_93, // @[:@130706.4]
  input  [63:0] io_ins_94, // @[:@130706.4]
  input  [63:0] io_ins_95, // @[:@130706.4]
  input  [63:0] io_ins_96, // @[:@130706.4]
  input  [63:0] io_ins_97, // @[:@130706.4]
  input  [63:0] io_ins_98, // @[:@130706.4]
  input  [63:0] io_ins_99, // @[:@130706.4]
  input  [63:0] io_ins_100, // @[:@130706.4]
  input  [63:0] io_ins_101, // @[:@130706.4]
  input  [63:0] io_ins_102, // @[:@130706.4]
  input  [63:0] io_ins_103, // @[:@130706.4]
  input  [63:0] io_ins_104, // @[:@130706.4]
  input  [63:0] io_ins_105, // @[:@130706.4]
  input  [63:0] io_ins_106, // @[:@130706.4]
  input  [63:0] io_ins_107, // @[:@130706.4]
  input  [63:0] io_ins_108, // @[:@130706.4]
  input  [63:0] io_ins_109, // @[:@130706.4]
  input  [63:0] io_ins_110, // @[:@130706.4]
  input  [63:0] io_ins_111, // @[:@130706.4]
  input  [63:0] io_ins_112, // @[:@130706.4]
  input  [63:0] io_ins_113, // @[:@130706.4]
  input  [63:0] io_ins_114, // @[:@130706.4]
  input  [63:0] io_ins_115, // @[:@130706.4]
  input  [63:0] io_ins_116, // @[:@130706.4]
  input  [63:0] io_ins_117, // @[:@130706.4]
  input  [63:0] io_ins_118, // @[:@130706.4]
  input  [63:0] io_ins_119, // @[:@130706.4]
  input  [63:0] io_ins_120, // @[:@130706.4]
  input  [63:0] io_ins_121, // @[:@130706.4]
  input  [63:0] io_ins_122, // @[:@130706.4]
  input  [63:0] io_ins_123, // @[:@130706.4]
  input  [63:0] io_ins_124, // @[:@130706.4]
  input  [63:0] io_ins_125, // @[:@130706.4]
  input  [63:0] io_ins_126, // @[:@130706.4]
  input  [63:0] io_ins_127, // @[:@130706.4]
  input  [63:0] io_ins_128, // @[:@130706.4]
  input  [63:0] io_ins_129, // @[:@130706.4]
  input  [63:0] io_ins_130, // @[:@130706.4]
  input  [63:0] io_ins_131, // @[:@130706.4]
  input  [63:0] io_ins_132, // @[:@130706.4]
  input  [63:0] io_ins_133, // @[:@130706.4]
  input  [63:0] io_ins_134, // @[:@130706.4]
  input  [63:0] io_ins_135, // @[:@130706.4]
  input  [63:0] io_ins_136, // @[:@130706.4]
  input  [63:0] io_ins_137, // @[:@130706.4]
  input  [63:0] io_ins_138, // @[:@130706.4]
  input  [63:0] io_ins_139, // @[:@130706.4]
  input  [63:0] io_ins_140, // @[:@130706.4]
  input  [63:0] io_ins_141, // @[:@130706.4]
  input  [63:0] io_ins_142, // @[:@130706.4]
  input  [63:0] io_ins_143, // @[:@130706.4]
  input  [63:0] io_ins_144, // @[:@130706.4]
  input  [63:0] io_ins_145, // @[:@130706.4]
  input  [63:0] io_ins_146, // @[:@130706.4]
  input  [63:0] io_ins_147, // @[:@130706.4]
  input  [63:0] io_ins_148, // @[:@130706.4]
  input  [63:0] io_ins_149, // @[:@130706.4]
  input  [63:0] io_ins_150, // @[:@130706.4]
  input  [63:0] io_ins_151, // @[:@130706.4]
  input  [63:0] io_ins_152, // @[:@130706.4]
  input  [63:0] io_ins_153, // @[:@130706.4]
  input  [63:0] io_ins_154, // @[:@130706.4]
  input  [63:0] io_ins_155, // @[:@130706.4]
  input  [63:0] io_ins_156, // @[:@130706.4]
  input  [63:0] io_ins_157, // @[:@130706.4]
  input  [63:0] io_ins_158, // @[:@130706.4]
  input  [63:0] io_ins_159, // @[:@130706.4]
  input  [63:0] io_ins_160, // @[:@130706.4]
  input  [63:0] io_ins_161, // @[:@130706.4]
  input  [63:0] io_ins_162, // @[:@130706.4]
  input  [63:0] io_ins_163, // @[:@130706.4]
  input  [63:0] io_ins_164, // @[:@130706.4]
  input  [63:0] io_ins_165, // @[:@130706.4]
  input  [63:0] io_ins_166, // @[:@130706.4]
  input  [63:0] io_ins_167, // @[:@130706.4]
  input  [63:0] io_ins_168, // @[:@130706.4]
  input  [63:0] io_ins_169, // @[:@130706.4]
  input  [63:0] io_ins_170, // @[:@130706.4]
  input  [63:0] io_ins_171, // @[:@130706.4]
  input  [63:0] io_ins_172, // @[:@130706.4]
  input  [63:0] io_ins_173, // @[:@130706.4]
  input  [63:0] io_ins_174, // @[:@130706.4]
  input  [63:0] io_ins_175, // @[:@130706.4]
  input  [63:0] io_ins_176, // @[:@130706.4]
  input  [63:0] io_ins_177, // @[:@130706.4]
  input  [63:0] io_ins_178, // @[:@130706.4]
  input  [63:0] io_ins_179, // @[:@130706.4]
  input  [63:0] io_ins_180, // @[:@130706.4]
  input  [63:0] io_ins_181, // @[:@130706.4]
  input  [63:0] io_ins_182, // @[:@130706.4]
  input  [63:0] io_ins_183, // @[:@130706.4]
  input  [63:0] io_ins_184, // @[:@130706.4]
  input  [63:0] io_ins_185, // @[:@130706.4]
  input  [63:0] io_ins_186, // @[:@130706.4]
  input  [63:0] io_ins_187, // @[:@130706.4]
  input  [63:0] io_ins_188, // @[:@130706.4]
  input  [63:0] io_ins_189, // @[:@130706.4]
  input  [63:0] io_ins_190, // @[:@130706.4]
  input  [63:0] io_ins_191, // @[:@130706.4]
  input  [63:0] io_ins_192, // @[:@130706.4]
  input  [63:0] io_ins_193, // @[:@130706.4]
  input  [63:0] io_ins_194, // @[:@130706.4]
  input  [63:0] io_ins_195, // @[:@130706.4]
  input  [63:0] io_ins_196, // @[:@130706.4]
  input  [63:0] io_ins_197, // @[:@130706.4]
  input  [63:0] io_ins_198, // @[:@130706.4]
  input  [63:0] io_ins_199, // @[:@130706.4]
  input  [63:0] io_ins_200, // @[:@130706.4]
  input  [63:0] io_ins_201, // @[:@130706.4]
  input  [63:0] io_ins_202, // @[:@130706.4]
  input  [63:0] io_ins_203, // @[:@130706.4]
  input  [63:0] io_ins_204, // @[:@130706.4]
  input  [63:0] io_ins_205, // @[:@130706.4]
  input  [63:0] io_ins_206, // @[:@130706.4]
  input  [63:0] io_ins_207, // @[:@130706.4]
  input  [63:0] io_ins_208, // @[:@130706.4]
  input  [63:0] io_ins_209, // @[:@130706.4]
  input  [63:0] io_ins_210, // @[:@130706.4]
  input  [63:0] io_ins_211, // @[:@130706.4]
  input  [63:0] io_ins_212, // @[:@130706.4]
  input  [63:0] io_ins_213, // @[:@130706.4]
  input  [63:0] io_ins_214, // @[:@130706.4]
  input  [63:0] io_ins_215, // @[:@130706.4]
  input  [63:0] io_ins_216, // @[:@130706.4]
  input  [63:0] io_ins_217, // @[:@130706.4]
  input  [63:0] io_ins_218, // @[:@130706.4]
  input  [63:0] io_ins_219, // @[:@130706.4]
  input  [63:0] io_ins_220, // @[:@130706.4]
  input  [63:0] io_ins_221, // @[:@130706.4]
  input  [63:0] io_ins_222, // @[:@130706.4]
  input  [63:0] io_ins_223, // @[:@130706.4]
  input  [63:0] io_ins_224, // @[:@130706.4]
  input  [63:0] io_ins_225, // @[:@130706.4]
  input  [63:0] io_ins_226, // @[:@130706.4]
  input  [63:0] io_ins_227, // @[:@130706.4]
  input  [63:0] io_ins_228, // @[:@130706.4]
  input  [63:0] io_ins_229, // @[:@130706.4]
  input  [63:0] io_ins_230, // @[:@130706.4]
  input  [63:0] io_ins_231, // @[:@130706.4]
  input  [63:0] io_ins_232, // @[:@130706.4]
  input  [63:0] io_ins_233, // @[:@130706.4]
  input  [63:0] io_ins_234, // @[:@130706.4]
  input  [63:0] io_ins_235, // @[:@130706.4]
  input  [63:0] io_ins_236, // @[:@130706.4]
  input  [63:0] io_ins_237, // @[:@130706.4]
  input  [63:0] io_ins_238, // @[:@130706.4]
  input  [63:0] io_ins_239, // @[:@130706.4]
  input  [63:0] io_ins_240, // @[:@130706.4]
  input  [63:0] io_ins_241, // @[:@130706.4]
  input  [63:0] io_ins_242, // @[:@130706.4]
  input  [63:0] io_ins_243, // @[:@130706.4]
  input  [63:0] io_ins_244, // @[:@130706.4]
  input  [63:0] io_ins_245, // @[:@130706.4]
  input  [63:0] io_ins_246, // @[:@130706.4]
  input  [63:0] io_ins_247, // @[:@130706.4]
  input  [63:0] io_ins_248, // @[:@130706.4]
  input  [63:0] io_ins_249, // @[:@130706.4]
  input  [63:0] io_ins_250, // @[:@130706.4]
  input  [63:0] io_ins_251, // @[:@130706.4]
  input  [63:0] io_ins_252, // @[:@130706.4]
  input  [63:0] io_ins_253, // @[:@130706.4]
  input  [63:0] io_ins_254, // @[:@130706.4]
  input  [63:0] io_ins_255, // @[:@130706.4]
  input  [63:0] io_ins_256, // @[:@130706.4]
  input  [63:0] io_ins_257, // @[:@130706.4]
  input  [63:0] io_ins_258, // @[:@130706.4]
  input  [63:0] io_ins_259, // @[:@130706.4]
  input  [63:0] io_ins_260, // @[:@130706.4]
  input  [63:0] io_ins_261, // @[:@130706.4]
  input  [63:0] io_ins_262, // @[:@130706.4]
  input  [63:0] io_ins_263, // @[:@130706.4]
  input  [63:0] io_ins_264, // @[:@130706.4]
  input  [63:0] io_ins_265, // @[:@130706.4]
  input  [63:0] io_ins_266, // @[:@130706.4]
  input  [63:0] io_ins_267, // @[:@130706.4]
  input  [63:0] io_ins_268, // @[:@130706.4]
  input  [63:0] io_ins_269, // @[:@130706.4]
  input  [63:0] io_ins_270, // @[:@130706.4]
  input  [63:0] io_ins_271, // @[:@130706.4]
  input  [63:0] io_ins_272, // @[:@130706.4]
  input  [63:0] io_ins_273, // @[:@130706.4]
  input  [63:0] io_ins_274, // @[:@130706.4]
  input  [63:0] io_ins_275, // @[:@130706.4]
  input  [63:0] io_ins_276, // @[:@130706.4]
  input  [63:0] io_ins_277, // @[:@130706.4]
  input  [63:0] io_ins_278, // @[:@130706.4]
  input  [63:0] io_ins_279, // @[:@130706.4]
  input  [63:0] io_ins_280, // @[:@130706.4]
  input  [63:0] io_ins_281, // @[:@130706.4]
  input  [63:0] io_ins_282, // @[:@130706.4]
  input  [63:0] io_ins_283, // @[:@130706.4]
  input  [63:0] io_ins_284, // @[:@130706.4]
  input  [63:0] io_ins_285, // @[:@130706.4]
  input  [63:0] io_ins_286, // @[:@130706.4]
  input  [63:0] io_ins_287, // @[:@130706.4]
  input  [63:0] io_ins_288, // @[:@130706.4]
  input  [63:0] io_ins_289, // @[:@130706.4]
  input  [63:0] io_ins_290, // @[:@130706.4]
  input  [63:0] io_ins_291, // @[:@130706.4]
  input  [63:0] io_ins_292, // @[:@130706.4]
  input  [63:0] io_ins_293, // @[:@130706.4]
  input  [63:0] io_ins_294, // @[:@130706.4]
  input  [63:0] io_ins_295, // @[:@130706.4]
  input  [63:0] io_ins_296, // @[:@130706.4]
  input  [63:0] io_ins_297, // @[:@130706.4]
  input  [63:0] io_ins_298, // @[:@130706.4]
  input  [63:0] io_ins_299, // @[:@130706.4]
  input  [63:0] io_ins_300, // @[:@130706.4]
  input  [63:0] io_ins_301, // @[:@130706.4]
  input  [63:0] io_ins_302, // @[:@130706.4]
  input  [63:0] io_ins_303, // @[:@130706.4]
  input  [63:0] io_ins_304, // @[:@130706.4]
  input  [63:0] io_ins_305, // @[:@130706.4]
  input  [63:0] io_ins_306, // @[:@130706.4]
  input  [63:0] io_ins_307, // @[:@130706.4]
  input  [63:0] io_ins_308, // @[:@130706.4]
  input  [63:0] io_ins_309, // @[:@130706.4]
  input  [63:0] io_ins_310, // @[:@130706.4]
  input  [63:0] io_ins_311, // @[:@130706.4]
  input  [63:0] io_ins_312, // @[:@130706.4]
  input  [63:0] io_ins_313, // @[:@130706.4]
  input  [63:0] io_ins_314, // @[:@130706.4]
  input  [63:0] io_ins_315, // @[:@130706.4]
  input  [63:0] io_ins_316, // @[:@130706.4]
  input  [63:0] io_ins_317, // @[:@130706.4]
  input  [63:0] io_ins_318, // @[:@130706.4]
  input  [63:0] io_ins_319, // @[:@130706.4]
  input  [63:0] io_ins_320, // @[:@130706.4]
  input  [63:0] io_ins_321, // @[:@130706.4]
  input  [63:0] io_ins_322, // @[:@130706.4]
  input  [63:0] io_ins_323, // @[:@130706.4]
  input  [63:0] io_ins_324, // @[:@130706.4]
  input  [63:0] io_ins_325, // @[:@130706.4]
  input  [63:0] io_ins_326, // @[:@130706.4]
  input  [63:0] io_ins_327, // @[:@130706.4]
  input  [63:0] io_ins_328, // @[:@130706.4]
  input  [63:0] io_ins_329, // @[:@130706.4]
  input  [63:0] io_ins_330, // @[:@130706.4]
  input  [63:0] io_ins_331, // @[:@130706.4]
  input  [63:0] io_ins_332, // @[:@130706.4]
  input  [63:0] io_ins_333, // @[:@130706.4]
  input  [63:0] io_ins_334, // @[:@130706.4]
  input  [63:0] io_ins_335, // @[:@130706.4]
  input  [63:0] io_ins_336, // @[:@130706.4]
  input  [63:0] io_ins_337, // @[:@130706.4]
  input  [63:0] io_ins_338, // @[:@130706.4]
  input  [63:0] io_ins_339, // @[:@130706.4]
  input  [63:0] io_ins_340, // @[:@130706.4]
  input  [63:0] io_ins_341, // @[:@130706.4]
  input  [63:0] io_ins_342, // @[:@130706.4]
  input  [63:0] io_ins_343, // @[:@130706.4]
  input  [63:0] io_ins_344, // @[:@130706.4]
  input  [63:0] io_ins_345, // @[:@130706.4]
  input  [63:0] io_ins_346, // @[:@130706.4]
  input  [63:0] io_ins_347, // @[:@130706.4]
  input  [63:0] io_ins_348, // @[:@130706.4]
  input  [63:0] io_ins_349, // @[:@130706.4]
  input  [63:0] io_ins_350, // @[:@130706.4]
  input  [63:0] io_ins_351, // @[:@130706.4]
  input  [63:0] io_ins_352, // @[:@130706.4]
  input  [63:0] io_ins_353, // @[:@130706.4]
  input  [63:0] io_ins_354, // @[:@130706.4]
  input  [63:0] io_ins_355, // @[:@130706.4]
  input  [63:0] io_ins_356, // @[:@130706.4]
  input  [63:0] io_ins_357, // @[:@130706.4]
  input  [63:0] io_ins_358, // @[:@130706.4]
  input  [63:0] io_ins_359, // @[:@130706.4]
  input  [63:0] io_ins_360, // @[:@130706.4]
  input  [63:0] io_ins_361, // @[:@130706.4]
  input  [63:0] io_ins_362, // @[:@130706.4]
  input  [63:0] io_ins_363, // @[:@130706.4]
  input  [63:0] io_ins_364, // @[:@130706.4]
  input  [63:0] io_ins_365, // @[:@130706.4]
  input  [63:0] io_ins_366, // @[:@130706.4]
  input  [63:0] io_ins_367, // @[:@130706.4]
  input  [63:0] io_ins_368, // @[:@130706.4]
  input  [63:0] io_ins_369, // @[:@130706.4]
  input  [63:0] io_ins_370, // @[:@130706.4]
  input  [63:0] io_ins_371, // @[:@130706.4]
  input  [63:0] io_ins_372, // @[:@130706.4]
  input  [63:0] io_ins_373, // @[:@130706.4]
  input  [63:0] io_ins_374, // @[:@130706.4]
  input  [63:0] io_ins_375, // @[:@130706.4]
  input  [63:0] io_ins_376, // @[:@130706.4]
  input  [63:0] io_ins_377, // @[:@130706.4]
  input  [63:0] io_ins_378, // @[:@130706.4]
  input  [63:0] io_ins_379, // @[:@130706.4]
  input  [63:0] io_ins_380, // @[:@130706.4]
  input  [63:0] io_ins_381, // @[:@130706.4]
  input  [63:0] io_ins_382, // @[:@130706.4]
  input  [63:0] io_ins_383, // @[:@130706.4]
  input  [63:0] io_ins_384, // @[:@130706.4]
  input  [63:0] io_ins_385, // @[:@130706.4]
  input  [63:0] io_ins_386, // @[:@130706.4]
  input  [63:0] io_ins_387, // @[:@130706.4]
  input  [63:0] io_ins_388, // @[:@130706.4]
  input  [63:0] io_ins_389, // @[:@130706.4]
  input  [63:0] io_ins_390, // @[:@130706.4]
  input  [63:0] io_ins_391, // @[:@130706.4]
  input  [63:0] io_ins_392, // @[:@130706.4]
  input  [63:0] io_ins_393, // @[:@130706.4]
  input  [63:0] io_ins_394, // @[:@130706.4]
  input  [63:0] io_ins_395, // @[:@130706.4]
  input  [63:0] io_ins_396, // @[:@130706.4]
  input  [63:0] io_ins_397, // @[:@130706.4]
  input  [63:0] io_ins_398, // @[:@130706.4]
  input  [63:0] io_ins_399, // @[:@130706.4]
  input  [63:0] io_ins_400, // @[:@130706.4]
  input  [63:0] io_ins_401, // @[:@130706.4]
  input  [63:0] io_ins_402, // @[:@130706.4]
  input  [63:0] io_ins_403, // @[:@130706.4]
  input  [63:0] io_ins_404, // @[:@130706.4]
  input  [63:0] io_ins_405, // @[:@130706.4]
  input  [63:0] io_ins_406, // @[:@130706.4]
  input  [63:0] io_ins_407, // @[:@130706.4]
  input  [63:0] io_ins_408, // @[:@130706.4]
  input  [63:0] io_ins_409, // @[:@130706.4]
  input  [63:0] io_ins_410, // @[:@130706.4]
  input  [63:0] io_ins_411, // @[:@130706.4]
  input  [63:0] io_ins_412, // @[:@130706.4]
  input  [63:0] io_ins_413, // @[:@130706.4]
  input  [63:0] io_ins_414, // @[:@130706.4]
  input  [63:0] io_ins_415, // @[:@130706.4]
  input  [63:0] io_ins_416, // @[:@130706.4]
  input  [63:0] io_ins_417, // @[:@130706.4]
  input  [63:0] io_ins_418, // @[:@130706.4]
  input  [63:0] io_ins_419, // @[:@130706.4]
  input  [63:0] io_ins_420, // @[:@130706.4]
  input  [63:0] io_ins_421, // @[:@130706.4]
  input  [63:0] io_ins_422, // @[:@130706.4]
  input  [63:0] io_ins_423, // @[:@130706.4]
  input  [63:0] io_ins_424, // @[:@130706.4]
  input  [63:0] io_ins_425, // @[:@130706.4]
  input  [63:0] io_ins_426, // @[:@130706.4]
  input  [63:0] io_ins_427, // @[:@130706.4]
  input  [63:0] io_ins_428, // @[:@130706.4]
  input  [63:0] io_ins_429, // @[:@130706.4]
  input  [63:0] io_ins_430, // @[:@130706.4]
  input  [63:0] io_ins_431, // @[:@130706.4]
  input  [63:0] io_ins_432, // @[:@130706.4]
  input  [63:0] io_ins_433, // @[:@130706.4]
  input  [63:0] io_ins_434, // @[:@130706.4]
  input  [63:0] io_ins_435, // @[:@130706.4]
  input  [63:0] io_ins_436, // @[:@130706.4]
  input  [63:0] io_ins_437, // @[:@130706.4]
  input  [63:0] io_ins_438, // @[:@130706.4]
  input  [63:0] io_ins_439, // @[:@130706.4]
  input  [63:0] io_ins_440, // @[:@130706.4]
  input  [63:0] io_ins_441, // @[:@130706.4]
  input  [63:0] io_ins_442, // @[:@130706.4]
  input  [63:0] io_ins_443, // @[:@130706.4]
  input  [63:0] io_ins_444, // @[:@130706.4]
  input  [63:0] io_ins_445, // @[:@130706.4]
  input  [63:0] io_ins_446, // @[:@130706.4]
  input  [63:0] io_ins_447, // @[:@130706.4]
  input  [63:0] io_ins_448, // @[:@130706.4]
  input  [63:0] io_ins_449, // @[:@130706.4]
  input  [63:0] io_ins_450, // @[:@130706.4]
  input  [63:0] io_ins_451, // @[:@130706.4]
  input  [63:0] io_ins_452, // @[:@130706.4]
  input  [63:0] io_ins_453, // @[:@130706.4]
  input  [63:0] io_ins_454, // @[:@130706.4]
  input  [63:0] io_ins_455, // @[:@130706.4]
  input  [63:0] io_ins_456, // @[:@130706.4]
  input  [63:0] io_ins_457, // @[:@130706.4]
  input  [63:0] io_ins_458, // @[:@130706.4]
  input  [63:0] io_ins_459, // @[:@130706.4]
  input  [63:0] io_ins_460, // @[:@130706.4]
  input  [63:0] io_ins_461, // @[:@130706.4]
  input  [63:0] io_ins_462, // @[:@130706.4]
  input  [63:0] io_ins_463, // @[:@130706.4]
  input  [63:0] io_ins_464, // @[:@130706.4]
  input  [63:0] io_ins_465, // @[:@130706.4]
  input  [63:0] io_ins_466, // @[:@130706.4]
  input  [63:0] io_ins_467, // @[:@130706.4]
  input  [63:0] io_ins_468, // @[:@130706.4]
  input  [63:0] io_ins_469, // @[:@130706.4]
  input  [63:0] io_ins_470, // @[:@130706.4]
  input  [63:0] io_ins_471, // @[:@130706.4]
  input  [63:0] io_ins_472, // @[:@130706.4]
  input  [63:0] io_ins_473, // @[:@130706.4]
  input  [63:0] io_ins_474, // @[:@130706.4]
  input  [63:0] io_ins_475, // @[:@130706.4]
  input  [63:0] io_ins_476, // @[:@130706.4]
  input  [63:0] io_ins_477, // @[:@130706.4]
  input  [63:0] io_ins_478, // @[:@130706.4]
  input  [63:0] io_ins_479, // @[:@130706.4]
  input  [63:0] io_ins_480, // @[:@130706.4]
  input  [63:0] io_ins_481, // @[:@130706.4]
  input  [63:0] io_ins_482, // @[:@130706.4]
  input  [63:0] io_ins_483, // @[:@130706.4]
  input  [63:0] io_ins_484, // @[:@130706.4]
  input  [63:0] io_ins_485, // @[:@130706.4]
  input  [63:0] io_ins_486, // @[:@130706.4]
  input  [63:0] io_ins_487, // @[:@130706.4]
  input  [63:0] io_ins_488, // @[:@130706.4]
  input  [63:0] io_ins_489, // @[:@130706.4]
  input  [63:0] io_ins_490, // @[:@130706.4]
  input  [63:0] io_ins_491, // @[:@130706.4]
  input  [63:0] io_ins_492, // @[:@130706.4]
  input  [63:0] io_ins_493, // @[:@130706.4]
  input  [63:0] io_ins_494, // @[:@130706.4]
  input  [63:0] io_ins_495, // @[:@130706.4]
  input  [63:0] io_ins_496, // @[:@130706.4]
  input  [63:0] io_ins_497, // @[:@130706.4]
  input  [63:0] io_ins_498, // @[:@130706.4]
  input  [63:0] io_ins_499, // @[:@130706.4]
  input  [63:0] io_ins_500, // @[:@130706.4]
  input  [63:0] io_ins_501, // @[:@130706.4]
  input  [63:0] io_ins_502, // @[:@130706.4]
  input  [8:0]  io_sel, // @[:@130706.4]
  output [63:0] io_out // @[:@130706.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@130708.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@130708.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@130708.4]
  assign io_out = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@130708.4]
endmodule
module RegFile( // @[:@130710.2]
  input         clock, // @[:@130711.4]
  input         reset, // @[:@130712.4]
  input  [31:0] io_raddr, // @[:@130713.4]
  input         io_wen, // @[:@130713.4]
  input  [31:0] io_waddr, // @[:@130713.4]
  input  [63:0] io_wdata, // @[:@130713.4]
  output [63:0] io_rdata, // @[:@130713.4]
  input         io_reset, // @[:@130713.4]
  output [63:0] io_argIns_0, // @[:@130713.4]
  output [63:0] io_argIns_1, // @[:@130713.4]
  output [63:0] io_argIns_2, // @[:@130713.4]
  output [63:0] io_argIns_3, // @[:@130713.4]
  input         io_argOuts_0_valid, // @[:@130713.4]
  input  [63:0] io_argOuts_0_bits, // @[:@130713.4]
  input         io_argOuts_1_valid, // @[:@130713.4]
  input  [63:0] io_argOuts_1_bits // @[:@130713.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@132723.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@132723.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@132723.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@132723.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@132723.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@132723.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@132735.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@132735.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@132735.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@132735.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@132735.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@132735.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@132754.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@132754.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@132754.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@132754.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@132754.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@132754.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@132766.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@132766.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@132766.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@132766.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@132766.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@132766.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@132778.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@132778.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@132778.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@132778.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@132778.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@132778.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@132792.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@132792.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@132792.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@132792.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@132792.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@132792.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@132806.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@132806.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@132806.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@132806.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@132806.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@132806.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@132820.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@132820.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@132820.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@132820.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@132820.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@132820.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@132834.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@132834.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@132834.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@132834.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@132834.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@132834.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@132848.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@132848.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@132848.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@132848.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@132848.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@132848.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@132862.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@132862.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@132862.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@132862.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@132862.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@132862.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@132876.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@132876.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@132876.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@132876.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@132876.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@132876.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@132890.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@132890.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@132890.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@132890.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@132890.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@132890.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@132904.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@132904.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@132904.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@132904.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@132904.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@132904.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@132918.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@132918.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@132918.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@132918.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@132918.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@132918.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@132932.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@132932.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@132932.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@132932.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@132932.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@132932.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@132946.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@132946.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@132946.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@132946.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@132946.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@132946.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@132960.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@132960.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@132960.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@132960.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@132960.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@132960.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@132974.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@132974.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@132974.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@132974.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@132974.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@132974.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@132988.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@132988.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@132988.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@132988.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@132988.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@132988.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@133002.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@133002.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@133002.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@133002.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@133002.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@133002.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@133016.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@133016.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@133016.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@133016.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@133016.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@133016.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@133030.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@133030.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@133030.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@133030.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@133030.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@133030.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@133044.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@133044.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@133044.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@133044.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@133044.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@133044.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@133058.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@133058.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@133058.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@133058.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@133058.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@133058.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@133072.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@133072.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@133072.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@133072.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@133072.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@133072.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@133086.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@133086.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@133086.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@133086.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@133086.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@133086.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@133100.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@133100.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@133100.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@133100.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@133100.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@133100.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@133114.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@133114.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@133114.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@133114.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@133114.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@133114.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@133128.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@133128.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@133128.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@133128.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@133128.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@133128.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@133142.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@133142.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@133142.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@133142.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@133142.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@133142.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@133156.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@133156.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@133156.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@133156.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@133156.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@133156.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@133170.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@133170.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@133170.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@133170.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@133170.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@133170.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@133184.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@133184.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@133184.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@133184.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@133184.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@133184.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@133198.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@133198.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@133198.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@133198.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@133198.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@133198.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@133212.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@133212.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@133212.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@133212.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@133212.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@133212.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@133226.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@133226.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@133226.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@133226.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@133226.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@133226.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@133240.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@133240.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@133240.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@133240.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@133240.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@133240.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@133254.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@133254.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@133254.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@133254.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@133254.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@133254.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@133268.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@133268.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@133268.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@133268.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@133268.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@133268.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@133282.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@133282.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@133282.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@133282.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@133282.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@133282.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@133296.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@133296.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@133296.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@133296.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@133296.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@133296.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@133310.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@133310.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@133310.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@133310.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@133310.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@133310.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@133324.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@133324.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@133324.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@133324.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@133324.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@133324.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@133338.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@133338.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@133338.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@133338.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@133338.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@133338.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@133352.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@133352.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@133352.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@133352.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@133352.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@133352.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@133366.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@133366.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@133366.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@133366.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@133366.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@133366.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@133380.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@133380.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@133380.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@133380.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@133380.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@133380.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@133394.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@133394.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@133394.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@133394.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@133394.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@133394.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@133408.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@133408.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@133408.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@133408.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@133408.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@133408.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@133422.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@133422.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@133422.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@133422.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@133422.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@133422.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@133436.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@133436.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@133436.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@133436.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@133436.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@133436.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@133450.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@133450.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@133450.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@133450.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@133450.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@133450.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@133464.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@133464.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@133464.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@133464.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@133464.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@133464.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@133478.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@133478.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@133478.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@133478.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@133478.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@133478.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@133492.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@133492.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@133492.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@133492.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@133492.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@133492.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@133506.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@133506.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@133506.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@133506.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@133506.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@133506.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@133520.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@133520.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@133520.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@133520.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@133520.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@133520.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@133534.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@133534.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@133534.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@133534.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@133534.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@133534.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@133548.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@133548.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@133548.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@133548.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@133548.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@133548.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@133562.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@133562.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@133562.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@133562.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@133562.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@133562.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@133576.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@133576.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@133576.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@133576.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@133576.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@133576.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@133590.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@133590.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@133590.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@133590.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@133590.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@133590.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@133604.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@133604.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@133604.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@133604.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@133604.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@133604.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@133618.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@133618.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@133618.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@133618.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@133618.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@133618.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@133632.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@133632.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@133632.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@133632.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@133632.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@133632.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@133646.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@133646.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@133646.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@133646.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@133646.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@133646.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@133660.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@133660.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@133660.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@133660.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@133660.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@133660.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@133674.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@133674.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@133674.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@133674.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@133674.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@133674.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@133688.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@133688.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@133688.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@133688.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@133688.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@133688.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@133702.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@133702.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@133702.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@133702.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@133702.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@133702.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@133716.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@133716.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@133716.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@133716.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@133716.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@133716.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@133730.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@133730.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@133730.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@133730.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@133730.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@133730.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@133744.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@133744.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@133744.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@133744.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@133744.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@133744.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@133758.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@133758.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@133758.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@133758.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@133758.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@133758.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@133772.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@133772.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@133772.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@133772.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@133772.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@133772.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@133786.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@133786.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@133786.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@133786.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@133786.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@133786.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@133800.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@133800.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@133800.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@133800.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@133800.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@133800.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@133814.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@133814.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@133814.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@133814.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@133814.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@133814.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@133828.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@133828.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@133828.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@133828.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@133828.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@133828.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@133842.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@133842.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@133842.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@133842.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@133842.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@133842.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@133856.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@133856.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@133856.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@133856.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@133856.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@133856.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@133870.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@133870.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@133870.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@133870.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@133870.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@133870.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@133884.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@133884.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@133884.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@133884.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@133884.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@133884.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@133898.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@133898.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@133898.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@133898.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@133898.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@133898.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@133912.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@133912.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@133912.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@133912.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@133912.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@133912.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@133926.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@133926.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@133926.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@133926.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@133926.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@133926.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@133940.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@133940.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@133940.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@133940.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@133940.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@133940.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@133954.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@133954.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@133954.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@133954.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@133954.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@133954.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@133968.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@133968.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@133968.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@133968.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@133968.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@133968.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@133982.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@133982.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@133982.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@133982.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@133982.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@133982.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@133996.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@133996.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@133996.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@133996.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@133996.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@133996.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@134010.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@134010.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@134010.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@134010.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@134010.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@134010.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@134024.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@134024.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@134024.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@134024.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@134024.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@134024.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@134038.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@134038.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@134038.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@134038.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@134038.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@134038.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@134052.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@134052.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@134052.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@134052.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@134052.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@134052.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@134066.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@134066.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@134066.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@134066.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@134066.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@134066.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@134080.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@134080.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@134080.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@134080.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@134080.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@134080.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@134094.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@134094.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@134094.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@134094.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@134094.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@134094.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@134108.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@134108.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@134108.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@134108.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@134108.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@134108.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@134122.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@134122.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@134122.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@134122.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@134122.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@134122.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@134136.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@134136.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@134136.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@134136.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@134136.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@134136.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@134150.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@134150.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@134150.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@134150.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@134150.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@134150.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@134164.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@134164.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@134164.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@134164.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@134164.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@134164.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@134178.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@134178.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@134178.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@134178.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@134178.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@134178.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@134192.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@134192.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@134192.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@134192.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@134192.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@134192.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@134206.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@134206.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@134206.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@134206.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@134206.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@134206.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@134220.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@134220.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@134220.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@134220.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@134220.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@134220.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@134234.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@134234.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@134234.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@134234.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@134234.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@134234.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@134248.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@134248.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@134248.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@134248.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@134248.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@134248.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@134262.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@134262.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@134262.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@134262.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@134262.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@134262.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@134276.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@134276.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@134276.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@134276.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@134276.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@134276.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@134290.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@134290.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@134290.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@134290.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@134290.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@134290.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@134304.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@134304.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@134304.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@134304.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@134304.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@134304.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@134318.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@134318.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@134318.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@134318.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@134318.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@134318.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@134332.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@134332.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@134332.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@134332.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@134332.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@134332.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@134346.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@134346.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@134346.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@134346.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@134346.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@134346.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@134360.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@134360.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@134360.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@134360.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@134360.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@134360.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@134374.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@134374.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@134374.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@134374.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@134374.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@134374.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@134388.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@134388.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@134388.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@134388.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@134388.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@134388.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@134402.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@134402.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@134402.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@134402.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@134402.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@134402.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@134416.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@134416.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@134416.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@134416.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@134416.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@134416.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@134430.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@134430.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@134430.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@134430.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@134430.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@134430.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@134444.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@134444.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@134444.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@134444.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@134444.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@134444.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@134458.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@134458.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@134458.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@134458.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@134458.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@134458.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@134472.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@134472.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@134472.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@134472.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@134472.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@134472.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@134486.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@134486.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@134486.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@134486.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@134486.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@134486.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@134500.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@134500.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@134500.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@134500.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@134500.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@134500.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@134514.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@134514.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@134514.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@134514.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@134514.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@134514.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@134528.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@134528.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@134528.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@134528.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@134528.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@134528.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@134542.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@134542.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@134542.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@134542.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@134542.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@134542.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@134556.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@134556.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@134556.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@134556.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@134556.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@134556.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@134570.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@134570.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@134570.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@134570.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@134570.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@134570.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@134584.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@134584.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@134584.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@134584.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@134584.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@134584.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@134598.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@134598.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@134598.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@134598.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@134598.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@134598.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@134612.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@134612.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@134612.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@134612.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@134612.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@134612.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@134626.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@134626.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@134626.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@134626.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@134626.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@134626.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@134640.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@134640.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@134640.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@134640.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@134640.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@134640.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@134654.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@134654.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@134654.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@134654.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@134654.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@134654.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@134668.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@134668.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@134668.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@134668.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@134668.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@134668.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@134682.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@134682.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@134682.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@134682.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@134682.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@134682.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@134696.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@134696.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@134696.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@134696.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@134696.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@134696.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@134710.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@134710.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@134710.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@134710.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@134710.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@134710.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@134724.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@134724.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@134724.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@134724.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@134724.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@134724.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@134738.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@134738.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@134738.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@134738.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@134738.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@134738.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@134752.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@134752.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@134752.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@134752.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@134752.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@134752.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@134766.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@134766.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@134766.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@134766.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@134766.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@134766.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@134780.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@134780.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@134780.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@134780.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@134780.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@134780.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@134794.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@134794.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@134794.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@134794.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@134794.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@134794.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@134808.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@134808.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@134808.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@134808.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@134808.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@134808.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@134822.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@134822.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@134822.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@134822.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@134822.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@134822.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@134836.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@134836.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@134836.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@134836.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@134836.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@134836.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@134850.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@134850.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@134850.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@134850.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@134850.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@134850.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@134864.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@134864.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@134864.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@134864.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@134864.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@134864.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@134878.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@134878.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@134878.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@134878.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@134878.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@134878.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@134892.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@134892.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@134892.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@134892.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@134892.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@134892.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@134906.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@134906.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@134906.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@134906.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@134906.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@134906.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@134920.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@134920.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@134920.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@134920.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@134920.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@134920.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@134934.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@134934.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@134934.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@134934.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@134934.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@134934.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@134948.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@134948.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@134948.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@134948.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@134948.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@134948.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@134962.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@134962.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@134962.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@134962.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@134962.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@134962.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@134976.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@134976.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@134976.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@134976.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@134976.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@134976.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@134990.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@134990.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@134990.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@134990.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@134990.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@134990.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@135004.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@135004.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@135004.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@135004.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@135004.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@135004.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@135018.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@135018.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@135018.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@135018.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@135018.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@135018.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@135032.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@135032.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@135032.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@135032.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@135032.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@135032.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@135046.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@135046.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@135046.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@135046.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@135046.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@135046.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@135060.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@135060.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@135060.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@135060.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@135060.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@135060.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@135074.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@135074.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@135074.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@135074.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@135074.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@135074.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@135088.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@135088.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@135088.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@135088.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@135088.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@135088.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@135102.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@135102.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@135102.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@135102.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@135102.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@135102.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@135116.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@135116.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@135116.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@135116.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@135116.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@135116.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@135130.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@135130.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@135130.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@135130.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@135130.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@135130.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@135144.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@135144.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@135144.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@135144.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@135144.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@135144.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@135158.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@135158.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@135158.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@135158.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@135158.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@135158.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@135172.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@135172.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@135172.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@135172.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@135172.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@135172.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@135186.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@135186.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@135186.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@135186.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@135186.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@135186.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@135200.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@135200.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@135200.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@135200.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@135200.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@135200.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@135214.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@135214.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@135214.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@135214.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@135214.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@135214.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@135228.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@135228.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@135228.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@135228.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@135228.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@135228.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@135242.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@135242.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@135242.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@135242.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@135242.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@135242.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@135256.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@135256.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@135256.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@135256.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@135256.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@135256.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@135270.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@135270.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@135270.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@135270.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@135270.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@135270.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@135284.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@135284.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@135284.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@135284.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@135284.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@135284.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@135298.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@135298.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@135298.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@135298.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@135298.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@135298.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@135312.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@135312.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@135312.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@135312.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@135312.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@135312.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@135326.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@135326.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@135326.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@135326.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@135326.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@135326.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@135340.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@135340.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@135340.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@135340.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@135340.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@135340.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@135354.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@135354.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@135354.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@135354.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@135354.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@135354.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@135368.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@135368.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@135368.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@135368.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@135368.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@135368.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@135382.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@135382.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@135382.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@135382.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@135382.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@135382.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@135396.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@135396.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@135396.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@135396.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@135396.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@135396.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@135410.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@135410.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@135410.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@135410.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@135410.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@135410.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@135424.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@135424.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@135424.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@135424.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@135424.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@135424.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@135438.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@135438.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@135438.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@135438.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@135438.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@135438.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@135452.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@135452.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@135452.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@135452.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@135452.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@135452.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@135466.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@135466.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@135466.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@135466.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@135466.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@135466.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@135480.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@135480.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@135480.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@135480.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@135480.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@135480.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@135494.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@135494.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@135494.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@135494.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@135494.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@135494.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@135508.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@135508.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@135508.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@135508.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@135508.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@135508.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@135522.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@135522.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@135522.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@135522.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@135522.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@135522.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@135536.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@135536.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@135536.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@135536.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@135536.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@135536.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@135550.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@135550.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@135550.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@135550.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@135550.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@135550.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@135564.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@135564.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@135564.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@135564.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@135564.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@135564.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@135578.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@135578.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@135578.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@135578.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@135578.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@135578.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@135592.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@135592.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@135592.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@135592.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@135592.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@135592.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@135606.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@135606.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@135606.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@135606.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@135606.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@135606.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@135620.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@135620.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@135620.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@135620.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@135620.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@135620.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@135634.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@135634.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@135634.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@135634.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@135634.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@135634.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@135648.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@135648.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@135648.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@135648.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@135648.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@135648.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@135662.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@135662.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@135662.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@135662.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@135662.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@135662.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@135676.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@135676.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@135676.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@135676.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@135676.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@135676.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@135690.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@135690.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@135690.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@135690.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@135690.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@135690.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@135704.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@135704.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@135704.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@135704.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@135704.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@135704.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@135718.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@135718.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@135718.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@135718.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@135718.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@135718.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@135732.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@135732.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@135732.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@135732.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@135732.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@135732.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@135746.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@135746.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@135746.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@135746.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@135746.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@135746.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@135760.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@135760.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@135760.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@135760.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@135760.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@135760.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@135774.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@135774.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@135774.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@135774.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@135774.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@135774.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@135788.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@135788.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@135788.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@135788.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@135788.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@135788.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@135802.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@135802.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@135802.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@135802.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@135802.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@135802.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@135816.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@135816.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@135816.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@135816.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@135816.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@135816.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@135830.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@135830.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@135830.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@135830.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@135830.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@135830.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@135844.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@135844.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@135844.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@135844.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@135844.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@135844.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@135858.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@135858.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@135858.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@135858.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@135858.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@135858.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@135872.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@135872.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@135872.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@135872.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@135872.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@135872.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@135886.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@135886.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@135886.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@135886.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@135886.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@135886.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@135900.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@135900.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@135900.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@135900.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@135900.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@135900.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@135914.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@135914.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@135914.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@135914.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@135914.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@135914.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@135928.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@135928.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@135928.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@135928.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@135928.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@135928.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@135942.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@135942.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@135942.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@135942.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@135942.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@135942.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@135956.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@135956.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@135956.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@135956.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@135956.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@135956.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@135970.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@135970.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@135970.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@135970.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@135970.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@135970.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@135984.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@135984.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@135984.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@135984.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@135984.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@135984.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@135998.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@135998.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@135998.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@135998.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@135998.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@135998.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@136012.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@136012.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@136012.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@136012.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@136012.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@136012.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@136026.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@136026.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@136026.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@136026.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@136026.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@136026.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@136040.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@136040.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@136040.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@136040.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@136040.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@136040.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@136054.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@136054.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@136054.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@136054.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@136054.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@136054.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@136068.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@136068.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@136068.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@136068.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@136068.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@136068.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@136082.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@136082.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@136082.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@136082.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@136082.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@136082.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@136096.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@136096.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@136096.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@136096.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@136096.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@136096.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@136110.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@136110.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@136110.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@136110.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@136110.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@136110.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@136124.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@136124.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@136124.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@136124.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@136124.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@136124.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@136138.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@136138.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@136138.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@136138.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@136138.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@136138.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@136152.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@136152.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@136152.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@136152.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@136152.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@136152.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@136166.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@136166.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@136166.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@136166.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@136166.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@136166.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@136180.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@136180.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@136180.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@136180.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@136180.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@136180.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@136194.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@136194.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@136194.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@136194.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@136194.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@136194.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@136208.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@136208.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@136208.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@136208.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@136208.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@136208.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@136222.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@136222.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@136222.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@136222.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@136222.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@136222.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@136236.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@136236.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@136236.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@136236.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@136236.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@136236.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@136250.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@136250.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@136250.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@136250.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@136250.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@136250.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@136264.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@136264.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@136264.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@136264.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@136264.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@136264.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@136278.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@136278.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@136278.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@136278.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@136278.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@136278.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@136292.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@136292.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@136292.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@136292.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@136292.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@136292.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@136306.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@136306.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@136306.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@136306.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@136306.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@136306.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@136320.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@136320.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@136320.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@136320.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@136320.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@136320.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@136334.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@136334.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@136334.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@136334.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@136334.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@136334.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@136348.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@136348.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@136348.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@136348.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@136348.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@136348.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@136362.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@136362.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@136362.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@136362.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@136362.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@136362.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@136376.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@136376.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@136376.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@136376.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@136376.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@136376.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@136390.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@136390.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@136390.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@136390.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@136390.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@136390.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@136404.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@136404.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@136404.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@136404.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@136404.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@136404.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@136418.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@136418.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@136418.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@136418.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@136418.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@136418.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@136432.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@136432.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@136432.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@136432.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@136432.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@136432.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@136446.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@136446.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@136446.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@136446.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@136446.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@136446.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@136460.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@136460.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@136460.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@136460.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@136460.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@136460.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@136474.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@136474.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@136474.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@136474.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@136474.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@136474.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@136488.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@136488.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@136488.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@136488.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@136488.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@136488.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@136502.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@136502.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@136502.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@136502.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@136502.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@136502.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@136516.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@136516.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@136516.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@136516.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@136516.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@136516.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@136530.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@136530.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@136530.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@136530.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@136530.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@136530.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@136544.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@136544.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@136544.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@136544.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@136544.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@136544.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@136558.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@136558.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@136558.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@136558.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@136558.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@136558.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@136572.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@136572.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@136572.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@136572.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@136572.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@136572.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@136586.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@136586.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@136586.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@136586.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@136586.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@136586.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@136600.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@136600.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@136600.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@136600.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@136600.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@136600.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@136614.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@136614.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@136614.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@136614.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@136614.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@136614.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@136628.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@136628.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@136628.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@136628.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@136628.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@136628.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@136642.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@136642.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@136642.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@136642.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@136642.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@136642.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@136656.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@136656.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@136656.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@136656.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@136656.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@136656.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@136670.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@136670.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@136670.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@136670.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@136670.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@136670.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@136684.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@136684.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@136684.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@136684.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@136684.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@136684.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@136698.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@136698.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@136698.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@136698.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@136698.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@136698.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@136712.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@136712.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@136712.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@136712.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@136712.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@136712.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@136726.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@136726.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@136726.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@136726.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@136726.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@136726.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@136740.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@136740.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@136740.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@136740.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@136740.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@136740.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@136754.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@136754.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@136754.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@136754.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@136754.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@136754.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@136768.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@136768.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@136768.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@136768.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@136768.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@136768.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@136782.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@136782.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@136782.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@136782.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@136782.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@136782.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@136796.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@136796.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@136796.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@136796.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@136796.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@136796.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@136810.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@136810.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@136810.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@136810.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@136810.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@136810.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@136824.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@136824.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@136824.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@136824.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@136824.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@136824.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@136838.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@136838.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@136838.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@136838.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@136838.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@136838.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@136852.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@136852.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@136852.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@136852.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@136852.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@136852.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@136866.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@136866.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@136866.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@136866.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@136866.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@136866.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@136880.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@136880.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@136880.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@136880.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@136880.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@136880.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@136894.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@136894.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@136894.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@136894.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@136894.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@136894.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@136908.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@136908.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@136908.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@136908.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@136908.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@136908.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@136922.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@136922.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@136922.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@136922.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@136922.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@136922.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@136936.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@136936.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@136936.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@136936.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@136936.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@136936.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@136950.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@136950.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@136950.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@136950.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@136950.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@136950.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@136964.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@136964.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@136964.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@136964.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@136964.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@136964.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@136978.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@136978.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@136978.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@136978.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@136978.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@136978.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@136992.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@136992.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@136992.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@136992.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@136992.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@136992.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@137006.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@137006.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@137006.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@137006.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@137006.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@137006.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@137020.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@137020.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@137020.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@137020.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@137020.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@137020.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@137034.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@137034.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@137034.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@137034.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@137034.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@137034.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@137048.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@137048.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@137048.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@137048.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@137048.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@137048.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@137062.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@137062.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@137062.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@137062.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@137062.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@137062.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@137076.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@137076.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@137076.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@137076.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@137076.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@137076.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@137090.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@137090.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@137090.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@137090.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@137090.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@137090.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@137104.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@137104.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@137104.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@137104.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@137104.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@137104.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@137118.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@137118.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@137118.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@137118.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@137118.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@137118.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@137132.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@137132.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@137132.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@137132.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@137132.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@137132.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@137146.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@137146.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@137146.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@137146.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@137146.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@137146.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@137160.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@137160.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@137160.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@137160.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@137160.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@137160.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@137174.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@137174.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@137174.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@137174.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@137174.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@137174.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@137188.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@137188.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@137188.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@137188.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@137188.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@137188.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@137202.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@137202.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@137202.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@137202.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@137202.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@137202.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@137216.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@137216.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@137216.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@137216.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@137216.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@137216.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@137230.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@137230.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@137230.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@137230.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@137230.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@137230.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@137244.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@137244.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@137244.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@137244.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@137244.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@137244.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@137258.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@137258.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@137258.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@137258.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@137258.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@137258.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@137272.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@137272.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@137272.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@137272.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@137272.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@137272.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@137286.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@137286.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@137286.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@137286.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@137286.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@137286.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@137300.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@137300.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@137300.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@137300.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@137300.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@137300.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@137314.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@137314.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@137314.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@137314.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@137314.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@137314.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@137328.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@137328.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@137328.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@137328.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@137328.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@137328.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@137342.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@137342.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@137342.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@137342.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@137342.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@137342.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@137356.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@137356.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@137356.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@137356.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@137356.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@137356.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@137370.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@137370.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@137370.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@137370.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@137370.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@137370.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@137384.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@137384.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@137384.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@137384.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@137384.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@137384.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@137398.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@137398.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@137398.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@137398.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@137398.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@137398.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@137412.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@137412.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@137412.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@137412.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@137412.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@137412.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@137426.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@137426.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@137426.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@137426.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@137426.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@137426.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@137440.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@137440.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@137440.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@137440.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@137440.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@137440.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@137454.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@137454.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@137454.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@137454.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@137454.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@137454.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@137468.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@137468.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@137468.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@137468.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@137468.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@137468.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@137482.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@137482.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@137482.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@137482.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@137482.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@137482.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@137496.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@137496.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@137496.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@137496.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@137496.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@137496.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@137510.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@137510.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@137510.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@137510.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@137510.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@137510.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@137524.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@137524.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@137524.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@137524.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@137524.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@137524.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@137538.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@137538.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@137538.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@137538.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@137538.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@137538.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@137552.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@137552.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@137552.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@137552.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@137552.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@137552.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@137566.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@137566.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@137566.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@137566.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@137566.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@137566.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@137580.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@137580.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@137580.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@137580.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@137580.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@137580.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@137594.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@137594.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@137594.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@137594.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@137594.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@137594.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@137608.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@137608.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@137608.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@137608.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@137608.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@137608.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@137622.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@137622.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@137622.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@137622.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@137622.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@137622.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@137636.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@137636.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@137636.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@137636.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@137636.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@137636.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@137650.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@137650.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@137650.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@137650.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@137650.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@137650.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@137664.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@137664.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@137664.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@137664.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@137664.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@137664.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@137678.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@137678.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@137678.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@137678.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@137678.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@137678.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@137692.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@137692.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@137692.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@137692.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@137692.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@137692.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@137706.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@137706.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@137706.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@137706.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@137706.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@137706.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@137720.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@137720.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@137720.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@137720.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@137720.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@137720.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@137734.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@137734.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@137734.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@137734.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@137734.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@137734.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@137748.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@137748.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@137748.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@137748.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@137748.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@137748.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@137762.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@137762.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@137762.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@137762.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@137762.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@137762.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@137776.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@137776.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@137776.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@137776.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@137776.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@137776.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@137790.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@137790.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@137790.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@137790.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@137790.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@137790.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@137804.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@137804.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@137804.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@137804.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@137804.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@137804.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@137818.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@137818.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@137818.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@137818.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@137818.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@137818.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@137832.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@137832.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@137832.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@137832.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@137832.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@137832.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@137846.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@137846.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@137846.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@137846.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@137846.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@137846.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@137860.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@137860.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@137860.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@137860.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@137860.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@137860.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@137874.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@137874.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@137874.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@137874.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@137874.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@137874.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@137888.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@137888.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@137888.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@137888.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@137888.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@137888.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@137902.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@137902.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@137902.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@137902.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@137902.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@137902.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@137916.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@137916.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@137916.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@137916.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@137916.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@137916.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@137930.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@137930.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@137930.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@137930.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@137930.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@137930.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@137944.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@137944.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@137944.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@137944.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@137944.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@137944.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@137958.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@137958.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@137958.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@137958.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@137958.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@137958.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@137972.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@137972.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@137972.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@137972.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@137972.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@137972.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@137986.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@137986.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@137986.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@137986.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@137986.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@137986.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@138000.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@138000.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@138000.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@138000.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@138000.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@138000.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@138014.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@138014.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@138014.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@138014.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@138014.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@138014.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@138028.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@138028.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@138028.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@138028.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@138028.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@138028.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@138042.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@138042.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@138042.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@138042.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@138042.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@138042.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@138056.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@138056.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@138056.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@138056.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@138056.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@138056.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@138070.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@138070.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@138070.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@138070.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@138070.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@138070.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@138084.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@138084.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@138084.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@138084.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@138084.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@138084.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@138098.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@138098.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@138098.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@138098.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@138098.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@138098.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@138112.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@138112.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@138112.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@138112.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@138112.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@138112.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@138126.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@138126.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@138126.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@138126.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@138126.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@138126.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@138140.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@138140.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@138140.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@138140.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@138140.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@138140.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@138154.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@138154.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@138154.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@138154.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@138154.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@138154.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@138168.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@138168.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@138168.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@138168.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@138168.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@138168.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@138182.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@138182.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@138182.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@138182.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@138182.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@138182.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@138196.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@138196.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@138196.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@138196.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@138196.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@138196.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@138210.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@138210.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@138210.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@138210.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@138210.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@138210.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@138224.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@138224.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@138224.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@138224.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@138224.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@138224.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@138238.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@138238.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@138238.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@138238.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@138238.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@138238.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@138252.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@138252.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@138252.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@138252.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@138252.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@138252.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@138266.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@138266.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@138266.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@138266.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@138266.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@138266.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@138280.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@138280.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@138280.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@138280.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@138280.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@138280.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@138294.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@138294.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@138294.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@138294.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@138294.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@138294.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@138308.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@138308.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@138308.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@138308.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@138308.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@138308.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@138322.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@138322.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@138322.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@138322.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@138322.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@138322.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@138336.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@138336.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@138336.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@138336.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@138336.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@138336.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@138350.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@138350.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@138350.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@138350.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@138350.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@138350.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@138364.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@138364.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@138364.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@138364.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@138364.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@138364.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@138378.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@138378.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@138378.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@138378.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@138378.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@138378.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@138392.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@138392.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@138392.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@138392.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@138392.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@138392.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@138406.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@138406.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@138406.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@138406.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@138406.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@138406.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@138420.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@138420.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@138420.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@138420.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@138420.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@138420.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@138434.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@138434.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@138434.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@138434.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@138434.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@138434.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@138448.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@138448.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@138448.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@138448.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@138448.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@138448.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@138462.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@138462.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@138462.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@138462.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@138462.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@138462.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@138476.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@138476.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@138476.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@138476.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@138476.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@138476.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@138490.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@138490.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@138490.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@138490.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@138490.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@138490.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@138504.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@138504.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@138504.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@138504.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@138504.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@138504.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@138518.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@138518.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@138518.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@138518.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@138518.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@138518.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@138532.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@138532.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@138532.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@138532.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@138532.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@138532.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@138546.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@138546.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@138546.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@138546.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@138546.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@138546.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@138560.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@138560.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@138560.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@138560.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@138560.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@138560.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@138574.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@138574.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@138574.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@138574.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@138574.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@138574.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@138588.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@138588.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@138588.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@138588.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@138588.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@138588.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@138602.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@138602.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@138602.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@138602.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@138602.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@138602.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@138616.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@138616.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@138616.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@138616.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@138616.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@138616.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@138630.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@138630.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@138630.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@138630.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@138630.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@138630.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@138644.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@138644.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@138644.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@138644.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@138644.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@138644.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@138658.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@138658.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@138658.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@138658.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@138658.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@138658.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@138672.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@138672.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@138672.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@138672.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@138672.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@138672.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@138686.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@138686.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@138686.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@138686.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@138686.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@138686.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@138700.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@138700.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@138700.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@138700.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@138700.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@138700.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@138714.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@138714.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@138714.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@138714.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@138714.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@138714.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@138728.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@138728.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@138728.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@138728.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@138728.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@138728.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@138742.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@138742.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@138742.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@138742.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@138742.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@138742.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@138756.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@138756.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@138756.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@138756.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@138756.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@138756.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@138770.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@138770.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@138770.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@138770.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@138770.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@138770.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@138784.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@138784.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@138784.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@138784.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@138784.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@138784.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@138798.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@138798.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@138798.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@138798.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@138798.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@138798.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@138812.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@138812.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@138812.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@138812.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@138812.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@138812.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@138826.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@138826.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@138826.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@138826.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@138826.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@138826.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@138840.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@138840.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@138840.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@138840.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@138840.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@138840.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@138854.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@138854.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@138854.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@138854.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@138854.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@138854.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@138868.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@138868.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@138868.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@138868.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@138868.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@138868.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@138882.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@138882.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@138882.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@138882.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@138882.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@138882.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@138896.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@138896.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@138896.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@138896.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@138896.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@138896.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@138910.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@138910.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@138910.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@138910.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@138910.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@138910.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@138924.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@138924.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@138924.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@138924.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@138924.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@138924.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@138938.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@138938.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@138938.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@138938.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@138938.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@138938.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@138952.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@138952.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@138952.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@138952.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@138952.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@138952.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@138966.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@138966.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@138966.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@138966.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@138966.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@138966.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@138980.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@138980.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@138980.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@138980.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@138980.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@138980.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@138994.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@138994.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@138994.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@138994.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@138994.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@138994.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@139008.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@139008.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@139008.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@139008.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@139008.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@139008.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@139022.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@139022.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@139022.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@139022.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@139022.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@139022.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@139036.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@139036.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@139036.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@139036.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@139036.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@139036.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@139050.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@139050.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@139050.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@139050.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@139050.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@139050.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@139064.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@139064.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@139064.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@139064.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@139064.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@139064.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@139078.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@139078.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@139078.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@139078.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@139078.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@139078.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@139092.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@139092.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@139092.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@139092.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@139092.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@139092.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@139106.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@139106.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@139106.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@139106.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@139106.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@139106.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@139120.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@139120.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@139120.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@139120.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@139120.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@139120.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@139134.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@139134.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@139134.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@139134.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@139134.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@139134.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@139148.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@139148.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@139148.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@139148.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@139148.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@139148.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@139162.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@139162.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@139162.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@139162.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@139162.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@139162.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@139176.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@139176.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@139176.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@139176.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@139176.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@139176.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@139190.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@139190.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@139190.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@139190.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@139190.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@139190.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@139204.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@139204.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@139204.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@139204.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@139204.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@139204.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@139218.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@139218.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@139218.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@139218.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@139218.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@139218.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@139232.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@139232.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@139232.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@139232.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@139232.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@139232.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@139246.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@139246.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@139246.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@139246.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@139246.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@139246.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@139260.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@139260.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@139260.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@139260.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@139260.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@139260.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@139274.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@139274.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@139274.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@139274.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@139274.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@139274.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@139288.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@139288.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@139288.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@139288.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@139288.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@139288.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@139302.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@139302.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@139302.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@139302.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@139302.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@139302.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@139316.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@139316.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@139316.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@139316.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@139316.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@139316.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@139330.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@139330.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@139330.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@139330.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@139330.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@139330.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@139344.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@139344.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@139344.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@139344.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@139344.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@139344.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@139358.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@139358.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@139358.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@139358.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@139358.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@139358.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@139372.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@139372.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@139372.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@139372.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@139372.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@139372.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@139386.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@139386.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@139386.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@139386.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@139386.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@139386.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@139400.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@139400.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@139400.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@139400.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@139400.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@139400.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@139414.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@139414.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@139414.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@139414.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@139414.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@139414.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@139428.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@139428.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@139428.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@139428.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@139428.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@139428.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@139442.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@139442.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@139442.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@139442.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@139442.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@139442.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@139456.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@139456.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@139456.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@139456.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@139456.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@139456.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@139470.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@139470.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@139470.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@139470.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@139470.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@139470.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@139484.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@139484.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@139484.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@139484.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@139484.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@139484.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@139498.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@139498.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@139498.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@139498.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@139498.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@139498.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@139512.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@139512.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@139512.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@139512.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@139512.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@139512.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@139526.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@139526.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@139526.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@139526.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@139526.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@139526.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@139540.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@139540.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@139540.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@139540.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@139540.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@139540.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@139554.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@139554.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@139554.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@139554.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@139554.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@139554.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@139568.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@139568.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@139568.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@139568.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@139568.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@139568.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@139582.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@139582.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@139582.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@139582.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@139582.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@139582.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@139596.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@139596.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@139596.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@139596.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@139596.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@139596.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@139610.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@139610.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@139610.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@139610.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@139610.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@139610.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@139624.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@139624.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@139624.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@139624.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@139624.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@139624.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@139638.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@139638.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@139638.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@139638.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@139638.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@139638.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@139652.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@139652.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@139652.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@139652.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@139652.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@139652.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@139666.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@139666.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@139666.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@139666.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@139666.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@139666.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@139680.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@139680.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@139680.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@139680.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@139680.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@139680.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@139694.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@139694.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@139694.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@139694.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@139694.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@139694.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@139708.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@139708.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@139708.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@139708.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@139708.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@139708.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@139722.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@139722.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@139722.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@139722.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@139722.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@139722.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@139736.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@139736.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@139736.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@139736.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@139736.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@139736.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@139750.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@139750.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@139750.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@139750.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@139750.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@139750.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@139764.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@139764.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@139764.4]
  wire  _T_3078; // @[RegFile.scala 80:42:@132726.4]
  wire  _T_3084; // @[RegFile.scala 68:46:@132738.4]
  wire  _T_3085; // @[RegFile.scala 68:34:@132739.4]
  wire  _T_3098; // @[RegFile.scala 80:42:@132757.4]
  wire  _T_3104; // @[RegFile.scala 80:42:@132769.4]
  wire  _T_3110; // @[RegFile.scala 74:80:@132781.4]
  wire  _T_3111; // @[RegFile.scala 74:68:@132782.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@132723.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@132735.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@132754.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@132766.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@132778.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@132792.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@132806.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@132820.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@132834.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@132848.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@132862.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@132876.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@132890.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@132904.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@132918.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@132932.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@132946.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@132960.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@132974.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@132988.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@133002.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@133016.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@133030.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@133044.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@133058.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@133072.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@133086.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@133100.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@133114.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@133128.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@133142.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@133156.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@133170.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@133184.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@133198.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@133212.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@133226.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@133240.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@133254.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@133268.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@133282.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@133296.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@133310.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@133324.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@133338.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@133352.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@133366.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@133380.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@133394.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@133408.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@133422.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@133436.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@133450.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@133464.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@133478.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@133492.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@133506.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@133520.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@133534.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@133548.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@133562.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@133576.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@133590.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@133604.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@133618.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@133632.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@133646.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@133660.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@133674.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@133688.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@133702.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@133716.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@133730.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@133744.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@133758.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@133772.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@133786.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@133800.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@133814.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@133828.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@133842.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@133856.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@133870.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@133884.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@133898.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@133912.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@133926.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@133940.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@133954.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@133968.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@133982.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@133996.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@134010.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@134024.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@134038.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@134052.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@134066.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@134080.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@134094.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@134108.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@134122.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@134136.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@134150.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@134164.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@134178.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@134192.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@134206.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@134220.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@134234.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@134248.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@134262.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@134276.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@134290.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@134304.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@134318.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@134332.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@134346.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@134360.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@134374.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@134388.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@134402.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@134416.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@134430.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@134444.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@134458.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@134472.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@134486.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@134500.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@134514.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@134528.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@134542.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@134556.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@134570.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@134584.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@134598.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@134612.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@134626.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@134640.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@134654.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@134668.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@134682.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@134696.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@134710.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@134724.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@134738.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@134752.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@134766.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@134780.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@134794.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@134808.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@134822.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@134836.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@134850.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@134864.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@134878.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@134892.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@134906.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@134920.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@134934.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@134948.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@134962.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@134976.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@134990.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@135004.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@135018.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@135032.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@135046.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@135060.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@135074.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@135088.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@135102.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@135116.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@135130.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@135144.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@135158.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@135172.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@135186.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@135200.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@135214.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@135228.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@135242.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@135256.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@135270.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@135284.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@135298.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@135312.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@135326.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@135340.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@135354.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@135368.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@135382.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@135396.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@135410.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@135424.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@135438.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@135452.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@135466.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@135480.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@135494.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@135508.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@135522.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@135536.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@135550.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@135564.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@135578.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@135592.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@135606.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@135620.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@135634.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@135648.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@135662.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@135676.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@135690.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@135704.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@135718.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@135732.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@135746.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@135760.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@135774.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@135788.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@135802.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@135816.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@135830.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@135844.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@135858.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@135872.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@135886.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@135900.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@135914.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@135928.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@135942.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@135956.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@135970.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@135984.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@135998.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@136012.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@136026.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@136040.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@136054.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@136068.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@136082.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@136096.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@136110.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@136124.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@136138.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@136152.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@136166.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@136180.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@136194.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@136208.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@136222.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@136236.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@136250.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@136264.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@136278.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@136292.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@136306.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@136320.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@136334.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@136348.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@136362.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@136376.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@136390.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@136404.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@136418.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@136432.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@136446.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@136460.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@136474.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@136488.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@136502.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@136516.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@136530.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@136544.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@136558.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@136572.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@136586.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@136600.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@136614.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@136628.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@136642.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@136656.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@136670.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@136684.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@136698.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@136712.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@136726.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@136740.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@136754.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@136768.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@136782.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@136796.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@136810.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@136824.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@136838.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@136852.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@136866.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@136880.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@136894.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@136908.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@136922.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@136936.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@136950.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@136964.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@136978.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@136992.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@137006.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@137020.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@137034.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@137048.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@137062.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@137076.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@137090.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@137104.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@137118.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@137132.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@137146.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@137160.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@137174.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@137188.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@137202.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@137216.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@137230.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@137244.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@137258.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@137272.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@137286.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@137300.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@137314.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@137328.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@137342.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@137356.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@137370.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@137384.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@137398.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@137412.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@137426.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@137440.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@137454.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@137468.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@137482.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@137496.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@137510.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@137524.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@137538.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@137552.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@137566.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@137580.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@137594.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@137608.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@137622.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@137636.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@137650.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@137664.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@137678.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@137692.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@137706.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@137720.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@137734.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@137748.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@137762.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@137776.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@137790.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@137804.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@137818.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@137832.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@137846.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@137860.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@137874.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@137888.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@137902.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@137916.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@137930.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@137944.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@137958.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@137972.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@137986.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@138000.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@138014.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@138028.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@138042.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@138056.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@138070.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@138084.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@138098.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@138112.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@138126.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@138140.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@138154.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@138168.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@138182.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@138196.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@138210.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@138224.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@138238.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@138252.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@138266.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@138280.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@138294.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@138308.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@138322.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@138336.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@138350.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@138364.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@138378.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@138392.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@138406.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@138420.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@138434.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@138448.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@138462.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@138476.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@138490.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@138504.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@138518.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@138532.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@138546.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@138560.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@138574.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@138588.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@138602.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@138616.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@138630.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@138644.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@138658.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@138672.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@138686.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@138700.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@138714.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@138728.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@138742.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@138756.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@138770.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@138784.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@138798.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@138812.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@138826.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@138840.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@138854.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@138868.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@138882.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@138896.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@138910.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@138924.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@138938.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@138952.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@138966.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@138980.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@138994.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@139008.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@139022.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@139036.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@139050.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@139064.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@139078.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@139092.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@139106.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@139120.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@139134.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@139148.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@139162.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@139176.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@139190.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@139204.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@139218.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@139232.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@139246.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@139260.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@139274.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@139288.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@139302.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@139316.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@139330.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@139344.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@139358.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@139372.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@139386.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@139400.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@139414.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@139428.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@139442.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@139456.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@139470.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@139484.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@139498.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@139512.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@139526.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@139540.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@139554.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@139568.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@139582.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@139596.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@139610.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@139624.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@139638.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@139652.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@139666.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@139680.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@139694.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@139708.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@139722.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@139736.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@139750.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@139764.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3078 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@132726.4]
  assign _T_3084 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@132738.4]
  assign _T_3085 = io_wen & _T_3084; // @[RegFile.scala 68:34:@132739.4]
  assign _T_3098 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@132757.4]
  assign _T_3104 = io_waddr == 32'h3; // @[RegFile.scala 80:42:@132769.4]
  assign _T_3110 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@132781.4]
  assign _T_3111 = io_wen & _T_3110; // @[RegFile.scala 74:68:@132782.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@140775.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@140781.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@140782.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@140783.4]
  assign io_argIns_3 = regs_3_io_out; // @[RegFile.scala 111:13:@140784.4]
  assign regs_0_clock = clock; // @[:@132724.4]
  assign regs_0_reset = reset; // @[:@132725.4 RegFile.scala 82:16:@132731.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@132729.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@132733.4]
  assign regs_0_io_enable = io_wen & _T_3078; // @[RegFile.scala 80:20:@132728.4]
  assign regs_1_clock = clock; // @[:@132736.4]
  assign regs_1_reset = reset; // @[:@132737.4 RegFile.scala 70:16:@132749.4]
  assign regs_1_io_in = _T_3085 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@132747.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@132752.4]
  assign regs_1_io_enable = _T_3085 ? _T_3085 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@132743.4]
  assign regs_2_clock = clock; // @[:@132755.4]
  assign regs_2_reset = reset; // @[:@132756.4 RegFile.scala 82:16:@132762.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@132760.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@132764.4]
  assign regs_2_io_enable = io_wen & _T_3098; // @[RegFile.scala 80:20:@132759.4]
  assign regs_3_clock = clock; // @[:@132767.4]
  assign regs_3_reset = reset; // @[:@132768.4 RegFile.scala 82:16:@132774.4]
  assign regs_3_io_in = io_wdata; // @[RegFile.scala 81:16:@132772.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 83:19:@132776.4]
  assign regs_3_io_enable = io_wen & _T_3104; // @[RegFile.scala 80:20:@132771.4]
  assign regs_4_clock = clock; // @[:@132779.4]
  assign regs_4_reset = io_reset; // @[:@132780.4 RegFile.scala 76:16:@132787.4]
  assign regs_4_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@132786.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@132790.4]
  assign regs_4_io_enable = io_argOuts_1_valid | _T_3111; // @[RegFile.scala 74:20:@132784.4]
  assign regs_5_clock = clock; // @[:@132793.4]
  assign regs_5_reset = io_reset; // @[:@132794.4 RegFile.scala 76:16:@132801.4]
  assign regs_5_io_in = 64'h0; // @[RegFile.scala 75:16:@132800.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@132804.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 74:20:@132798.4]
  assign regs_6_clock = clock; // @[:@132807.4]
  assign regs_6_reset = io_reset; // @[:@132808.4 RegFile.scala 76:16:@132815.4]
  assign regs_6_io_in = 64'h0; // @[RegFile.scala 75:16:@132814.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@132818.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 74:20:@132812.4]
  assign regs_7_clock = clock; // @[:@132821.4]
  assign regs_7_reset = io_reset; // @[:@132822.4 RegFile.scala 76:16:@132829.4]
  assign regs_7_io_in = 64'h0; // @[RegFile.scala 75:16:@132828.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@132832.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 74:20:@132826.4]
  assign regs_8_clock = clock; // @[:@132835.4]
  assign regs_8_reset = io_reset; // @[:@132836.4 RegFile.scala 76:16:@132843.4]
  assign regs_8_io_in = 64'h0; // @[RegFile.scala 75:16:@132842.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@132846.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 74:20:@132840.4]
  assign regs_9_clock = clock; // @[:@132849.4]
  assign regs_9_reset = io_reset; // @[:@132850.4 RegFile.scala 76:16:@132857.4]
  assign regs_9_io_in = 64'h0; // @[RegFile.scala 75:16:@132856.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@132860.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 74:20:@132854.4]
  assign regs_10_clock = clock; // @[:@132863.4]
  assign regs_10_reset = io_reset; // @[:@132864.4 RegFile.scala 76:16:@132871.4]
  assign regs_10_io_in = 64'h0; // @[RegFile.scala 75:16:@132870.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@132874.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 74:20:@132868.4]
  assign regs_11_clock = clock; // @[:@132877.4]
  assign regs_11_reset = io_reset; // @[:@132878.4 RegFile.scala 76:16:@132885.4]
  assign regs_11_io_in = 64'h0; // @[RegFile.scala 75:16:@132884.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@132888.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 74:20:@132882.4]
  assign regs_12_clock = clock; // @[:@132891.4]
  assign regs_12_reset = io_reset; // @[:@132892.4 RegFile.scala 76:16:@132899.4]
  assign regs_12_io_in = 64'h0; // @[RegFile.scala 75:16:@132898.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@132902.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 74:20:@132896.4]
  assign regs_13_clock = clock; // @[:@132905.4]
  assign regs_13_reset = io_reset; // @[:@132906.4 RegFile.scala 76:16:@132913.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 75:16:@132912.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@132916.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@132910.4]
  assign regs_14_clock = clock; // @[:@132919.4]
  assign regs_14_reset = io_reset; // @[:@132920.4 RegFile.scala 76:16:@132927.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 75:16:@132926.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@132930.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@132924.4]
  assign regs_15_clock = clock; // @[:@132933.4]
  assign regs_15_reset = io_reset; // @[:@132934.4 RegFile.scala 76:16:@132941.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 75:16:@132940.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@132944.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@132938.4]
  assign regs_16_clock = clock; // @[:@132947.4]
  assign regs_16_reset = io_reset; // @[:@132948.4 RegFile.scala 76:16:@132955.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 75:16:@132954.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@132958.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@132952.4]
  assign regs_17_clock = clock; // @[:@132961.4]
  assign regs_17_reset = io_reset; // @[:@132962.4 RegFile.scala 76:16:@132969.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 75:16:@132968.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@132972.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@132966.4]
  assign regs_18_clock = clock; // @[:@132975.4]
  assign regs_18_reset = io_reset; // @[:@132976.4 RegFile.scala 76:16:@132983.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 75:16:@132982.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@132986.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@132980.4]
  assign regs_19_clock = clock; // @[:@132989.4]
  assign regs_19_reset = io_reset; // @[:@132990.4 RegFile.scala 76:16:@132997.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 75:16:@132996.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@133000.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@132994.4]
  assign regs_20_clock = clock; // @[:@133003.4]
  assign regs_20_reset = io_reset; // @[:@133004.4 RegFile.scala 76:16:@133011.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 75:16:@133010.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@133014.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@133008.4]
  assign regs_21_clock = clock; // @[:@133017.4]
  assign regs_21_reset = io_reset; // @[:@133018.4 RegFile.scala 76:16:@133025.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 75:16:@133024.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@133028.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@133022.4]
  assign regs_22_clock = clock; // @[:@133031.4]
  assign regs_22_reset = io_reset; // @[:@133032.4 RegFile.scala 76:16:@133039.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 75:16:@133038.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@133042.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@133036.4]
  assign regs_23_clock = clock; // @[:@133045.4]
  assign regs_23_reset = io_reset; // @[:@133046.4 RegFile.scala 76:16:@133053.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@133052.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@133056.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@133050.4]
  assign regs_24_clock = clock; // @[:@133059.4]
  assign regs_24_reset = io_reset; // @[:@133060.4 RegFile.scala 76:16:@133067.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@133066.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@133070.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@133064.4]
  assign regs_25_clock = clock; // @[:@133073.4]
  assign regs_25_reset = io_reset; // @[:@133074.4 RegFile.scala 76:16:@133081.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@133080.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@133084.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@133078.4]
  assign regs_26_clock = clock; // @[:@133087.4]
  assign regs_26_reset = io_reset; // @[:@133088.4 RegFile.scala 76:16:@133095.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@133094.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@133098.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@133092.4]
  assign regs_27_clock = clock; // @[:@133101.4]
  assign regs_27_reset = io_reset; // @[:@133102.4 RegFile.scala 76:16:@133109.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@133108.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@133112.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@133106.4]
  assign regs_28_clock = clock; // @[:@133115.4]
  assign regs_28_reset = io_reset; // @[:@133116.4 RegFile.scala 76:16:@133123.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@133122.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@133126.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@133120.4]
  assign regs_29_clock = clock; // @[:@133129.4]
  assign regs_29_reset = io_reset; // @[:@133130.4 RegFile.scala 76:16:@133137.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@133136.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@133140.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@133134.4]
  assign regs_30_clock = clock; // @[:@133143.4]
  assign regs_30_reset = io_reset; // @[:@133144.4 RegFile.scala 76:16:@133151.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@133150.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@133154.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@133148.4]
  assign regs_31_clock = clock; // @[:@133157.4]
  assign regs_31_reset = io_reset; // @[:@133158.4 RegFile.scala 76:16:@133165.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@133164.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@133168.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@133162.4]
  assign regs_32_clock = clock; // @[:@133171.4]
  assign regs_32_reset = io_reset; // @[:@133172.4 RegFile.scala 76:16:@133179.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@133178.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@133182.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@133176.4]
  assign regs_33_clock = clock; // @[:@133185.4]
  assign regs_33_reset = io_reset; // @[:@133186.4 RegFile.scala 76:16:@133193.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@133192.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@133196.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@133190.4]
  assign regs_34_clock = clock; // @[:@133199.4]
  assign regs_34_reset = io_reset; // @[:@133200.4 RegFile.scala 76:16:@133207.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@133206.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@133210.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@133204.4]
  assign regs_35_clock = clock; // @[:@133213.4]
  assign regs_35_reset = io_reset; // @[:@133214.4 RegFile.scala 76:16:@133221.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@133220.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@133224.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@133218.4]
  assign regs_36_clock = clock; // @[:@133227.4]
  assign regs_36_reset = io_reset; // @[:@133228.4 RegFile.scala 76:16:@133235.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@133234.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@133238.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@133232.4]
  assign regs_37_clock = clock; // @[:@133241.4]
  assign regs_37_reset = io_reset; // @[:@133242.4 RegFile.scala 76:16:@133249.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@133248.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@133252.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@133246.4]
  assign regs_38_clock = clock; // @[:@133255.4]
  assign regs_38_reset = io_reset; // @[:@133256.4 RegFile.scala 76:16:@133263.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@133262.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@133266.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@133260.4]
  assign regs_39_clock = clock; // @[:@133269.4]
  assign regs_39_reset = io_reset; // @[:@133270.4 RegFile.scala 76:16:@133277.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@133276.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@133280.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@133274.4]
  assign regs_40_clock = clock; // @[:@133283.4]
  assign regs_40_reset = io_reset; // @[:@133284.4 RegFile.scala 76:16:@133291.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@133290.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@133294.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@133288.4]
  assign regs_41_clock = clock; // @[:@133297.4]
  assign regs_41_reset = io_reset; // @[:@133298.4 RegFile.scala 76:16:@133305.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@133304.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@133308.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@133302.4]
  assign regs_42_clock = clock; // @[:@133311.4]
  assign regs_42_reset = io_reset; // @[:@133312.4 RegFile.scala 76:16:@133319.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@133318.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@133322.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@133316.4]
  assign regs_43_clock = clock; // @[:@133325.4]
  assign regs_43_reset = io_reset; // @[:@133326.4 RegFile.scala 76:16:@133333.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@133332.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@133336.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@133330.4]
  assign regs_44_clock = clock; // @[:@133339.4]
  assign regs_44_reset = io_reset; // @[:@133340.4 RegFile.scala 76:16:@133347.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@133346.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@133350.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@133344.4]
  assign regs_45_clock = clock; // @[:@133353.4]
  assign regs_45_reset = io_reset; // @[:@133354.4 RegFile.scala 76:16:@133361.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@133360.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@133364.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@133358.4]
  assign regs_46_clock = clock; // @[:@133367.4]
  assign regs_46_reset = io_reset; // @[:@133368.4 RegFile.scala 76:16:@133375.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@133374.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@133378.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@133372.4]
  assign regs_47_clock = clock; // @[:@133381.4]
  assign regs_47_reset = io_reset; // @[:@133382.4 RegFile.scala 76:16:@133389.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@133388.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@133392.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@133386.4]
  assign regs_48_clock = clock; // @[:@133395.4]
  assign regs_48_reset = io_reset; // @[:@133396.4 RegFile.scala 76:16:@133403.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@133402.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@133406.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@133400.4]
  assign regs_49_clock = clock; // @[:@133409.4]
  assign regs_49_reset = io_reset; // @[:@133410.4 RegFile.scala 76:16:@133417.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@133416.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@133420.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@133414.4]
  assign regs_50_clock = clock; // @[:@133423.4]
  assign regs_50_reset = io_reset; // @[:@133424.4 RegFile.scala 76:16:@133431.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@133430.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@133434.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@133428.4]
  assign regs_51_clock = clock; // @[:@133437.4]
  assign regs_51_reset = io_reset; // @[:@133438.4 RegFile.scala 76:16:@133445.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@133444.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@133448.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@133442.4]
  assign regs_52_clock = clock; // @[:@133451.4]
  assign regs_52_reset = io_reset; // @[:@133452.4 RegFile.scala 76:16:@133459.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@133458.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@133462.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@133456.4]
  assign regs_53_clock = clock; // @[:@133465.4]
  assign regs_53_reset = io_reset; // @[:@133466.4 RegFile.scala 76:16:@133473.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@133472.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@133476.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@133470.4]
  assign regs_54_clock = clock; // @[:@133479.4]
  assign regs_54_reset = io_reset; // @[:@133480.4 RegFile.scala 76:16:@133487.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@133486.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@133490.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@133484.4]
  assign regs_55_clock = clock; // @[:@133493.4]
  assign regs_55_reset = io_reset; // @[:@133494.4 RegFile.scala 76:16:@133501.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@133500.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@133504.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@133498.4]
  assign regs_56_clock = clock; // @[:@133507.4]
  assign regs_56_reset = io_reset; // @[:@133508.4 RegFile.scala 76:16:@133515.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@133514.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@133518.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@133512.4]
  assign regs_57_clock = clock; // @[:@133521.4]
  assign regs_57_reset = io_reset; // @[:@133522.4 RegFile.scala 76:16:@133529.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@133528.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@133532.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@133526.4]
  assign regs_58_clock = clock; // @[:@133535.4]
  assign regs_58_reset = io_reset; // @[:@133536.4 RegFile.scala 76:16:@133543.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@133542.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@133546.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@133540.4]
  assign regs_59_clock = clock; // @[:@133549.4]
  assign regs_59_reset = io_reset; // @[:@133550.4 RegFile.scala 76:16:@133557.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@133556.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@133560.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@133554.4]
  assign regs_60_clock = clock; // @[:@133563.4]
  assign regs_60_reset = io_reset; // @[:@133564.4 RegFile.scala 76:16:@133571.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@133570.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@133574.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@133568.4]
  assign regs_61_clock = clock; // @[:@133577.4]
  assign regs_61_reset = io_reset; // @[:@133578.4 RegFile.scala 76:16:@133585.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@133584.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@133588.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@133582.4]
  assign regs_62_clock = clock; // @[:@133591.4]
  assign regs_62_reset = io_reset; // @[:@133592.4 RegFile.scala 76:16:@133599.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@133598.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@133602.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@133596.4]
  assign regs_63_clock = clock; // @[:@133605.4]
  assign regs_63_reset = io_reset; // @[:@133606.4 RegFile.scala 76:16:@133613.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@133612.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@133616.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@133610.4]
  assign regs_64_clock = clock; // @[:@133619.4]
  assign regs_64_reset = io_reset; // @[:@133620.4 RegFile.scala 76:16:@133627.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@133626.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@133630.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@133624.4]
  assign regs_65_clock = clock; // @[:@133633.4]
  assign regs_65_reset = io_reset; // @[:@133634.4 RegFile.scala 76:16:@133641.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@133640.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@133644.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@133638.4]
  assign regs_66_clock = clock; // @[:@133647.4]
  assign regs_66_reset = io_reset; // @[:@133648.4 RegFile.scala 76:16:@133655.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@133654.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@133658.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@133652.4]
  assign regs_67_clock = clock; // @[:@133661.4]
  assign regs_67_reset = io_reset; // @[:@133662.4 RegFile.scala 76:16:@133669.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@133668.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@133672.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@133666.4]
  assign regs_68_clock = clock; // @[:@133675.4]
  assign regs_68_reset = io_reset; // @[:@133676.4 RegFile.scala 76:16:@133683.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@133682.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@133686.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@133680.4]
  assign regs_69_clock = clock; // @[:@133689.4]
  assign regs_69_reset = io_reset; // @[:@133690.4 RegFile.scala 76:16:@133697.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@133696.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@133700.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@133694.4]
  assign regs_70_clock = clock; // @[:@133703.4]
  assign regs_70_reset = io_reset; // @[:@133704.4 RegFile.scala 76:16:@133711.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@133710.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@133714.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@133708.4]
  assign regs_71_clock = clock; // @[:@133717.4]
  assign regs_71_reset = io_reset; // @[:@133718.4 RegFile.scala 76:16:@133725.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@133724.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@133728.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@133722.4]
  assign regs_72_clock = clock; // @[:@133731.4]
  assign regs_72_reset = io_reset; // @[:@133732.4 RegFile.scala 76:16:@133739.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@133738.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@133742.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@133736.4]
  assign regs_73_clock = clock; // @[:@133745.4]
  assign regs_73_reset = io_reset; // @[:@133746.4 RegFile.scala 76:16:@133753.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@133752.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@133756.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@133750.4]
  assign regs_74_clock = clock; // @[:@133759.4]
  assign regs_74_reset = io_reset; // @[:@133760.4 RegFile.scala 76:16:@133767.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@133766.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@133770.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@133764.4]
  assign regs_75_clock = clock; // @[:@133773.4]
  assign regs_75_reset = io_reset; // @[:@133774.4 RegFile.scala 76:16:@133781.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@133780.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@133784.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@133778.4]
  assign regs_76_clock = clock; // @[:@133787.4]
  assign regs_76_reset = io_reset; // @[:@133788.4 RegFile.scala 76:16:@133795.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@133794.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@133798.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@133792.4]
  assign regs_77_clock = clock; // @[:@133801.4]
  assign regs_77_reset = io_reset; // @[:@133802.4 RegFile.scala 76:16:@133809.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@133808.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@133812.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@133806.4]
  assign regs_78_clock = clock; // @[:@133815.4]
  assign regs_78_reset = io_reset; // @[:@133816.4 RegFile.scala 76:16:@133823.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@133822.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@133826.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@133820.4]
  assign regs_79_clock = clock; // @[:@133829.4]
  assign regs_79_reset = io_reset; // @[:@133830.4 RegFile.scala 76:16:@133837.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@133836.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@133840.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@133834.4]
  assign regs_80_clock = clock; // @[:@133843.4]
  assign regs_80_reset = io_reset; // @[:@133844.4 RegFile.scala 76:16:@133851.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@133850.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@133854.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@133848.4]
  assign regs_81_clock = clock; // @[:@133857.4]
  assign regs_81_reset = io_reset; // @[:@133858.4 RegFile.scala 76:16:@133865.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@133864.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@133868.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@133862.4]
  assign regs_82_clock = clock; // @[:@133871.4]
  assign regs_82_reset = io_reset; // @[:@133872.4 RegFile.scala 76:16:@133879.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@133878.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@133882.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@133876.4]
  assign regs_83_clock = clock; // @[:@133885.4]
  assign regs_83_reset = io_reset; // @[:@133886.4 RegFile.scala 76:16:@133893.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@133892.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@133896.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@133890.4]
  assign regs_84_clock = clock; // @[:@133899.4]
  assign regs_84_reset = io_reset; // @[:@133900.4 RegFile.scala 76:16:@133907.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@133906.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@133910.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@133904.4]
  assign regs_85_clock = clock; // @[:@133913.4]
  assign regs_85_reset = io_reset; // @[:@133914.4 RegFile.scala 76:16:@133921.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@133920.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@133924.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@133918.4]
  assign regs_86_clock = clock; // @[:@133927.4]
  assign regs_86_reset = io_reset; // @[:@133928.4 RegFile.scala 76:16:@133935.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@133934.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@133938.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@133932.4]
  assign regs_87_clock = clock; // @[:@133941.4]
  assign regs_87_reset = io_reset; // @[:@133942.4 RegFile.scala 76:16:@133949.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@133948.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@133952.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@133946.4]
  assign regs_88_clock = clock; // @[:@133955.4]
  assign regs_88_reset = io_reset; // @[:@133956.4 RegFile.scala 76:16:@133963.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@133962.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@133966.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@133960.4]
  assign regs_89_clock = clock; // @[:@133969.4]
  assign regs_89_reset = io_reset; // @[:@133970.4 RegFile.scala 76:16:@133977.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@133976.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@133980.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@133974.4]
  assign regs_90_clock = clock; // @[:@133983.4]
  assign regs_90_reset = io_reset; // @[:@133984.4 RegFile.scala 76:16:@133991.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@133990.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@133994.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@133988.4]
  assign regs_91_clock = clock; // @[:@133997.4]
  assign regs_91_reset = io_reset; // @[:@133998.4 RegFile.scala 76:16:@134005.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@134004.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@134008.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@134002.4]
  assign regs_92_clock = clock; // @[:@134011.4]
  assign regs_92_reset = io_reset; // @[:@134012.4 RegFile.scala 76:16:@134019.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@134018.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@134022.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@134016.4]
  assign regs_93_clock = clock; // @[:@134025.4]
  assign regs_93_reset = io_reset; // @[:@134026.4 RegFile.scala 76:16:@134033.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@134032.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@134036.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@134030.4]
  assign regs_94_clock = clock; // @[:@134039.4]
  assign regs_94_reset = io_reset; // @[:@134040.4 RegFile.scala 76:16:@134047.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@134046.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@134050.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@134044.4]
  assign regs_95_clock = clock; // @[:@134053.4]
  assign regs_95_reset = io_reset; // @[:@134054.4 RegFile.scala 76:16:@134061.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@134060.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@134064.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@134058.4]
  assign regs_96_clock = clock; // @[:@134067.4]
  assign regs_96_reset = io_reset; // @[:@134068.4 RegFile.scala 76:16:@134075.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@134074.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@134078.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@134072.4]
  assign regs_97_clock = clock; // @[:@134081.4]
  assign regs_97_reset = io_reset; // @[:@134082.4 RegFile.scala 76:16:@134089.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@134088.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@134092.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@134086.4]
  assign regs_98_clock = clock; // @[:@134095.4]
  assign regs_98_reset = io_reset; // @[:@134096.4 RegFile.scala 76:16:@134103.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@134102.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@134106.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@134100.4]
  assign regs_99_clock = clock; // @[:@134109.4]
  assign regs_99_reset = io_reset; // @[:@134110.4 RegFile.scala 76:16:@134117.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@134116.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@134120.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@134114.4]
  assign regs_100_clock = clock; // @[:@134123.4]
  assign regs_100_reset = io_reset; // @[:@134124.4 RegFile.scala 76:16:@134131.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@134130.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@134134.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@134128.4]
  assign regs_101_clock = clock; // @[:@134137.4]
  assign regs_101_reset = io_reset; // @[:@134138.4 RegFile.scala 76:16:@134145.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@134144.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@134148.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@134142.4]
  assign regs_102_clock = clock; // @[:@134151.4]
  assign regs_102_reset = io_reset; // @[:@134152.4 RegFile.scala 76:16:@134159.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@134158.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@134162.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@134156.4]
  assign regs_103_clock = clock; // @[:@134165.4]
  assign regs_103_reset = io_reset; // @[:@134166.4 RegFile.scala 76:16:@134173.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@134172.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@134176.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@134170.4]
  assign regs_104_clock = clock; // @[:@134179.4]
  assign regs_104_reset = io_reset; // @[:@134180.4 RegFile.scala 76:16:@134187.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@134186.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@134190.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@134184.4]
  assign regs_105_clock = clock; // @[:@134193.4]
  assign regs_105_reset = io_reset; // @[:@134194.4 RegFile.scala 76:16:@134201.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@134200.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@134204.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@134198.4]
  assign regs_106_clock = clock; // @[:@134207.4]
  assign regs_106_reset = io_reset; // @[:@134208.4 RegFile.scala 76:16:@134215.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@134214.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@134218.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@134212.4]
  assign regs_107_clock = clock; // @[:@134221.4]
  assign regs_107_reset = io_reset; // @[:@134222.4 RegFile.scala 76:16:@134229.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@134228.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@134232.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@134226.4]
  assign regs_108_clock = clock; // @[:@134235.4]
  assign regs_108_reset = io_reset; // @[:@134236.4 RegFile.scala 76:16:@134243.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@134242.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@134246.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@134240.4]
  assign regs_109_clock = clock; // @[:@134249.4]
  assign regs_109_reset = io_reset; // @[:@134250.4 RegFile.scala 76:16:@134257.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@134256.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@134260.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@134254.4]
  assign regs_110_clock = clock; // @[:@134263.4]
  assign regs_110_reset = io_reset; // @[:@134264.4 RegFile.scala 76:16:@134271.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@134270.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@134274.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@134268.4]
  assign regs_111_clock = clock; // @[:@134277.4]
  assign regs_111_reset = io_reset; // @[:@134278.4 RegFile.scala 76:16:@134285.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@134284.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@134288.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@134282.4]
  assign regs_112_clock = clock; // @[:@134291.4]
  assign regs_112_reset = io_reset; // @[:@134292.4 RegFile.scala 76:16:@134299.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@134298.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@134302.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@134296.4]
  assign regs_113_clock = clock; // @[:@134305.4]
  assign regs_113_reset = io_reset; // @[:@134306.4 RegFile.scala 76:16:@134313.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@134312.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@134316.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@134310.4]
  assign regs_114_clock = clock; // @[:@134319.4]
  assign regs_114_reset = io_reset; // @[:@134320.4 RegFile.scala 76:16:@134327.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@134326.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@134330.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@134324.4]
  assign regs_115_clock = clock; // @[:@134333.4]
  assign regs_115_reset = io_reset; // @[:@134334.4 RegFile.scala 76:16:@134341.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@134340.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@134344.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@134338.4]
  assign regs_116_clock = clock; // @[:@134347.4]
  assign regs_116_reset = io_reset; // @[:@134348.4 RegFile.scala 76:16:@134355.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@134354.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@134358.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@134352.4]
  assign regs_117_clock = clock; // @[:@134361.4]
  assign regs_117_reset = io_reset; // @[:@134362.4 RegFile.scala 76:16:@134369.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@134368.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@134372.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@134366.4]
  assign regs_118_clock = clock; // @[:@134375.4]
  assign regs_118_reset = io_reset; // @[:@134376.4 RegFile.scala 76:16:@134383.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@134382.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@134386.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@134380.4]
  assign regs_119_clock = clock; // @[:@134389.4]
  assign regs_119_reset = io_reset; // @[:@134390.4 RegFile.scala 76:16:@134397.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@134396.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@134400.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@134394.4]
  assign regs_120_clock = clock; // @[:@134403.4]
  assign regs_120_reset = io_reset; // @[:@134404.4 RegFile.scala 76:16:@134411.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@134410.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@134414.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@134408.4]
  assign regs_121_clock = clock; // @[:@134417.4]
  assign regs_121_reset = io_reset; // @[:@134418.4 RegFile.scala 76:16:@134425.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@134424.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@134428.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@134422.4]
  assign regs_122_clock = clock; // @[:@134431.4]
  assign regs_122_reset = io_reset; // @[:@134432.4 RegFile.scala 76:16:@134439.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@134438.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@134442.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@134436.4]
  assign regs_123_clock = clock; // @[:@134445.4]
  assign regs_123_reset = io_reset; // @[:@134446.4 RegFile.scala 76:16:@134453.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@134452.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@134456.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@134450.4]
  assign regs_124_clock = clock; // @[:@134459.4]
  assign regs_124_reset = io_reset; // @[:@134460.4 RegFile.scala 76:16:@134467.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@134466.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@134470.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@134464.4]
  assign regs_125_clock = clock; // @[:@134473.4]
  assign regs_125_reset = io_reset; // @[:@134474.4 RegFile.scala 76:16:@134481.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@134480.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@134484.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@134478.4]
  assign regs_126_clock = clock; // @[:@134487.4]
  assign regs_126_reset = io_reset; // @[:@134488.4 RegFile.scala 76:16:@134495.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@134494.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@134498.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@134492.4]
  assign regs_127_clock = clock; // @[:@134501.4]
  assign regs_127_reset = io_reset; // @[:@134502.4 RegFile.scala 76:16:@134509.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@134508.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@134512.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@134506.4]
  assign regs_128_clock = clock; // @[:@134515.4]
  assign regs_128_reset = io_reset; // @[:@134516.4 RegFile.scala 76:16:@134523.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@134522.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@134526.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@134520.4]
  assign regs_129_clock = clock; // @[:@134529.4]
  assign regs_129_reset = io_reset; // @[:@134530.4 RegFile.scala 76:16:@134537.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@134536.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@134540.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@134534.4]
  assign regs_130_clock = clock; // @[:@134543.4]
  assign regs_130_reset = io_reset; // @[:@134544.4 RegFile.scala 76:16:@134551.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@134550.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@134554.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@134548.4]
  assign regs_131_clock = clock; // @[:@134557.4]
  assign regs_131_reset = io_reset; // @[:@134558.4 RegFile.scala 76:16:@134565.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@134564.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@134568.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@134562.4]
  assign regs_132_clock = clock; // @[:@134571.4]
  assign regs_132_reset = io_reset; // @[:@134572.4 RegFile.scala 76:16:@134579.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@134578.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@134582.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@134576.4]
  assign regs_133_clock = clock; // @[:@134585.4]
  assign regs_133_reset = io_reset; // @[:@134586.4 RegFile.scala 76:16:@134593.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@134592.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@134596.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@134590.4]
  assign regs_134_clock = clock; // @[:@134599.4]
  assign regs_134_reset = io_reset; // @[:@134600.4 RegFile.scala 76:16:@134607.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@134606.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@134610.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@134604.4]
  assign regs_135_clock = clock; // @[:@134613.4]
  assign regs_135_reset = io_reset; // @[:@134614.4 RegFile.scala 76:16:@134621.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@134620.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@134624.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@134618.4]
  assign regs_136_clock = clock; // @[:@134627.4]
  assign regs_136_reset = io_reset; // @[:@134628.4 RegFile.scala 76:16:@134635.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@134634.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@134638.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@134632.4]
  assign regs_137_clock = clock; // @[:@134641.4]
  assign regs_137_reset = io_reset; // @[:@134642.4 RegFile.scala 76:16:@134649.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@134648.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@134652.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@134646.4]
  assign regs_138_clock = clock; // @[:@134655.4]
  assign regs_138_reset = io_reset; // @[:@134656.4 RegFile.scala 76:16:@134663.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@134662.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@134666.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@134660.4]
  assign regs_139_clock = clock; // @[:@134669.4]
  assign regs_139_reset = io_reset; // @[:@134670.4 RegFile.scala 76:16:@134677.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@134676.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@134680.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@134674.4]
  assign regs_140_clock = clock; // @[:@134683.4]
  assign regs_140_reset = io_reset; // @[:@134684.4 RegFile.scala 76:16:@134691.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@134690.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@134694.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@134688.4]
  assign regs_141_clock = clock; // @[:@134697.4]
  assign regs_141_reset = io_reset; // @[:@134698.4 RegFile.scala 76:16:@134705.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@134704.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@134708.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@134702.4]
  assign regs_142_clock = clock; // @[:@134711.4]
  assign regs_142_reset = io_reset; // @[:@134712.4 RegFile.scala 76:16:@134719.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@134718.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@134722.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@134716.4]
  assign regs_143_clock = clock; // @[:@134725.4]
  assign regs_143_reset = io_reset; // @[:@134726.4 RegFile.scala 76:16:@134733.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@134732.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@134736.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@134730.4]
  assign regs_144_clock = clock; // @[:@134739.4]
  assign regs_144_reset = io_reset; // @[:@134740.4 RegFile.scala 76:16:@134747.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@134746.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@134750.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@134744.4]
  assign regs_145_clock = clock; // @[:@134753.4]
  assign regs_145_reset = io_reset; // @[:@134754.4 RegFile.scala 76:16:@134761.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@134760.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@134764.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@134758.4]
  assign regs_146_clock = clock; // @[:@134767.4]
  assign regs_146_reset = io_reset; // @[:@134768.4 RegFile.scala 76:16:@134775.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@134774.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@134778.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@134772.4]
  assign regs_147_clock = clock; // @[:@134781.4]
  assign regs_147_reset = io_reset; // @[:@134782.4 RegFile.scala 76:16:@134789.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@134788.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@134792.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@134786.4]
  assign regs_148_clock = clock; // @[:@134795.4]
  assign regs_148_reset = io_reset; // @[:@134796.4 RegFile.scala 76:16:@134803.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@134802.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@134806.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@134800.4]
  assign regs_149_clock = clock; // @[:@134809.4]
  assign regs_149_reset = io_reset; // @[:@134810.4 RegFile.scala 76:16:@134817.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@134816.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@134820.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@134814.4]
  assign regs_150_clock = clock; // @[:@134823.4]
  assign regs_150_reset = io_reset; // @[:@134824.4 RegFile.scala 76:16:@134831.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@134830.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@134834.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@134828.4]
  assign regs_151_clock = clock; // @[:@134837.4]
  assign regs_151_reset = io_reset; // @[:@134838.4 RegFile.scala 76:16:@134845.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@134844.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@134848.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@134842.4]
  assign regs_152_clock = clock; // @[:@134851.4]
  assign regs_152_reset = io_reset; // @[:@134852.4 RegFile.scala 76:16:@134859.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@134858.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@134862.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@134856.4]
  assign regs_153_clock = clock; // @[:@134865.4]
  assign regs_153_reset = io_reset; // @[:@134866.4 RegFile.scala 76:16:@134873.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@134872.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@134876.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@134870.4]
  assign regs_154_clock = clock; // @[:@134879.4]
  assign regs_154_reset = io_reset; // @[:@134880.4 RegFile.scala 76:16:@134887.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@134886.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@134890.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@134884.4]
  assign regs_155_clock = clock; // @[:@134893.4]
  assign regs_155_reset = io_reset; // @[:@134894.4 RegFile.scala 76:16:@134901.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@134900.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@134904.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@134898.4]
  assign regs_156_clock = clock; // @[:@134907.4]
  assign regs_156_reset = io_reset; // @[:@134908.4 RegFile.scala 76:16:@134915.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@134914.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@134918.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@134912.4]
  assign regs_157_clock = clock; // @[:@134921.4]
  assign regs_157_reset = io_reset; // @[:@134922.4 RegFile.scala 76:16:@134929.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@134928.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@134932.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@134926.4]
  assign regs_158_clock = clock; // @[:@134935.4]
  assign regs_158_reset = io_reset; // @[:@134936.4 RegFile.scala 76:16:@134943.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@134942.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@134946.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@134940.4]
  assign regs_159_clock = clock; // @[:@134949.4]
  assign regs_159_reset = io_reset; // @[:@134950.4 RegFile.scala 76:16:@134957.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@134956.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@134960.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@134954.4]
  assign regs_160_clock = clock; // @[:@134963.4]
  assign regs_160_reset = io_reset; // @[:@134964.4 RegFile.scala 76:16:@134971.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@134970.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@134974.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@134968.4]
  assign regs_161_clock = clock; // @[:@134977.4]
  assign regs_161_reset = io_reset; // @[:@134978.4 RegFile.scala 76:16:@134985.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@134984.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@134988.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@134982.4]
  assign regs_162_clock = clock; // @[:@134991.4]
  assign regs_162_reset = io_reset; // @[:@134992.4 RegFile.scala 76:16:@134999.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@134998.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@135002.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@134996.4]
  assign regs_163_clock = clock; // @[:@135005.4]
  assign regs_163_reset = io_reset; // @[:@135006.4 RegFile.scala 76:16:@135013.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@135012.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@135016.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@135010.4]
  assign regs_164_clock = clock; // @[:@135019.4]
  assign regs_164_reset = io_reset; // @[:@135020.4 RegFile.scala 76:16:@135027.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@135026.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@135030.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@135024.4]
  assign regs_165_clock = clock; // @[:@135033.4]
  assign regs_165_reset = io_reset; // @[:@135034.4 RegFile.scala 76:16:@135041.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@135040.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@135044.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@135038.4]
  assign regs_166_clock = clock; // @[:@135047.4]
  assign regs_166_reset = io_reset; // @[:@135048.4 RegFile.scala 76:16:@135055.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@135054.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@135058.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@135052.4]
  assign regs_167_clock = clock; // @[:@135061.4]
  assign regs_167_reset = io_reset; // @[:@135062.4 RegFile.scala 76:16:@135069.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@135068.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@135072.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@135066.4]
  assign regs_168_clock = clock; // @[:@135075.4]
  assign regs_168_reset = io_reset; // @[:@135076.4 RegFile.scala 76:16:@135083.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@135082.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@135086.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@135080.4]
  assign regs_169_clock = clock; // @[:@135089.4]
  assign regs_169_reset = io_reset; // @[:@135090.4 RegFile.scala 76:16:@135097.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@135096.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@135100.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@135094.4]
  assign regs_170_clock = clock; // @[:@135103.4]
  assign regs_170_reset = io_reset; // @[:@135104.4 RegFile.scala 76:16:@135111.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@135110.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@135114.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@135108.4]
  assign regs_171_clock = clock; // @[:@135117.4]
  assign regs_171_reset = io_reset; // @[:@135118.4 RegFile.scala 76:16:@135125.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@135124.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@135128.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@135122.4]
  assign regs_172_clock = clock; // @[:@135131.4]
  assign regs_172_reset = io_reset; // @[:@135132.4 RegFile.scala 76:16:@135139.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@135138.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@135142.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@135136.4]
  assign regs_173_clock = clock; // @[:@135145.4]
  assign regs_173_reset = io_reset; // @[:@135146.4 RegFile.scala 76:16:@135153.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@135152.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@135156.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@135150.4]
  assign regs_174_clock = clock; // @[:@135159.4]
  assign regs_174_reset = io_reset; // @[:@135160.4 RegFile.scala 76:16:@135167.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@135166.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@135170.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@135164.4]
  assign regs_175_clock = clock; // @[:@135173.4]
  assign regs_175_reset = io_reset; // @[:@135174.4 RegFile.scala 76:16:@135181.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@135180.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@135184.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@135178.4]
  assign regs_176_clock = clock; // @[:@135187.4]
  assign regs_176_reset = io_reset; // @[:@135188.4 RegFile.scala 76:16:@135195.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@135194.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@135198.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@135192.4]
  assign regs_177_clock = clock; // @[:@135201.4]
  assign regs_177_reset = io_reset; // @[:@135202.4 RegFile.scala 76:16:@135209.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@135208.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@135212.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@135206.4]
  assign regs_178_clock = clock; // @[:@135215.4]
  assign regs_178_reset = io_reset; // @[:@135216.4 RegFile.scala 76:16:@135223.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@135222.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@135226.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@135220.4]
  assign regs_179_clock = clock; // @[:@135229.4]
  assign regs_179_reset = io_reset; // @[:@135230.4 RegFile.scala 76:16:@135237.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@135236.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@135240.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@135234.4]
  assign regs_180_clock = clock; // @[:@135243.4]
  assign regs_180_reset = io_reset; // @[:@135244.4 RegFile.scala 76:16:@135251.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@135250.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@135254.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@135248.4]
  assign regs_181_clock = clock; // @[:@135257.4]
  assign regs_181_reset = io_reset; // @[:@135258.4 RegFile.scala 76:16:@135265.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@135264.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@135268.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@135262.4]
  assign regs_182_clock = clock; // @[:@135271.4]
  assign regs_182_reset = io_reset; // @[:@135272.4 RegFile.scala 76:16:@135279.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@135278.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@135282.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@135276.4]
  assign regs_183_clock = clock; // @[:@135285.4]
  assign regs_183_reset = io_reset; // @[:@135286.4 RegFile.scala 76:16:@135293.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@135292.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@135296.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@135290.4]
  assign regs_184_clock = clock; // @[:@135299.4]
  assign regs_184_reset = io_reset; // @[:@135300.4 RegFile.scala 76:16:@135307.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@135306.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@135310.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@135304.4]
  assign regs_185_clock = clock; // @[:@135313.4]
  assign regs_185_reset = io_reset; // @[:@135314.4 RegFile.scala 76:16:@135321.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@135320.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@135324.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@135318.4]
  assign regs_186_clock = clock; // @[:@135327.4]
  assign regs_186_reset = io_reset; // @[:@135328.4 RegFile.scala 76:16:@135335.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@135334.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@135338.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@135332.4]
  assign regs_187_clock = clock; // @[:@135341.4]
  assign regs_187_reset = io_reset; // @[:@135342.4 RegFile.scala 76:16:@135349.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@135348.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@135352.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@135346.4]
  assign regs_188_clock = clock; // @[:@135355.4]
  assign regs_188_reset = io_reset; // @[:@135356.4 RegFile.scala 76:16:@135363.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@135362.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@135366.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@135360.4]
  assign regs_189_clock = clock; // @[:@135369.4]
  assign regs_189_reset = io_reset; // @[:@135370.4 RegFile.scala 76:16:@135377.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@135376.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@135380.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@135374.4]
  assign regs_190_clock = clock; // @[:@135383.4]
  assign regs_190_reset = io_reset; // @[:@135384.4 RegFile.scala 76:16:@135391.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@135390.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@135394.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@135388.4]
  assign regs_191_clock = clock; // @[:@135397.4]
  assign regs_191_reset = io_reset; // @[:@135398.4 RegFile.scala 76:16:@135405.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@135404.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@135408.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@135402.4]
  assign regs_192_clock = clock; // @[:@135411.4]
  assign regs_192_reset = io_reset; // @[:@135412.4 RegFile.scala 76:16:@135419.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@135418.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@135422.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@135416.4]
  assign regs_193_clock = clock; // @[:@135425.4]
  assign regs_193_reset = io_reset; // @[:@135426.4 RegFile.scala 76:16:@135433.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@135432.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@135436.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@135430.4]
  assign regs_194_clock = clock; // @[:@135439.4]
  assign regs_194_reset = io_reset; // @[:@135440.4 RegFile.scala 76:16:@135447.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@135446.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@135450.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@135444.4]
  assign regs_195_clock = clock; // @[:@135453.4]
  assign regs_195_reset = io_reset; // @[:@135454.4 RegFile.scala 76:16:@135461.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@135460.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@135464.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@135458.4]
  assign regs_196_clock = clock; // @[:@135467.4]
  assign regs_196_reset = io_reset; // @[:@135468.4 RegFile.scala 76:16:@135475.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@135474.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@135478.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@135472.4]
  assign regs_197_clock = clock; // @[:@135481.4]
  assign regs_197_reset = io_reset; // @[:@135482.4 RegFile.scala 76:16:@135489.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@135488.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@135492.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@135486.4]
  assign regs_198_clock = clock; // @[:@135495.4]
  assign regs_198_reset = io_reset; // @[:@135496.4 RegFile.scala 76:16:@135503.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@135502.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@135506.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@135500.4]
  assign regs_199_clock = clock; // @[:@135509.4]
  assign regs_199_reset = io_reset; // @[:@135510.4 RegFile.scala 76:16:@135517.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@135516.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@135520.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@135514.4]
  assign regs_200_clock = clock; // @[:@135523.4]
  assign regs_200_reset = io_reset; // @[:@135524.4 RegFile.scala 76:16:@135531.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@135530.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@135534.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@135528.4]
  assign regs_201_clock = clock; // @[:@135537.4]
  assign regs_201_reset = io_reset; // @[:@135538.4 RegFile.scala 76:16:@135545.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@135544.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@135548.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@135542.4]
  assign regs_202_clock = clock; // @[:@135551.4]
  assign regs_202_reset = io_reset; // @[:@135552.4 RegFile.scala 76:16:@135559.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@135558.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@135562.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@135556.4]
  assign regs_203_clock = clock; // @[:@135565.4]
  assign regs_203_reset = io_reset; // @[:@135566.4 RegFile.scala 76:16:@135573.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@135572.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@135576.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@135570.4]
  assign regs_204_clock = clock; // @[:@135579.4]
  assign regs_204_reset = io_reset; // @[:@135580.4 RegFile.scala 76:16:@135587.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@135586.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@135590.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@135584.4]
  assign regs_205_clock = clock; // @[:@135593.4]
  assign regs_205_reset = io_reset; // @[:@135594.4 RegFile.scala 76:16:@135601.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@135600.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@135604.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@135598.4]
  assign regs_206_clock = clock; // @[:@135607.4]
  assign regs_206_reset = io_reset; // @[:@135608.4 RegFile.scala 76:16:@135615.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@135614.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@135618.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@135612.4]
  assign regs_207_clock = clock; // @[:@135621.4]
  assign regs_207_reset = io_reset; // @[:@135622.4 RegFile.scala 76:16:@135629.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@135628.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@135632.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@135626.4]
  assign regs_208_clock = clock; // @[:@135635.4]
  assign regs_208_reset = io_reset; // @[:@135636.4 RegFile.scala 76:16:@135643.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@135642.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@135646.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@135640.4]
  assign regs_209_clock = clock; // @[:@135649.4]
  assign regs_209_reset = io_reset; // @[:@135650.4 RegFile.scala 76:16:@135657.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@135656.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@135660.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@135654.4]
  assign regs_210_clock = clock; // @[:@135663.4]
  assign regs_210_reset = io_reset; // @[:@135664.4 RegFile.scala 76:16:@135671.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@135670.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@135674.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@135668.4]
  assign regs_211_clock = clock; // @[:@135677.4]
  assign regs_211_reset = io_reset; // @[:@135678.4 RegFile.scala 76:16:@135685.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@135684.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@135688.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@135682.4]
  assign regs_212_clock = clock; // @[:@135691.4]
  assign regs_212_reset = io_reset; // @[:@135692.4 RegFile.scala 76:16:@135699.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@135698.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@135702.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@135696.4]
  assign regs_213_clock = clock; // @[:@135705.4]
  assign regs_213_reset = io_reset; // @[:@135706.4 RegFile.scala 76:16:@135713.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@135712.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@135716.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@135710.4]
  assign regs_214_clock = clock; // @[:@135719.4]
  assign regs_214_reset = io_reset; // @[:@135720.4 RegFile.scala 76:16:@135727.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@135726.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@135730.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@135724.4]
  assign regs_215_clock = clock; // @[:@135733.4]
  assign regs_215_reset = io_reset; // @[:@135734.4 RegFile.scala 76:16:@135741.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@135740.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@135744.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@135738.4]
  assign regs_216_clock = clock; // @[:@135747.4]
  assign regs_216_reset = io_reset; // @[:@135748.4 RegFile.scala 76:16:@135755.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@135754.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@135758.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@135752.4]
  assign regs_217_clock = clock; // @[:@135761.4]
  assign regs_217_reset = io_reset; // @[:@135762.4 RegFile.scala 76:16:@135769.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@135768.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@135772.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@135766.4]
  assign regs_218_clock = clock; // @[:@135775.4]
  assign regs_218_reset = io_reset; // @[:@135776.4 RegFile.scala 76:16:@135783.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@135782.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@135786.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@135780.4]
  assign regs_219_clock = clock; // @[:@135789.4]
  assign regs_219_reset = io_reset; // @[:@135790.4 RegFile.scala 76:16:@135797.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@135796.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@135800.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@135794.4]
  assign regs_220_clock = clock; // @[:@135803.4]
  assign regs_220_reset = io_reset; // @[:@135804.4 RegFile.scala 76:16:@135811.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@135810.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@135814.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@135808.4]
  assign regs_221_clock = clock; // @[:@135817.4]
  assign regs_221_reset = io_reset; // @[:@135818.4 RegFile.scala 76:16:@135825.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@135824.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@135828.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@135822.4]
  assign regs_222_clock = clock; // @[:@135831.4]
  assign regs_222_reset = io_reset; // @[:@135832.4 RegFile.scala 76:16:@135839.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@135838.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@135842.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@135836.4]
  assign regs_223_clock = clock; // @[:@135845.4]
  assign regs_223_reset = io_reset; // @[:@135846.4 RegFile.scala 76:16:@135853.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@135852.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@135856.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@135850.4]
  assign regs_224_clock = clock; // @[:@135859.4]
  assign regs_224_reset = io_reset; // @[:@135860.4 RegFile.scala 76:16:@135867.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@135866.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@135870.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@135864.4]
  assign regs_225_clock = clock; // @[:@135873.4]
  assign regs_225_reset = io_reset; // @[:@135874.4 RegFile.scala 76:16:@135881.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@135880.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@135884.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@135878.4]
  assign regs_226_clock = clock; // @[:@135887.4]
  assign regs_226_reset = io_reset; // @[:@135888.4 RegFile.scala 76:16:@135895.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@135894.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@135898.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@135892.4]
  assign regs_227_clock = clock; // @[:@135901.4]
  assign regs_227_reset = io_reset; // @[:@135902.4 RegFile.scala 76:16:@135909.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@135908.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@135912.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@135906.4]
  assign regs_228_clock = clock; // @[:@135915.4]
  assign regs_228_reset = io_reset; // @[:@135916.4 RegFile.scala 76:16:@135923.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@135922.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@135926.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@135920.4]
  assign regs_229_clock = clock; // @[:@135929.4]
  assign regs_229_reset = io_reset; // @[:@135930.4 RegFile.scala 76:16:@135937.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@135936.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@135940.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@135934.4]
  assign regs_230_clock = clock; // @[:@135943.4]
  assign regs_230_reset = io_reset; // @[:@135944.4 RegFile.scala 76:16:@135951.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@135950.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@135954.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@135948.4]
  assign regs_231_clock = clock; // @[:@135957.4]
  assign regs_231_reset = io_reset; // @[:@135958.4 RegFile.scala 76:16:@135965.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@135964.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@135968.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@135962.4]
  assign regs_232_clock = clock; // @[:@135971.4]
  assign regs_232_reset = io_reset; // @[:@135972.4 RegFile.scala 76:16:@135979.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@135978.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@135982.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@135976.4]
  assign regs_233_clock = clock; // @[:@135985.4]
  assign regs_233_reset = io_reset; // @[:@135986.4 RegFile.scala 76:16:@135993.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@135992.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@135996.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@135990.4]
  assign regs_234_clock = clock; // @[:@135999.4]
  assign regs_234_reset = io_reset; // @[:@136000.4 RegFile.scala 76:16:@136007.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@136006.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@136010.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@136004.4]
  assign regs_235_clock = clock; // @[:@136013.4]
  assign regs_235_reset = io_reset; // @[:@136014.4 RegFile.scala 76:16:@136021.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@136020.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@136024.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@136018.4]
  assign regs_236_clock = clock; // @[:@136027.4]
  assign regs_236_reset = io_reset; // @[:@136028.4 RegFile.scala 76:16:@136035.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@136034.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@136038.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@136032.4]
  assign regs_237_clock = clock; // @[:@136041.4]
  assign regs_237_reset = io_reset; // @[:@136042.4 RegFile.scala 76:16:@136049.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@136048.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@136052.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@136046.4]
  assign regs_238_clock = clock; // @[:@136055.4]
  assign regs_238_reset = io_reset; // @[:@136056.4 RegFile.scala 76:16:@136063.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@136062.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@136066.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@136060.4]
  assign regs_239_clock = clock; // @[:@136069.4]
  assign regs_239_reset = io_reset; // @[:@136070.4 RegFile.scala 76:16:@136077.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@136076.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@136080.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@136074.4]
  assign regs_240_clock = clock; // @[:@136083.4]
  assign regs_240_reset = io_reset; // @[:@136084.4 RegFile.scala 76:16:@136091.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@136090.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@136094.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@136088.4]
  assign regs_241_clock = clock; // @[:@136097.4]
  assign regs_241_reset = io_reset; // @[:@136098.4 RegFile.scala 76:16:@136105.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@136104.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@136108.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@136102.4]
  assign regs_242_clock = clock; // @[:@136111.4]
  assign regs_242_reset = io_reset; // @[:@136112.4 RegFile.scala 76:16:@136119.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@136118.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@136122.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@136116.4]
  assign regs_243_clock = clock; // @[:@136125.4]
  assign regs_243_reset = io_reset; // @[:@136126.4 RegFile.scala 76:16:@136133.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@136132.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@136136.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@136130.4]
  assign regs_244_clock = clock; // @[:@136139.4]
  assign regs_244_reset = io_reset; // @[:@136140.4 RegFile.scala 76:16:@136147.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@136146.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@136150.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@136144.4]
  assign regs_245_clock = clock; // @[:@136153.4]
  assign regs_245_reset = io_reset; // @[:@136154.4 RegFile.scala 76:16:@136161.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@136160.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@136164.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@136158.4]
  assign regs_246_clock = clock; // @[:@136167.4]
  assign regs_246_reset = io_reset; // @[:@136168.4 RegFile.scala 76:16:@136175.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@136174.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@136178.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@136172.4]
  assign regs_247_clock = clock; // @[:@136181.4]
  assign regs_247_reset = io_reset; // @[:@136182.4 RegFile.scala 76:16:@136189.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@136188.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@136192.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@136186.4]
  assign regs_248_clock = clock; // @[:@136195.4]
  assign regs_248_reset = io_reset; // @[:@136196.4 RegFile.scala 76:16:@136203.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@136202.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@136206.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@136200.4]
  assign regs_249_clock = clock; // @[:@136209.4]
  assign regs_249_reset = io_reset; // @[:@136210.4 RegFile.scala 76:16:@136217.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@136216.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@136220.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@136214.4]
  assign regs_250_clock = clock; // @[:@136223.4]
  assign regs_250_reset = io_reset; // @[:@136224.4 RegFile.scala 76:16:@136231.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@136230.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@136234.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@136228.4]
  assign regs_251_clock = clock; // @[:@136237.4]
  assign regs_251_reset = io_reset; // @[:@136238.4 RegFile.scala 76:16:@136245.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@136244.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@136248.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@136242.4]
  assign regs_252_clock = clock; // @[:@136251.4]
  assign regs_252_reset = io_reset; // @[:@136252.4 RegFile.scala 76:16:@136259.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@136258.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@136262.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@136256.4]
  assign regs_253_clock = clock; // @[:@136265.4]
  assign regs_253_reset = io_reset; // @[:@136266.4 RegFile.scala 76:16:@136273.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@136272.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@136276.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@136270.4]
  assign regs_254_clock = clock; // @[:@136279.4]
  assign regs_254_reset = io_reset; // @[:@136280.4 RegFile.scala 76:16:@136287.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@136286.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@136290.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@136284.4]
  assign regs_255_clock = clock; // @[:@136293.4]
  assign regs_255_reset = io_reset; // @[:@136294.4 RegFile.scala 76:16:@136301.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@136300.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@136304.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@136298.4]
  assign regs_256_clock = clock; // @[:@136307.4]
  assign regs_256_reset = io_reset; // @[:@136308.4 RegFile.scala 76:16:@136315.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@136314.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@136318.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@136312.4]
  assign regs_257_clock = clock; // @[:@136321.4]
  assign regs_257_reset = io_reset; // @[:@136322.4 RegFile.scala 76:16:@136329.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@136328.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@136332.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@136326.4]
  assign regs_258_clock = clock; // @[:@136335.4]
  assign regs_258_reset = io_reset; // @[:@136336.4 RegFile.scala 76:16:@136343.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@136342.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@136346.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@136340.4]
  assign regs_259_clock = clock; // @[:@136349.4]
  assign regs_259_reset = io_reset; // @[:@136350.4 RegFile.scala 76:16:@136357.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@136356.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@136360.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@136354.4]
  assign regs_260_clock = clock; // @[:@136363.4]
  assign regs_260_reset = io_reset; // @[:@136364.4 RegFile.scala 76:16:@136371.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@136370.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@136374.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@136368.4]
  assign regs_261_clock = clock; // @[:@136377.4]
  assign regs_261_reset = io_reset; // @[:@136378.4 RegFile.scala 76:16:@136385.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@136384.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@136388.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@136382.4]
  assign regs_262_clock = clock; // @[:@136391.4]
  assign regs_262_reset = io_reset; // @[:@136392.4 RegFile.scala 76:16:@136399.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@136398.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@136402.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@136396.4]
  assign regs_263_clock = clock; // @[:@136405.4]
  assign regs_263_reset = io_reset; // @[:@136406.4 RegFile.scala 76:16:@136413.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@136412.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@136416.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@136410.4]
  assign regs_264_clock = clock; // @[:@136419.4]
  assign regs_264_reset = io_reset; // @[:@136420.4 RegFile.scala 76:16:@136427.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@136426.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@136430.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@136424.4]
  assign regs_265_clock = clock; // @[:@136433.4]
  assign regs_265_reset = io_reset; // @[:@136434.4 RegFile.scala 76:16:@136441.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@136440.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@136444.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@136438.4]
  assign regs_266_clock = clock; // @[:@136447.4]
  assign regs_266_reset = io_reset; // @[:@136448.4 RegFile.scala 76:16:@136455.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@136454.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@136458.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@136452.4]
  assign regs_267_clock = clock; // @[:@136461.4]
  assign regs_267_reset = io_reset; // @[:@136462.4 RegFile.scala 76:16:@136469.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@136468.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@136472.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@136466.4]
  assign regs_268_clock = clock; // @[:@136475.4]
  assign regs_268_reset = io_reset; // @[:@136476.4 RegFile.scala 76:16:@136483.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@136482.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@136486.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@136480.4]
  assign regs_269_clock = clock; // @[:@136489.4]
  assign regs_269_reset = io_reset; // @[:@136490.4 RegFile.scala 76:16:@136497.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@136496.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@136500.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@136494.4]
  assign regs_270_clock = clock; // @[:@136503.4]
  assign regs_270_reset = io_reset; // @[:@136504.4 RegFile.scala 76:16:@136511.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@136510.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@136514.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@136508.4]
  assign regs_271_clock = clock; // @[:@136517.4]
  assign regs_271_reset = io_reset; // @[:@136518.4 RegFile.scala 76:16:@136525.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@136524.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@136528.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@136522.4]
  assign regs_272_clock = clock; // @[:@136531.4]
  assign regs_272_reset = io_reset; // @[:@136532.4 RegFile.scala 76:16:@136539.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@136538.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@136542.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@136536.4]
  assign regs_273_clock = clock; // @[:@136545.4]
  assign regs_273_reset = io_reset; // @[:@136546.4 RegFile.scala 76:16:@136553.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@136552.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@136556.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@136550.4]
  assign regs_274_clock = clock; // @[:@136559.4]
  assign regs_274_reset = io_reset; // @[:@136560.4 RegFile.scala 76:16:@136567.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@136566.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@136570.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@136564.4]
  assign regs_275_clock = clock; // @[:@136573.4]
  assign regs_275_reset = io_reset; // @[:@136574.4 RegFile.scala 76:16:@136581.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@136580.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@136584.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@136578.4]
  assign regs_276_clock = clock; // @[:@136587.4]
  assign regs_276_reset = io_reset; // @[:@136588.4 RegFile.scala 76:16:@136595.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@136594.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@136598.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@136592.4]
  assign regs_277_clock = clock; // @[:@136601.4]
  assign regs_277_reset = io_reset; // @[:@136602.4 RegFile.scala 76:16:@136609.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@136608.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@136612.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@136606.4]
  assign regs_278_clock = clock; // @[:@136615.4]
  assign regs_278_reset = io_reset; // @[:@136616.4 RegFile.scala 76:16:@136623.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@136622.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@136626.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@136620.4]
  assign regs_279_clock = clock; // @[:@136629.4]
  assign regs_279_reset = io_reset; // @[:@136630.4 RegFile.scala 76:16:@136637.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@136636.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@136640.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@136634.4]
  assign regs_280_clock = clock; // @[:@136643.4]
  assign regs_280_reset = io_reset; // @[:@136644.4 RegFile.scala 76:16:@136651.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@136650.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@136654.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@136648.4]
  assign regs_281_clock = clock; // @[:@136657.4]
  assign regs_281_reset = io_reset; // @[:@136658.4 RegFile.scala 76:16:@136665.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@136664.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@136668.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@136662.4]
  assign regs_282_clock = clock; // @[:@136671.4]
  assign regs_282_reset = io_reset; // @[:@136672.4 RegFile.scala 76:16:@136679.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@136678.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@136682.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@136676.4]
  assign regs_283_clock = clock; // @[:@136685.4]
  assign regs_283_reset = io_reset; // @[:@136686.4 RegFile.scala 76:16:@136693.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@136692.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@136696.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@136690.4]
  assign regs_284_clock = clock; // @[:@136699.4]
  assign regs_284_reset = io_reset; // @[:@136700.4 RegFile.scala 76:16:@136707.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@136706.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@136710.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@136704.4]
  assign regs_285_clock = clock; // @[:@136713.4]
  assign regs_285_reset = io_reset; // @[:@136714.4 RegFile.scala 76:16:@136721.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@136720.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@136724.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@136718.4]
  assign regs_286_clock = clock; // @[:@136727.4]
  assign regs_286_reset = io_reset; // @[:@136728.4 RegFile.scala 76:16:@136735.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@136734.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@136738.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@136732.4]
  assign regs_287_clock = clock; // @[:@136741.4]
  assign regs_287_reset = io_reset; // @[:@136742.4 RegFile.scala 76:16:@136749.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@136748.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@136752.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@136746.4]
  assign regs_288_clock = clock; // @[:@136755.4]
  assign regs_288_reset = io_reset; // @[:@136756.4 RegFile.scala 76:16:@136763.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@136762.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@136766.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@136760.4]
  assign regs_289_clock = clock; // @[:@136769.4]
  assign regs_289_reset = io_reset; // @[:@136770.4 RegFile.scala 76:16:@136777.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@136776.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@136780.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@136774.4]
  assign regs_290_clock = clock; // @[:@136783.4]
  assign regs_290_reset = io_reset; // @[:@136784.4 RegFile.scala 76:16:@136791.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@136790.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@136794.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@136788.4]
  assign regs_291_clock = clock; // @[:@136797.4]
  assign regs_291_reset = io_reset; // @[:@136798.4 RegFile.scala 76:16:@136805.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@136804.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@136808.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@136802.4]
  assign regs_292_clock = clock; // @[:@136811.4]
  assign regs_292_reset = io_reset; // @[:@136812.4 RegFile.scala 76:16:@136819.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@136818.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@136822.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@136816.4]
  assign regs_293_clock = clock; // @[:@136825.4]
  assign regs_293_reset = io_reset; // @[:@136826.4 RegFile.scala 76:16:@136833.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@136832.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@136836.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@136830.4]
  assign regs_294_clock = clock; // @[:@136839.4]
  assign regs_294_reset = io_reset; // @[:@136840.4 RegFile.scala 76:16:@136847.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@136846.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@136850.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@136844.4]
  assign regs_295_clock = clock; // @[:@136853.4]
  assign regs_295_reset = io_reset; // @[:@136854.4 RegFile.scala 76:16:@136861.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@136860.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@136864.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@136858.4]
  assign regs_296_clock = clock; // @[:@136867.4]
  assign regs_296_reset = io_reset; // @[:@136868.4 RegFile.scala 76:16:@136875.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@136874.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@136878.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@136872.4]
  assign regs_297_clock = clock; // @[:@136881.4]
  assign regs_297_reset = io_reset; // @[:@136882.4 RegFile.scala 76:16:@136889.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@136888.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@136892.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@136886.4]
  assign regs_298_clock = clock; // @[:@136895.4]
  assign regs_298_reset = io_reset; // @[:@136896.4 RegFile.scala 76:16:@136903.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@136902.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@136906.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@136900.4]
  assign regs_299_clock = clock; // @[:@136909.4]
  assign regs_299_reset = io_reset; // @[:@136910.4 RegFile.scala 76:16:@136917.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@136916.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@136920.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@136914.4]
  assign regs_300_clock = clock; // @[:@136923.4]
  assign regs_300_reset = io_reset; // @[:@136924.4 RegFile.scala 76:16:@136931.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@136930.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@136934.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@136928.4]
  assign regs_301_clock = clock; // @[:@136937.4]
  assign regs_301_reset = io_reset; // @[:@136938.4 RegFile.scala 76:16:@136945.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@136944.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@136948.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@136942.4]
  assign regs_302_clock = clock; // @[:@136951.4]
  assign regs_302_reset = io_reset; // @[:@136952.4 RegFile.scala 76:16:@136959.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@136958.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@136962.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@136956.4]
  assign regs_303_clock = clock; // @[:@136965.4]
  assign regs_303_reset = io_reset; // @[:@136966.4 RegFile.scala 76:16:@136973.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@136972.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@136976.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@136970.4]
  assign regs_304_clock = clock; // @[:@136979.4]
  assign regs_304_reset = io_reset; // @[:@136980.4 RegFile.scala 76:16:@136987.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@136986.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@136990.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@136984.4]
  assign regs_305_clock = clock; // @[:@136993.4]
  assign regs_305_reset = io_reset; // @[:@136994.4 RegFile.scala 76:16:@137001.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@137000.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@137004.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@136998.4]
  assign regs_306_clock = clock; // @[:@137007.4]
  assign regs_306_reset = io_reset; // @[:@137008.4 RegFile.scala 76:16:@137015.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@137014.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@137018.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@137012.4]
  assign regs_307_clock = clock; // @[:@137021.4]
  assign regs_307_reset = io_reset; // @[:@137022.4 RegFile.scala 76:16:@137029.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@137028.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@137032.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@137026.4]
  assign regs_308_clock = clock; // @[:@137035.4]
  assign regs_308_reset = io_reset; // @[:@137036.4 RegFile.scala 76:16:@137043.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@137042.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@137046.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@137040.4]
  assign regs_309_clock = clock; // @[:@137049.4]
  assign regs_309_reset = io_reset; // @[:@137050.4 RegFile.scala 76:16:@137057.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@137056.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@137060.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@137054.4]
  assign regs_310_clock = clock; // @[:@137063.4]
  assign regs_310_reset = io_reset; // @[:@137064.4 RegFile.scala 76:16:@137071.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@137070.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@137074.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@137068.4]
  assign regs_311_clock = clock; // @[:@137077.4]
  assign regs_311_reset = io_reset; // @[:@137078.4 RegFile.scala 76:16:@137085.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@137084.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@137088.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@137082.4]
  assign regs_312_clock = clock; // @[:@137091.4]
  assign regs_312_reset = io_reset; // @[:@137092.4 RegFile.scala 76:16:@137099.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@137098.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@137102.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@137096.4]
  assign regs_313_clock = clock; // @[:@137105.4]
  assign regs_313_reset = io_reset; // @[:@137106.4 RegFile.scala 76:16:@137113.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@137112.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@137116.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@137110.4]
  assign regs_314_clock = clock; // @[:@137119.4]
  assign regs_314_reset = io_reset; // @[:@137120.4 RegFile.scala 76:16:@137127.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@137126.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@137130.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@137124.4]
  assign regs_315_clock = clock; // @[:@137133.4]
  assign regs_315_reset = io_reset; // @[:@137134.4 RegFile.scala 76:16:@137141.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@137140.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@137144.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@137138.4]
  assign regs_316_clock = clock; // @[:@137147.4]
  assign regs_316_reset = io_reset; // @[:@137148.4 RegFile.scala 76:16:@137155.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@137154.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@137158.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@137152.4]
  assign regs_317_clock = clock; // @[:@137161.4]
  assign regs_317_reset = io_reset; // @[:@137162.4 RegFile.scala 76:16:@137169.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@137168.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@137172.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@137166.4]
  assign regs_318_clock = clock; // @[:@137175.4]
  assign regs_318_reset = io_reset; // @[:@137176.4 RegFile.scala 76:16:@137183.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@137182.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@137186.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@137180.4]
  assign regs_319_clock = clock; // @[:@137189.4]
  assign regs_319_reset = io_reset; // @[:@137190.4 RegFile.scala 76:16:@137197.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@137196.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@137200.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@137194.4]
  assign regs_320_clock = clock; // @[:@137203.4]
  assign regs_320_reset = io_reset; // @[:@137204.4 RegFile.scala 76:16:@137211.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@137210.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@137214.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@137208.4]
  assign regs_321_clock = clock; // @[:@137217.4]
  assign regs_321_reset = io_reset; // @[:@137218.4 RegFile.scala 76:16:@137225.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@137224.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@137228.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@137222.4]
  assign regs_322_clock = clock; // @[:@137231.4]
  assign regs_322_reset = io_reset; // @[:@137232.4 RegFile.scala 76:16:@137239.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@137238.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@137242.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@137236.4]
  assign regs_323_clock = clock; // @[:@137245.4]
  assign regs_323_reset = io_reset; // @[:@137246.4 RegFile.scala 76:16:@137253.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@137252.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@137256.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@137250.4]
  assign regs_324_clock = clock; // @[:@137259.4]
  assign regs_324_reset = io_reset; // @[:@137260.4 RegFile.scala 76:16:@137267.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@137266.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@137270.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@137264.4]
  assign regs_325_clock = clock; // @[:@137273.4]
  assign regs_325_reset = io_reset; // @[:@137274.4 RegFile.scala 76:16:@137281.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@137280.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@137284.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@137278.4]
  assign regs_326_clock = clock; // @[:@137287.4]
  assign regs_326_reset = io_reset; // @[:@137288.4 RegFile.scala 76:16:@137295.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@137294.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@137298.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@137292.4]
  assign regs_327_clock = clock; // @[:@137301.4]
  assign regs_327_reset = io_reset; // @[:@137302.4 RegFile.scala 76:16:@137309.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@137308.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@137312.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@137306.4]
  assign regs_328_clock = clock; // @[:@137315.4]
  assign regs_328_reset = io_reset; // @[:@137316.4 RegFile.scala 76:16:@137323.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@137322.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@137326.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@137320.4]
  assign regs_329_clock = clock; // @[:@137329.4]
  assign regs_329_reset = io_reset; // @[:@137330.4 RegFile.scala 76:16:@137337.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@137336.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@137340.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@137334.4]
  assign regs_330_clock = clock; // @[:@137343.4]
  assign regs_330_reset = io_reset; // @[:@137344.4 RegFile.scala 76:16:@137351.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@137350.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@137354.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@137348.4]
  assign regs_331_clock = clock; // @[:@137357.4]
  assign regs_331_reset = io_reset; // @[:@137358.4 RegFile.scala 76:16:@137365.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@137364.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@137368.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@137362.4]
  assign regs_332_clock = clock; // @[:@137371.4]
  assign regs_332_reset = io_reset; // @[:@137372.4 RegFile.scala 76:16:@137379.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@137378.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@137382.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@137376.4]
  assign regs_333_clock = clock; // @[:@137385.4]
  assign regs_333_reset = io_reset; // @[:@137386.4 RegFile.scala 76:16:@137393.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@137392.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@137396.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@137390.4]
  assign regs_334_clock = clock; // @[:@137399.4]
  assign regs_334_reset = io_reset; // @[:@137400.4 RegFile.scala 76:16:@137407.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@137406.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@137410.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@137404.4]
  assign regs_335_clock = clock; // @[:@137413.4]
  assign regs_335_reset = io_reset; // @[:@137414.4 RegFile.scala 76:16:@137421.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@137420.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@137424.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@137418.4]
  assign regs_336_clock = clock; // @[:@137427.4]
  assign regs_336_reset = io_reset; // @[:@137428.4 RegFile.scala 76:16:@137435.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@137434.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@137438.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@137432.4]
  assign regs_337_clock = clock; // @[:@137441.4]
  assign regs_337_reset = io_reset; // @[:@137442.4 RegFile.scala 76:16:@137449.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@137448.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@137452.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@137446.4]
  assign regs_338_clock = clock; // @[:@137455.4]
  assign regs_338_reset = io_reset; // @[:@137456.4 RegFile.scala 76:16:@137463.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@137462.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@137466.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@137460.4]
  assign regs_339_clock = clock; // @[:@137469.4]
  assign regs_339_reset = io_reset; // @[:@137470.4 RegFile.scala 76:16:@137477.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@137476.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@137480.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@137474.4]
  assign regs_340_clock = clock; // @[:@137483.4]
  assign regs_340_reset = io_reset; // @[:@137484.4 RegFile.scala 76:16:@137491.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@137490.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@137494.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@137488.4]
  assign regs_341_clock = clock; // @[:@137497.4]
  assign regs_341_reset = io_reset; // @[:@137498.4 RegFile.scala 76:16:@137505.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@137504.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@137508.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@137502.4]
  assign regs_342_clock = clock; // @[:@137511.4]
  assign regs_342_reset = io_reset; // @[:@137512.4 RegFile.scala 76:16:@137519.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@137518.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@137522.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@137516.4]
  assign regs_343_clock = clock; // @[:@137525.4]
  assign regs_343_reset = io_reset; // @[:@137526.4 RegFile.scala 76:16:@137533.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@137532.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@137536.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@137530.4]
  assign regs_344_clock = clock; // @[:@137539.4]
  assign regs_344_reset = io_reset; // @[:@137540.4 RegFile.scala 76:16:@137547.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@137546.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@137550.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@137544.4]
  assign regs_345_clock = clock; // @[:@137553.4]
  assign regs_345_reset = io_reset; // @[:@137554.4 RegFile.scala 76:16:@137561.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@137560.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@137564.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@137558.4]
  assign regs_346_clock = clock; // @[:@137567.4]
  assign regs_346_reset = io_reset; // @[:@137568.4 RegFile.scala 76:16:@137575.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@137574.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@137578.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@137572.4]
  assign regs_347_clock = clock; // @[:@137581.4]
  assign regs_347_reset = io_reset; // @[:@137582.4 RegFile.scala 76:16:@137589.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@137588.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@137592.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@137586.4]
  assign regs_348_clock = clock; // @[:@137595.4]
  assign regs_348_reset = io_reset; // @[:@137596.4 RegFile.scala 76:16:@137603.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@137602.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@137606.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@137600.4]
  assign regs_349_clock = clock; // @[:@137609.4]
  assign regs_349_reset = io_reset; // @[:@137610.4 RegFile.scala 76:16:@137617.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@137616.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@137620.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@137614.4]
  assign regs_350_clock = clock; // @[:@137623.4]
  assign regs_350_reset = io_reset; // @[:@137624.4 RegFile.scala 76:16:@137631.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@137630.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@137634.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@137628.4]
  assign regs_351_clock = clock; // @[:@137637.4]
  assign regs_351_reset = io_reset; // @[:@137638.4 RegFile.scala 76:16:@137645.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@137644.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@137648.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@137642.4]
  assign regs_352_clock = clock; // @[:@137651.4]
  assign regs_352_reset = io_reset; // @[:@137652.4 RegFile.scala 76:16:@137659.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@137658.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@137662.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@137656.4]
  assign regs_353_clock = clock; // @[:@137665.4]
  assign regs_353_reset = io_reset; // @[:@137666.4 RegFile.scala 76:16:@137673.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@137672.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@137676.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@137670.4]
  assign regs_354_clock = clock; // @[:@137679.4]
  assign regs_354_reset = io_reset; // @[:@137680.4 RegFile.scala 76:16:@137687.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@137686.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@137690.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@137684.4]
  assign regs_355_clock = clock; // @[:@137693.4]
  assign regs_355_reset = io_reset; // @[:@137694.4 RegFile.scala 76:16:@137701.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@137700.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@137704.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@137698.4]
  assign regs_356_clock = clock; // @[:@137707.4]
  assign regs_356_reset = io_reset; // @[:@137708.4 RegFile.scala 76:16:@137715.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@137714.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@137718.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@137712.4]
  assign regs_357_clock = clock; // @[:@137721.4]
  assign regs_357_reset = io_reset; // @[:@137722.4 RegFile.scala 76:16:@137729.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@137728.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@137732.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@137726.4]
  assign regs_358_clock = clock; // @[:@137735.4]
  assign regs_358_reset = io_reset; // @[:@137736.4 RegFile.scala 76:16:@137743.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@137742.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@137746.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@137740.4]
  assign regs_359_clock = clock; // @[:@137749.4]
  assign regs_359_reset = io_reset; // @[:@137750.4 RegFile.scala 76:16:@137757.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@137756.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@137760.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@137754.4]
  assign regs_360_clock = clock; // @[:@137763.4]
  assign regs_360_reset = io_reset; // @[:@137764.4 RegFile.scala 76:16:@137771.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@137770.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@137774.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@137768.4]
  assign regs_361_clock = clock; // @[:@137777.4]
  assign regs_361_reset = io_reset; // @[:@137778.4 RegFile.scala 76:16:@137785.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@137784.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@137788.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@137782.4]
  assign regs_362_clock = clock; // @[:@137791.4]
  assign regs_362_reset = io_reset; // @[:@137792.4 RegFile.scala 76:16:@137799.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@137798.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@137802.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@137796.4]
  assign regs_363_clock = clock; // @[:@137805.4]
  assign regs_363_reset = io_reset; // @[:@137806.4 RegFile.scala 76:16:@137813.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@137812.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@137816.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@137810.4]
  assign regs_364_clock = clock; // @[:@137819.4]
  assign regs_364_reset = io_reset; // @[:@137820.4 RegFile.scala 76:16:@137827.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@137826.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@137830.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@137824.4]
  assign regs_365_clock = clock; // @[:@137833.4]
  assign regs_365_reset = io_reset; // @[:@137834.4 RegFile.scala 76:16:@137841.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@137840.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@137844.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@137838.4]
  assign regs_366_clock = clock; // @[:@137847.4]
  assign regs_366_reset = io_reset; // @[:@137848.4 RegFile.scala 76:16:@137855.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@137854.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@137858.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@137852.4]
  assign regs_367_clock = clock; // @[:@137861.4]
  assign regs_367_reset = io_reset; // @[:@137862.4 RegFile.scala 76:16:@137869.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@137868.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@137872.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@137866.4]
  assign regs_368_clock = clock; // @[:@137875.4]
  assign regs_368_reset = io_reset; // @[:@137876.4 RegFile.scala 76:16:@137883.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@137882.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@137886.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@137880.4]
  assign regs_369_clock = clock; // @[:@137889.4]
  assign regs_369_reset = io_reset; // @[:@137890.4 RegFile.scala 76:16:@137897.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@137896.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@137900.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@137894.4]
  assign regs_370_clock = clock; // @[:@137903.4]
  assign regs_370_reset = io_reset; // @[:@137904.4 RegFile.scala 76:16:@137911.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@137910.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@137914.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@137908.4]
  assign regs_371_clock = clock; // @[:@137917.4]
  assign regs_371_reset = io_reset; // @[:@137918.4 RegFile.scala 76:16:@137925.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@137924.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@137928.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@137922.4]
  assign regs_372_clock = clock; // @[:@137931.4]
  assign regs_372_reset = io_reset; // @[:@137932.4 RegFile.scala 76:16:@137939.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@137938.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@137942.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@137936.4]
  assign regs_373_clock = clock; // @[:@137945.4]
  assign regs_373_reset = io_reset; // @[:@137946.4 RegFile.scala 76:16:@137953.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@137952.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@137956.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@137950.4]
  assign regs_374_clock = clock; // @[:@137959.4]
  assign regs_374_reset = io_reset; // @[:@137960.4 RegFile.scala 76:16:@137967.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@137966.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@137970.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@137964.4]
  assign regs_375_clock = clock; // @[:@137973.4]
  assign regs_375_reset = io_reset; // @[:@137974.4 RegFile.scala 76:16:@137981.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@137980.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@137984.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@137978.4]
  assign regs_376_clock = clock; // @[:@137987.4]
  assign regs_376_reset = io_reset; // @[:@137988.4 RegFile.scala 76:16:@137995.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@137994.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@137998.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@137992.4]
  assign regs_377_clock = clock; // @[:@138001.4]
  assign regs_377_reset = io_reset; // @[:@138002.4 RegFile.scala 76:16:@138009.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@138008.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@138012.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@138006.4]
  assign regs_378_clock = clock; // @[:@138015.4]
  assign regs_378_reset = io_reset; // @[:@138016.4 RegFile.scala 76:16:@138023.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@138022.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@138026.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@138020.4]
  assign regs_379_clock = clock; // @[:@138029.4]
  assign regs_379_reset = io_reset; // @[:@138030.4 RegFile.scala 76:16:@138037.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@138036.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@138040.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@138034.4]
  assign regs_380_clock = clock; // @[:@138043.4]
  assign regs_380_reset = io_reset; // @[:@138044.4 RegFile.scala 76:16:@138051.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@138050.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@138054.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@138048.4]
  assign regs_381_clock = clock; // @[:@138057.4]
  assign regs_381_reset = io_reset; // @[:@138058.4 RegFile.scala 76:16:@138065.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@138064.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@138068.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@138062.4]
  assign regs_382_clock = clock; // @[:@138071.4]
  assign regs_382_reset = io_reset; // @[:@138072.4 RegFile.scala 76:16:@138079.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@138078.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@138082.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@138076.4]
  assign regs_383_clock = clock; // @[:@138085.4]
  assign regs_383_reset = io_reset; // @[:@138086.4 RegFile.scala 76:16:@138093.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@138092.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@138096.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@138090.4]
  assign regs_384_clock = clock; // @[:@138099.4]
  assign regs_384_reset = io_reset; // @[:@138100.4 RegFile.scala 76:16:@138107.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@138106.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@138110.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@138104.4]
  assign regs_385_clock = clock; // @[:@138113.4]
  assign regs_385_reset = io_reset; // @[:@138114.4 RegFile.scala 76:16:@138121.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@138120.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@138124.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@138118.4]
  assign regs_386_clock = clock; // @[:@138127.4]
  assign regs_386_reset = io_reset; // @[:@138128.4 RegFile.scala 76:16:@138135.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@138134.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@138138.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@138132.4]
  assign regs_387_clock = clock; // @[:@138141.4]
  assign regs_387_reset = io_reset; // @[:@138142.4 RegFile.scala 76:16:@138149.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@138148.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@138152.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@138146.4]
  assign regs_388_clock = clock; // @[:@138155.4]
  assign regs_388_reset = io_reset; // @[:@138156.4 RegFile.scala 76:16:@138163.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@138162.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@138166.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@138160.4]
  assign regs_389_clock = clock; // @[:@138169.4]
  assign regs_389_reset = io_reset; // @[:@138170.4 RegFile.scala 76:16:@138177.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@138176.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@138180.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@138174.4]
  assign regs_390_clock = clock; // @[:@138183.4]
  assign regs_390_reset = io_reset; // @[:@138184.4 RegFile.scala 76:16:@138191.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@138190.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@138194.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@138188.4]
  assign regs_391_clock = clock; // @[:@138197.4]
  assign regs_391_reset = io_reset; // @[:@138198.4 RegFile.scala 76:16:@138205.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@138204.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@138208.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@138202.4]
  assign regs_392_clock = clock; // @[:@138211.4]
  assign regs_392_reset = io_reset; // @[:@138212.4 RegFile.scala 76:16:@138219.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@138218.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@138222.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@138216.4]
  assign regs_393_clock = clock; // @[:@138225.4]
  assign regs_393_reset = io_reset; // @[:@138226.4 RegFile.scala 76:16:@138233.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@138232.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@138236.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@138230.4]
  assign regs_394_clock = clock; // @[:@138239.4]
  assign regs_394_reset = io_reset; // @[:@138240.4 RegFile.scala 76:16:@138247.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@138246.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@138250.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@138244.4]
  assign regs_395_clock = clock; // @[:@138253.4]
  assign regs_395_reset = io_reset; // @[:@138254.4 RegFile.scala 76:16:@138261.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@138260.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@138264.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@138258.4]
  assign regs_396_clock = clock; // @[:@138267.4]
  assign regs_396_reset = io_reset; // @[:@138268.4 RegFile.scala 76:16:@138275.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@138274.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@138278.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@138272.4]
  assign regs_397_clock = clock; // @[:@138281.4]
  assign regs_397_reset = io_reset; // @[:@138282.4 RegFile.scala 76:16:@138289.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@138288.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@138292.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@138286.4]
  assign regs_398_clock = clock; // @[:@138295.4]
  assign regs_398_reset = io_reset; // @[:@138296.4 RegFile.scala 76:16:@138303.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@138302.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@138306.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@138300.4]
  assign regs_399_clock = clock; // @[:@138309.4]
  assign regs_399_reset = io_reset; // @[:@138310.4 RegFile.scala 76:16:@138317.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@138316.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@138320.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@138314.4]
  assign regs_400_clock = clock; // @[:@138323.4]
  assign regs_400_reset = io_reset; // @[:@138324.4 RegFile.scala 76:16:@138331.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@138330.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@138334.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@138328.4]
  assign regs_401_clock = clock; // @[:@138337.4]
  assign regs_401_reset = io_reset; // @[:@138338.4 RegFile.scala 76:16:@138345.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@138344.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@138348.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@138342.4]
  assign regs_402_clock = clock; // @[:@138351.4]
  assign regs_402_reset = io_reset; // @[:@138352.4 RegFile.scala 76:16:@138359.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@138358.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@138362.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@138356.4]
  assign regs_403_clock = clock; // @[:@138365.4]
  assign regs_403_reset = io_reset; // @[:@138366.4 RegFile.scala 76:16:@138373.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@138372.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@138376.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@138370.4]
  assign regs_404_clock = clock; // @[:@138379.4]
  assign regs_404_reset = io_reset; // @[:@138380.4 RegFile.scala 76:16:@138387.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@138386.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@138390.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@138384.4]
  assign regs_405_clock = clock; // @[:@138393.4]
  assign regs_405_reset = io_reset; // @[:@138394.4 RegFile.scala 76:16:@138401.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@138400.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@138404.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@138398.4]
  assign regs_406_clock = clock; // @[:@138407.4]
  assign regs_406_reset = io_reset; // @[:@138408.4 RegFile.scala 76:16:@138415.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@138414.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@138418.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@138412.4]
  assign regs_407_clock = clock; // @[:@138421.4]
  assign regs_407_reset = io_reset; // @[:@138422.4 RegFile.scala 76:16:@138429.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@138428.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@138432.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@138426.4]
  assign regs_408_clock = clock; // @[:@138435.4]
  assign regs_408_reset = io_reset; // @[:@138436.4 RegFile.scala 76:16:@138443.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@138442.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@138446.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@138440.4]
  assign regs_409_clock = clock; // @[:@138449.4]
  assign regs_409_reset = io_reset; // @[:@138450.4 RegFile.scala 76:16:@138457.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@138456.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@138460.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@138454.4]
  assign regs_410_clock = clock; // @[:@138463.4]
  assign regs_410_reset = io_reset; // @[:@138464.4 RegFile.scala 76:16:@138471.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@138470.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@138474.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@138468.4]
  assign regs_411_clock = clock; // @[:@138477.4]
  assign regs_411_reset = io_reset; // @[:@138478.4 RegFile.scala 76:16:@138485.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@138484.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@138488.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@138482.4]
  assign regs_412_clock = clock; // @[:@138491.4]
  assign regs_412_reset = io_reset; // @[:@138492.4 RegFile.scala 76:16:@138499.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@138498.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@138502.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@138496.4]
  assign regs_413_clock = clock; // @[:@138505.4]
  assign regs_413_reset = io_reset; // @[:@138506.4 RegFile.scala 76:16:@138513.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@138512.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@138516.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@138510.4]
  assign regs_414_clock = clock; // @[:@138519.4]
  assign regs_414_reset = io_reset; // @[:@138520.4 RegFile.scala 76:16:@138527.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@138526.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@138530.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@138524.4]
  assign regs_415_clock = clock; // @[:@138533.4]
  assign regs_415_reset = io_reset; // @[:@138534.4 RegFile.scala 76:16:@138541.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@138540.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@138544.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@138538.4]
  assign regs_416_clock = clock; // @[:@138547.4]
  assign regs_416_reset = io_reset; // @[:@138548.4 RegFile.scala 76:16:@138555.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@138554.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@138558.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@138552.4]
  assign regs_417_clock = clock; // @[:@138561.4]
  assign regs_417_reset = io_reset; // @[:@138562.4 RegFile.scala 76:16:@138569.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@138568.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@138572.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@138566.4]
  assign regs_418_clock = clock; // @[:@138575.4]
  assign regs_418_reset = io_reset; // @[:@138576.4 RegFile.scala 76:16:@138583.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@138582.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@138586.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@138580.4]
  assign regs_419_clock = clock; // @[:@138589.4]
  assign regs_419_reset = io_reset; // @[:@138590.4 RegFile.scala 76:16:@138597.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@138596.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@138600.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@138594.4]
  assign regs_420_clock = clock; // @[:@138603.4]
  assign regs_420_reset = io_reset; // @[:@138604.4 RegFile.scala 76:16:@138611.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@138610.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@138614.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@138608.4]
  assign regs_421_clock = clock; // @[:@138617.4]
  assign regs_421_reset = io_reset; // @[:@138618.4 RegFile.scala 76:16:@138625.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@138624.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@138628.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@138622.4]
  assign regs_422_clock = clock; // @[:@138631.4]
  assign regs_422_reset = io_reset; // @[:@138632.4 RegFile.scala 76:16:@138639.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@138638.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@138642.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@138636.4]
  assign regs_423_clock = clock; // @[:@138645.4]
  assign regs_423_reset = io_reset; // @[:@138646.4 RegFile.scala 76:16:@138653.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@138652.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@138656.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@138650.4]
  assign regs_424_clock = clock; // @[:@138659.4]
  assign regs_424_reset = io_reset; // @[:@138660.4 RegFile.scala 76:16:@138667.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@138666.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@138670.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@138664.4]
  assign regs_425_clock = clock; // @[:@138673.4]
  assign regs_425_reset = io_reset; // @[:@138674.4 RegFile.scala 76:16:@138681.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@138680.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@138684.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@138678.4]
  assign regs_426_clock = clock; // @[:@138687.4]
  assign regs_426_reset = io_reset; // @[:@138688.4 RegFile.scala 76:16:@138695.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@138694.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@138698.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@138692.4]
  assign regs_427_clock = clock; // @[:@138701.4]
  assign regs_427_reset = io_reset; // @[:@138702.4 RegFile.scala 76:16:@138709.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@138708.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@138712.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@138706.4]
  assign regs_428_clock = clock; // @[:@138715.4]
  assign regs_428_reset = io_reset; // @[:@138716.4 RegFile.scala 76:16:@138723.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@138722.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@138726.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@138720.4]
  assign regs_429_clock = clock; // @[:@138729.4]
  assign regs_429_reset = io_reset; // @[:@138730.4 RegFile.scala 76:16:@138737.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@138736.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@138740.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@138734.4]
  assign regs_430_clock = clock; // @[:@138743.4]
  assign regs_430_reset = io_reset; // @[:@138744.4 RegFile.scala 76:16:@138751.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@138750.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@138754.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@138748.4]
  assign regs_431_clock = clock; // @[:@138757.4]
  assign regs_431_reset = io_reset; // @[:@138758.4 RegFile.scala 76:16:@138765.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@138764.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@138768.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@138762.4]
  assign regs_432_clock = clock; // @[:@138771.4]
  assign regs_432_reset = io_reset; // @[:@138772.4 RegFile.scala 76:16:@138779.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@138778.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@138782.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@138776.4]
  assign regs_433_clock = clock; // @[:@138785.4]
  assign regs_433_reset = io_reset; // @[:@138786.4 RegFile.scala 76:16:@138793.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@138792.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@138796.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@138790.4]
  assign regs_434_clock = clock; // @[:@138799.4]
  assign regs_434_reset = io_reset; // @[:@138800.4 RegFile.scala 76:16:@138807.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@138806.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@138810.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@138804.4]
  assign regs_435_clock = clock; // @[:@138813.4]
  assign regs_435_reset = io_reset; // @[:@138814.4 RegFile.scala 76:16:@138821.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@138820.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@138824.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@138818.4]
  assign regs_436_clock = clock; // @[:@138827.4]
  assign regs_436_reset = io_reset; // @[:@138828.4 RegFile.scala 76:16:@138835.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@138834.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@138838.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@138832.4]
  assign regs_437_clock = clock; // @[:@138841.4]
  assign regs_437_reset = io_reset; // @[:@138842.4 RegFile.scala 76:16:@138849.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@138848.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@138852.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@138846.4]
  assign regs_438_clock = clock; // @[:@138855.4]
  assign regs_438_reset = io_reset; // @[:@138856.4 RegFile.scala 76:16:@138863.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@138862.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@138866.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@138860.4]
  assign regs_439_clock = clock; // @[:@138869.4]
  assign regs_439_reset = io_reset; // @[:@138870.4 RegFile.scala 76:16:@138877.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@138876.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@138880.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@138874.4]
  assign regs_440_clock = clock; // @[:@138883.4]
  assign regs_440_reset = io_reset; // @[:@138884.4 RegFile.scala 76:16:@138891.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@138890.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@138894.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@138888.4]
  assign regs_441_clock = clock; // @[:@138897.4]
  assign regs_441_reset = io_reset; // @[:@138898.4 RegFile.scala 76:16:@138905.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@138904.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@138908.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@138902.4]
  assign regs_442_clock = clock; // @[:@138911.4]
  assign regs_442_reset = io_reset; // @[:@138912.4 RegFile.scala 76:16:@138919.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@138918.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@138922.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@138916.4]
  assign regs_443_clock = clock; // @[:@138925.4]
  assign regs_443_reset = io_reset; // @[:@138926.4 RegFile.scala 76:16:@138933.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@138932.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@138936.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@138930.4]
  assign regs_444_clock = clock; // @[:@138939.4]
  assign regs_444_reset = io_reset; // @[:@138940.4 RegFile.scala 76:16:@138947.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@138946.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@138950.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@138944.4]
  assign regs_445_clock = clock; // @[:@138953.4]
  assign regs_445_reset = io_reset; // @[:@138954.4 RegFile.scala 76:16:@138961.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@138960.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@138964.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@138958.4]
  assign regs_446_clock = clock; // @[:@138967.4]
  assign regs_446_reset = io_reset; // @[:@138968.4 RegFile.scala 76:16:@138975.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@138974.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@138978.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@138972.4]
  assign regs_447_clock = clock; // @[:@138981.4]
  assign regs_447_reset = io_reset; // @[:@138982.4 RegFile.scala 76:16:@138989.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@138988.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@138992.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@138986.4]
  assign regs_448_clock = clock; // @[:@138995.4]
  assign regs_448_reset = io_reset; // @[:@138996.4 RegFile.scala 76:16:@139003.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@139002.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@139006.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@139000.4]
  assign regs_449_clock = clock; // @[:@139009.4]
  assign regs_449_reset = io_reset; // @[:@139010.4 RegFile.scala 76:16:@139017.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@139016.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@139020.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@139014.4]
  assign regs_450_clock = clock; // @[:@139023.4]
  assign regs_450_reset = io_reset; // @[:@139024.4 RegFile.scala 76:16:@139031.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@139030.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@139034.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@139028.4]
  assign regs_451_clock = clock; // @[:@139037.4]
  assign regs_451_reset = io_reset; // @[:@139038.4 RegFile.scala 76:16:@139045.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@139044.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@139048.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@139042.4]
  assign regs_452_clock = clock; // @[:@139051.4]
  assign regs_452_reset = io_reset; // @[:@139052.4 RegFile.scala 76:16:@139059.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@139058.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@139062.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@139056.4]
  assign regs_453_clock = clock; // @[:@139065.4]
  assign regs_453_reset = io_reset; // @[:@139066.4 RegFile.scala 76:16:@139073.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@139072.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@139076.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@139070.4]
  assign regs_454_clock = clock; // @[:@139079.4]
  assign regs_454_reset = io_reset; // @[:@139080.4 RegFile.scala 76:16:@139087.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@139086.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@139090.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@139084.4]
  assign regs_455_clock = clock; // @[:@139093.4]
  assign regs_455_reset = io_reset; // @[:@139094.4 RegFile.scala 76:16:@139101.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@139100.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@139104.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@139098.4]
  assign regs_456_clock = clock; // @[:@139107.4]
  assign regs_456_reset = io_reset; // @[:@139108.4 RegFile.scala 76:16:@139115.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@139114.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@139118.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@139112.4]
  assign regs_457_clock = clock; // @[:@139121.4]
  assign regs_457_reset = io_reset; // @[:@139122.4 RegFile.scala 76:16:@139129.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@139128.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@139132.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@139126.4]
  assign regs_458_clock = clock; // @[:@139135.4]
  assign regs_458_reset = io_reset; // @[:@139136.4 RegFile.scala 76:16:@139143.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@139142.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@139146.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@139140.4]
  assign regs_459_clock = clock; // @[:@139149.4]
  assign regs_459_reset = io_reset; // @[:@139150.4 RegFile.scala 76:16:@139157.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@139156.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@139160.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@139154.4]
  assign regs_460_clock = clock; // @[:@139163.4]
  assign regs_460_reset = io_reset; // @[:@139164.4 RegFile.scala 76:16:@139171.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@139170.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@139174.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@139168.4]
  assign regs_461_clock = clock; // @[:@139177.4]
  assign regs_461_reset = io_reset; // @[:@139178.4 RegFile.scala 76:16:@139185.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@139184.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@139188.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@139182.4]
  assign regs_462_clock = clock; // @[:@139191.4]
  assign regs_462_reset = io_reset; // @[:@139192.4 RegFile.scala 76:16:@139199.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@139198.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@139202.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@139196.4]
  assign regs_463_clock = clock; // @[:@139205.4]
  assign regs_463_reset = io_reset; // @[:@139206.4 RegFile.scala 76:16:@139213.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@139212.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@139216.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@139210.4]
  assign regs_464_clock = clock; // @[:@139219.4]
  assign regs_464_reset = io_reset; // @[:@139220.4 RegFile.scala 76:16:@139227.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@139226.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@139230.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@139224.4]
  assign regs_465_clock = clock; // @[:@139233.4]
  assign regs_465_reset = io_reset; // @[:@139234.4 RegFile.scala 76:16:@139241.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@139240.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@139244.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@139238.4]
  assign regs_466_clock = clock; // @[:@139247.4]
  assign regs_466_reset = io_reset; // @[:@139248.4 RegFile.scala 76:16:@139255.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@139254.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@139258.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@139252.4]
  assign regs_467_clock = clock; // @[:@139261.4]
  assign regs_467_reset = io_reset; // @[:@139262.4 RegFile.scala 76:16:@139269.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@139268.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@139272.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@139266.4]
  assign regs_468_clock = clock; // @[:@139275.4]
  assign regs_468_reset = io_reset; // @[:@139276.4 RegFile.scala 76:16:@139283.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@139282.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@139286.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@139280.4]
  assign regs_469_clock = clock; // @[:@139289.4]
  assign regs_469_reset = io_reset; // @[:@139290.4 RegFile.scala 76:16:@139297.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@139296.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@139300.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@139294.4]
  assign regs_470_clock = clock; // @[:@139303.4]
  assign regs_470_reset = io_reset; // @[:@139304.4 RegFile.scala 76:16:@139311.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@139310.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@139314.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@139308.4]
  assign regs_471_clock = clock; // @[:@139317.4]
  assign regs_471_reset = io_reset; // @[:@139318.4 RegFile.scala 76:16:@139325.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@139324.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@139328.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@139322.4]
  assign regs_472_clock = clock; // @[:@139331.4]
  assign regs_472_reset = io_reset; // @[:@139332.4 RegFile.scala 76:16:@139339.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@139338.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@139342.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@139336.4]
  assign regs_473_clock = clock; // @[:@139345.4]
  assign regs_473_reset = io_reset; // @[:@139346.4 RegFile.scala 76:16:@139353.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@139352.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@139356.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@139350.4]
  assign regs_474_clock = clock; // @[:@139359.4]
  assign regs_474_reset = io_reset; // @[:@139360.4 RegFile.scala 76:16:@139367.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@139366.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@139370.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@139364.4]
  assign regs_475_clock = clock; // @[:@139373.4]
  assign regs_475_reset = io_reset; // @[:@139374.4 RegFile.scala 76:16:@139381.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@139380.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@139384.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@139378.4]
  assign regs_476_clock = clock; // @[:@139387.4]
  assign regs_476_reset = io_reset; // @[:@139388.4 RegFile.scala 76:16:@139395.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@139394.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@139398.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@139392.4]
  assign regs_477_clock = clock; // @[:@139401.4]
  assign regs_477_reset = io_reset; // @[:@139402.4 RegFile.scala 76:16:@139409.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@139408.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@139412.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@139406.4]
  assign regs_478_clock = clock; // @[:@139415.4]
  assign regs_478_reset = io_reset; // @[:@139416.4 RegFile.scala 76:16:@139423.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@139422.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@139426.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@139420.4]
  assign regs_479_clock = clock; // @[:@139429.4]
  assign regs_479_reset = io_reset; // @[:@139430.4 RegFile.scala 76:16:@139437.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@139436.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@139440.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@139434.4]
  assign regs_480_clock = clock; // @[:@139443.4]
  assign regs_480_reset = io_reset; // @[:@139444.4 RegFile.scala 76:16:@139451.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@139450.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@139454.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@139448.4]
  assign regs_481_clock = clock; // @[:@139457.4]
  assign regs_481_reset = io_reset; // @[:@139458.4 RegFile.scala 76:16:@139465.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@139464.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@139468.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@139462.4]
  assign regs_482_clock = clock; // @[:@139471.4]
  assign regs_482_reset = io_reset; // @[:@139472.4 RegFile.scala 76:16:@139479.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@139478.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@139482.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@139476.4]
  assign regs_483_clock = clock; // @[:@139485.4]
  assign regs_483_reset = io_reset; // @[:@139486.4 RegFile.scala 76:16:@139493.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@139492.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@139496.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@139490.4]
  assign regs_484_clock = clock; // @[:@139499.4]
  assign regs_484_reset = io_reset; // @[:@139500.4 RegFile.scala 76:16:@139507.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@139506.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@139510.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@139504.4]
  assign regs_485_clock = clock; // @[:@139513.4]
  assign regs_485_reset = io_reset; // @[:@139514.4 RegFile.scala 76:16:@139521.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@139520.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@139524.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@139518.4]
  assign regs_486_clock = clock; // @[:@139527.4]
  assign regs_486_reset = io_reset; // @[:@139528.4 RegFile.scala 76:16:@139535.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@139534.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@139538.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@139532.4]
  assign regs_487_clock = clock; // @[:@139541.4]
  assign regs_487_reset = io_reset; // @[:@139542.4 RegFile.scala 76:16:@139549.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@139548.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@139552.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@139546.4]
  assign regs_488_clock = clock; // @[:@139555.4]
  assign regs_488_reset = io_reset; // @[:@139556.4 RegFile.scala 76:16:@139563.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@139562.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@139566.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@139560.4]
  assign regs_489_clock = clock; // @[:@139569.4]
  assign regs_489_reset = io_reset; // @[:@139570.4 RegFile.scala 76:16:@139577.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@139576.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@139580.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@139574.4]
  assign regs_490_clock = clock; // @[:@139583.4]
  assign regs_490_reset = io_reset; // @[:@139584.4 RegFile.scala 76:16:@139591.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@139590.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@139594.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@139588.4]
  assign regs_491_clock = clock; // @[:@139597.4]
  assign regs_491_reset = io_reset; // @[:@139598.4 RegFile.scala 76:16:@139605.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@139604.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@139608.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@139602.4]
  assign regs_492_clock = clock; // @[:@139611.4]
  assign regs_492_reset = io_reset; // @[:@139612.4 RegFile.scala 76:16:@139619.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@139618.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@139622.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@139616.4]
  assign regs_493_clock = clock; // @[:@139625.4]
  assign regs_493_reset = io_reset; // @[:@139626.4 RegFile.scala 76:16:@139633.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@139632.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@139636.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@139630.4]
  assign regs_494_clock = clock; // @[:@139639.4]
  assign regs_494_reset = io_reset; // @[:@139640.4 RegFile.scala 76:16:@139647.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@139646.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@139650.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@139644.4]
  assign regs_495_clock = clock; // @[:@139653.4]
  assign regs_495_reset = io_reset; // @[:@139654.4 RegFile.scala 76:16:@139661.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@139660.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@139664.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@139658.4]
  assign regs_496_clock = clock; // @[:@139667.4]
  assign regs_496_reset = io_reset; // @[:@139668.4 RegFile.scala 76:16:@139675.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@139674.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@139678.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@139672.4]
  assign regs_497_clock = clock; // @[:@139681.4]
  assign regs_497_reset = io_reset; // @[:@139682.4 RegFile.scala 76:16:@139689.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@139688.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@139692.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@139686.4]
  assign regs_498_clock = clock; // @[:@139695.4]
  assign regs_498_reset = io_reset; // @[:@139696.4 RegFile.scala 76:16:@139703.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@139702.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@139706.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@139700.4]
  assign regs_499_clock = clock; // @[:@139709.4]
  assign regs_499_reset = io_reset; // @[:@139710.4 RegFile.scala 76:16:@139717.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@139716.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@139720.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@139714.4]
  assign regs_500_clock = clock; // @[:@139723.4]
  assign regs_500_reset = io_reset; // @[:@139724.4 RegFile.scala 76:16:@139731.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@139730.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@139734.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@139728.4]
  assign regs_501_clock = clock; // @[:@139737.4]
  assign regs_501_reset = io_reset; // @[:@139738.4 RegFile.scala 76:16:@139745.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@139744.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@139748.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@139742.4]
  assign regs_502_clock = clock; // @[:@139751.4]
  assign regs_502_reset = io_reset; // @[:@139752.4 RegFile.scala 76:16:@139759.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@139758.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@139762.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@139756.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@140271.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@140272.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@140273.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@140274.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@140275.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@140276.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@140277.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@140278.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@140279.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@140280.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@140281.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@140282.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@140283.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@140284.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@140285.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@140286.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@140287.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@140288.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@140289.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@140290.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@140291.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@140292.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@140293.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@140294.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@140295.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@140296.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@140297.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@140298.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@140299.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@140300.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@140301.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@140302.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@140303.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@140304.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@140305.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@140306.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@140307.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@140308.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@140309.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@140310.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@140311.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@140312.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@140313.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@140314.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@140315.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@140316.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@140317.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@140318.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@140319.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@140320.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@140321.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@140322.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@140323.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@140324.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@140325.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@140326.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@140327.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@140328.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@140329.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@140330.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@140331.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@140332.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@140333.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@140334.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@140335.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@140336.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@140337.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@140338.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@140339.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@140340.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@140341.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@140342.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@140343.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@140344.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@140345.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@140346.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@140347.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@140348.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@140349.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@140350.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@140351.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@140352.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@140353.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@140354.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@140355.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@140356.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@140357.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@140358.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@140359.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@140360.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@140361.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@140362.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@140363.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@140364.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@140365.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@140366.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@140367.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@140368.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@140369.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@140370.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@140371.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@140372.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@140373.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@140374.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@140375.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@140376.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@140377.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@140378.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@140379.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@140380.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@140381.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@140382.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@140383.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@140384.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@140385.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@140386.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@140387.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@140388.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@140389.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@140390.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@140391.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@140392.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@140393.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@140394.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@140395.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@140396.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@140397.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@140398.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@140399.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@140400.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@140401.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@140402.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@140403.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@140404.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@140405.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@140406.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@140407.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@140408.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@140409.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@140410.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@140411.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@140412.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@140413.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@140414.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@140415.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@140416.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@140417.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@140418.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@140419.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@140420.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@140421.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@140422.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@140423.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@140424.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@140425.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@140426.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@140427.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@140428.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@140429.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@140430.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@140431.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@140432.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@140433.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@140434.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@140435.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@140436.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@140437.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@140438.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@140439.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@140440.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@140441.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@140442.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@140443.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@140444.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@140445.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@140446.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@140447.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@140448.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@140449.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@140450.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@140451.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@140452.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@140453.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@140454.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@140455.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@140456.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@140457.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@140458.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@140459.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@140460.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@140461.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@140462.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@140463.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@140464.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@140465.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@140466.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@140467.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@140468.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@140469.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@140470.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@140471.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@140472.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@140473.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@140474.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@140475.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@140476.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@140477.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@140478.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@140479.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@140480.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@140481.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@140482.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@140483.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@140484.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@140485.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@140486.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@140487.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@140488.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@140489.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@140490.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@140491.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@140492.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@140493.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@140494.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@140495.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@140496.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@140497.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@140498.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@140499.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@140500.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@140501.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@140502.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@140503.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@140504.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@140505.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@140506.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@140507.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@140508.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@140509.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@140510.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@140511.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@140512.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@140513.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@140514.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@140515.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@140516.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@140517.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@140518.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@140519.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@140520.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@140521.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@140522.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@140523.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@140524.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@140525.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@140526.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@140527.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@140528.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@140529.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@140530.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@140531.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@140532.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@140533.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@140534.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@140535.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@140536.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@140537.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@140538.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@140539.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@140540.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@140541.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@140542.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@140543.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@140544.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@140545.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@140546.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@140547.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@140548.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@140549.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@140550.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@140551.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@140552.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@140553.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@140554.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@140555.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@140556.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@140557.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@140558.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@140559.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@140560.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@140561.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@140562.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@140563.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@140564.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@140565.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@140566.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@140567.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@140568.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@140569.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@140570.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@140571.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@140572.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@140573.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@140574.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@140575.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@140576.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@140577.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@140578.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@140579.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@140580.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@140581.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@140582.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@140583.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@140584.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@140585.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@140586.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@140587.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@140588.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@140589.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@140590.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@140591.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@140592.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@140593.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@140594.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@140595.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@140596.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@140597.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@140598.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@140599.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@140600.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@140601.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@140602.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@140603.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@140604.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@140605.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@140606.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@140607.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@140608.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@140609.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@140610.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@140611.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@140612.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@140613.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@140614.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@140615.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@140616.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@140617.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@140618.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@140619.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@140620.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@140621.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@140622.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@140623.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@140624.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@140625.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@140626.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@140627.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@140628.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@140629.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@140630.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@140631.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@140632.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@140633.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@140634.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@140635.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@140636.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@140637.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@140638.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@140639.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@140640.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@140641.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@140642.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@140643.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@140644.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@140645.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@140646.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@140647.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@140648.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@140649.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@140650.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@140651.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@140652.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@140653.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@140654.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@140655.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@140656.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@140657.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@140658.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@140659.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@140660.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@140661.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@140662.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@140663.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@140664.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@140665.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@140666.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@140667.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@140668.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@140669.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@140670.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@140671.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@140672.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@140673.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@140674.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@140675.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@140676.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@140677.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@140678.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@140679.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@140680.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@140681.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@140682.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@140683.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@140684.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@140685.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@140686.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@140687.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@140688.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@140689.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@140690.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@140691.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@140692.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@140693.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@140694.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@140695.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@140696.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@140697.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@140698.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@140699.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@140700.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@140701.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@140702.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@140703.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@140704.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@140705.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@140706.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@140707.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@140708.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@140709.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@140710.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@140711.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@140712.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@140713.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@140714.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@140715.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@140716.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@140717.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@140718.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@140719.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@140720.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@140721.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@140722.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@140723.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@140724.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@140725.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@140726.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@140727.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@140728.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@140729.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@140730.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@140731.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@140732.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@140733.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@140734.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@140735.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@140736.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@140737.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@140738.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@140739.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@140740.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@140741.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@140742.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@140743.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@140744.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@140745.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@140746.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@140747.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@140748.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@140749.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@140750.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@140751.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@140752.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@140753.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@140754.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@140755.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@140756.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@140757.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@140758.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@140759.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@140760.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@140761.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@140762.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@140763.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@140764.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@140765.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@140766.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@140767.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@140768.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@140769.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@140770.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@140771.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@140772.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@140773.4]
  assign rport_io_sel = io_raddr[8:0]; // @[RegFile.scala 106:18:@140774.4]
endmodule
module RetimeWrapper_927( // @[:@140798.2]
  input         clock, // @[:@140799.4]
  input         reset, // @[:@140800.4]
  input  [39:0] io_in, // @[:@140801.4]
  output [39:0] io_out // @[:@140801.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@140803.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@140803.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@140803.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@140803.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@140803.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@140803.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@140803.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@140816.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@140815.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@140814.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@140813.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@140812.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@140810.4]
endmodule
module FringeFF_503( // @[:@140818.2]
  input         clock, // @[:@140819.4]
  input         reset, // @[:@140820.4]
  input  [39:0] io_in, // @[:@140821.4]
  output [39:0] io_out, // @[:@140821.4]
  input         io_enable // @[:@140821.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@140824.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@140824.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@140824.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@140824.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@140829.4 package.scala 96:25:@140830.4]
  RetimeWrapper_927 RetimeWrapper ( // @[package.scala 93:22:@140824.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@140829.4 package.scala 96:25:@140830.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@140841.4]
  assign RetimeWrapper_clock = clock; // @[:@140825.4]
  assign RetimeWrapper_reset = reset; // @[:@140826.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@140827.4]
endmodule
module FringeCounter( // @[:@140843.2]
  input   clock, // @[:@140844.4]
  input   reset, // @[:@140845.4]
  input   io_enable, // @[:@140846.4]
  output  io_done // @[:@140846.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@140848.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@140848.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@140848.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@140848.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@140848.4]
  wire [40:0] count; // @[Cat.scala 30:58:@140855.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@140856.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@140857.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@140858.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@140860.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@140848.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@140855.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@140856.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@140857.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@140858.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@140860.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@140871.4]
  assign reg$_clock = clock; // @[:@140849.4]
  assign reg$_reset = reset; // @[:@140850.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@140862.6 FringeCounter.scala 37:15:@140865.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@140853.4]
endmodule
module FringeFF_504( // @[:@140905.2]
  input   clock, // @[:@140906.4]
  input   reset, // @[:@140907.4]
  input   io_in, // @[:@140908.4]
  input   io_reset, // @[:@140908.4]
  output  io_out, // @[:@140908.4]
  input   io_enable // @[:@140908.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@140911.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@140911.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@140911.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@140911.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@140911.4]
  wire  _T_18; // @[package.scala 96:25:@140916.4 package.scala 96:25:@140917.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@140922.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@140911.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@140916.4 package.scala 96:25:@140917.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@140922.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@140928.4]
  assign RetimeWrapper_clock = clock; // @[:@140912.4]
  assign RetimeWrapper_reset = reset; // @[:@140913.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@140915.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@140914.4]
endmodule
module Depulser( // @[:@140930.2]
  input   clock, // @[:@140931.4]
  input   reset, // @[:@140932.4]
  input   io_in, // @[:@140933.4]
  input   io_rst, // @[:@140933.4]
  output  io_out // @[:@140933.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@140935.4]
  wire  r_reset; // @[Depulser.scala 14:17:@140935.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@140935.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@140935.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@140935.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@140935.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@140935.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@140944.4]
  assign r_clock = clock; // @[:@140936.4]
  assign r_reset = reset; // @[:@140937.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@140939.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@140943.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@140942.4]
endmodule
module Fringe( // @[:@140946.2]
  input         clock, // @[:@140947.4]
  input         reset, // @[:@140948.4]
  input  [31:0] io_raddr, // @[:@140949.4]
  input         io_wen, // @[:@140949.4]
  input  [31:0] io_waddr, // @[:@140949.4]
  input  [63:0] io_wdata, // @[:@140949.4]
  output [63:0] io_rdata, // @[:@140949.4]
  output        io_enable, // @[:@140949.4]
  input         io_done, // @[:@140949.4]
  output        io_reset, // @[:@140949.4]
  output [63:0] io_argIns_0, // @[:@140949.4]
  output [63:0] io_argIns_1, // @[:@140949.4]
  input         io_argOuts_0_valid, // @[:@140949.4]
  input  [63:0] io_argOuts_0_bits, // @[:@140949.4]
  output        io_memStreams_stores_0_cmd_ready, // @[:@140949.4]
  input         io_memStreams_stores_0_cmd_valid, // @[:@140949.4]
  input  [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@140949.4]
  input  [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@140949.4]
  output        io_memStreams_stores_0_data_ready, // @[:@140949.4]
  input         io_memStreams_stores_0_data_valid, // @[:@140949.4]
  input  [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@140949.4]
  input         io_memStreams_stores_0_data_bits_wstrb, // @[:@140949.4]
  input         io_memStreams_stores_0_wresp_ready, // @[:@140949.4]
  output        io_memStreams_stores_0_wresp_valid, // @[:@140949.4]
  output        io_memStreams_stores_0_wresp_bits, // @[:@140949.4]
  input         io_dram_0_cmd_ready, // @[:@140949.4]
  output        io_dram_0_cmd_valid, // @[:@140949.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@140949.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@140949.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@140949.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@140949.4]
  input         io_dram_0_wdata_ready, // @[:@140949.4]
  output        io_dram_0_wdata_valid, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_0, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_1, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_2, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_3, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_4, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_5, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_6, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_7, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_8, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_9, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_10, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_11, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_12, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_13, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_14, // @[:@140949.4]
  output [31:0] io_dram_0_wdata_bits_wdata_15, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@140949.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@140949.4]
  output        io_dram_0_rresp_ready, // @[:@140949.4]
  output        io_dram_0_wresp_ready, // @[:@140949.4]
  input         io_dram_0_wresp_valid, // @[:@140949.4]
  input  [31:0] io_dram_0_wresp_bits_tag, // @[:@140949.4]
  input         io_dram_1_cmd_ready, // @[:@140949.4]
  output        io_dram_1_cmd_valid, // @[:@140949.4]
  output [63:0] io_dram_1_cmd_bits_addr, // @[:@140949.4]
  output [31:0] io_dram_1_cmd_bits_size, // @[:@140949.4]
  output        io_dram_1_cmd_bits_isWr, // @[:@140949.4]
  output [31:0] io_dram_1_cmd_bits_tag, // @[:@140949.4]
  input         io_dram_1_wdata_ready, // @[:@140949.4]
  output        io_dram_1_wdata_valid, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_0, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_1, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_2, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_3, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_4, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_5, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_6, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_7, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_8, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_9, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_10, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_11, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_12, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_13, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_14, // @[:@140949.4]
  output [31:0] io_dram_1_wdata_bits_wdata_15, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_0, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_1, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_2, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_3, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_4, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_5, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_6, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_7, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_8, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_9, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_10, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_11, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_12, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_13, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_14, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_15, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_16, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_17, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_18, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_19, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_20, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_21, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_22, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_23, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_24, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_25, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_26, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_27, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_28, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_29, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_30, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_31, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_32, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_33, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_34, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_35, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_36, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_37, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_38, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_39, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_40, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_41, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_42, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_43, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_44, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_45, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_46, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_47, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_48, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_49, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_50, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_51, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_52, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_53, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_54, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_55, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_56, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_57, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_58, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_59, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_60, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_61, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_62, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wstrb_63, // @[:@140949.4]
  output        io_dram_1_wdata_bits_wlast, // @[:@140949.4]
  output        io_dram_1_rresp_ready, // @[:@140949.4]
  output        io_dram_1_wresp_ready, // @[:@140949.4]
  input         io_dram_1_wresp_valid, // @[:@140949.4]
  input  [31:0] io_dram_1_wresp_bits_tag, // @[:@140949.4]
  input         io_dram_2_cmd_ready, // @[:@140949.4]
  output        io_dram_2_cmd_valid, // @[:@140949.4]
  output [63:0] io_dram_2_cmd_bits_addr, // @[:@140949.4]
  output [31:0] io_dram_2_cmd_bits_size, // @[:@140949.4]
  output        io_dram_2_cmd_bits_isWr, // @[:@140949.4]
  output [31:0] io_dram_2_cmd_bits_tag, // @[:@140949.4]
  input         io_dram_2_wdata_ready, // @[:@140949.4]
  output        io_dram_2_wdata_valid, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_0, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_1, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_2, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_3, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_4, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_5, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_6, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_7, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_8, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_9, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_10, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_11, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_12, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_13, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_14, // @[:@140949.4]
  output [31:0] io_dram_2_wdata_bits_wdata_15, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_0, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_1, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_2, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_3, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_4, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_5, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_6, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_7, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_8, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_9, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_10, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_11, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_12, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_13, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_14, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_15, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_16, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_17, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_18, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_19, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_20, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_21, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_22, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_23, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_24, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_25, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_26, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_27, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_28, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_29, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_30, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_31, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_32, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_33, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_34, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_35, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_36, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_37, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_38, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_39, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_40, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_41, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_42, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_43, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_44, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_45, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_46, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_47, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_48, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_49, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_50, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_51, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_52, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_53, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_54, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_55, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_56, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_57, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_58, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_59, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_60, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_61, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_62, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wstrb_63, // @[:@140949.4]
  output        io_dram_2_wdata_bits_wlast, // @[:@140949.4]
  output        io_dram_2_rresp_ready, // @[:@140949.4]
  output        io_dram_2_wresp_ready, // @[:@140949.4]
  input         io_dram_2_wresp_valid, // @[:@140949.4]
  input  [31:0] io_dram_2_wresp_bits_tag, // @[:@140949.4]
  input         io_dram_3_cmd_ready, // @[:@140949.4]
  output        io_dram_3_cmd_valid, // @[:@140949.4]
  output [63:0] io_dram_3_cmd_bits_addr, // @[:@140949.4]
  output [31:0] io_dram_3_cmd_bits_size, // @[:@140949.4]
  output        io_dram_3_cmd_bits_isWr, // @[:@140949.4]
  output [31:0] io_dram_3_cmd_bits_tag, // @[:@140949.4]
  input         io_dram_3_wdata_ready, // @[:@140949.4]
  output        io_dram_3_wdata_valid, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_0, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_1, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_2, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_3, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_4, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_5, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_6, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_7, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_8, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_9, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_10, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_11, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_12, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_13, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_14, // @[:@140949.4]
  output [31:0] io_dram_3_wdata_bits_wdata_15, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_0, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_1, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_2, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_3, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_4, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_5, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_6, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_7, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_8, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_9, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_10, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_11, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_12, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_13, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_14, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_15, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_16, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_17, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_18, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_19, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_20, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_21, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_22, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_23, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_24, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_25, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_26, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_27, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_28, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_29, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_30, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_31, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_32, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_33, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_34, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_35, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_36, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_37, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_38, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_39, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_40, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_41, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_42, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_43, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_44, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_45, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_46, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_47, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_48, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_49, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_50, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_51, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_52, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_53, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_54, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_55, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_56, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_57, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_58, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_59, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_60, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_61, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_62, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wstrb_63, // @[:@140949.4]
  output        io_dram_3_wdata_bits_wlast, // @[:@140949.4]
  output        io_dram_3_rresp_ready, // @[:@140949.4]
  output        io_dram_3_wresp_ready, // @[:@140949.4]
  input         io_dram_3_wresp_valid, // @[:@140949.4]
  input  [31:0] io_dram_3_wresp_bits_tag, // @[:@140949.4]
  input         io_heap_0_req_valid, // @[:@140949.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@140949.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@140949.4]
  output        io_heap_0_resp_valid, // @[:@140949.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@140949.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@140949.4]
);
  wire  dramArbs_0_clock; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_reset; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_enable; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@140955.4]
  wire [63:0] dramArbs_0_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_app_stores_0_wresp_ready; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_cmd_ready; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 91:25:@140955.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_ready; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_0_io_dram_wresp_valid; // @[Fringe.scala 91:25:@140955.4]
  wire [31:0] dramArbs_0_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@140955.4]
  wire  dramArbs_1_clock; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_reset; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_enable; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_cmd_ready; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 91:25:@141948.4]
  wire [63:0] dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_ready; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_1_io_dram_wresp_valid; // @[Fringe.scala 91:25:@141948.4]
  wire [31:0] dramArbs_1_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@141948.4]
  wire  dramArbs_2_clock; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_reset; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_enable; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_cmd_ready; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 91:25:@142908.4]
  wire [63:0] dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_ready; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_io_dram_wresp_valid; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_2_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_3_clock; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_reset; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_enable; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_cmd_ready; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 91:25:@143868.4]
  wire [63:0] dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_ready; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_io_dram_wresp_valid; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_3_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@143868.4]
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@144828.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@144828.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@144828.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@144828.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@144828.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@144828.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@144828.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@144828.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@144828.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@144828.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@144828.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@144828.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@144837.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@144837.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@144837.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@144837.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@144837.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@144837.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@144837.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@144837.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@144837.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@144837.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@144837.4]
  wire [63:0] regs_io_argIns_3; // @[Fringe.scala 116:20:@144837.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@144837.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@144837.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@144837.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@144837.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@146887.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@146887.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@146887.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@146887.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@146906.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@146906.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@146906.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@146906.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@146906.4]
  wire [63:0] _T_1020; // @[:@146864.4 :@146865.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@146866.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@146868.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@146870.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@146872.4]
  wire  _T_1025; // @[Fringe.scala 134:28:@146874.4]
  wire  _T_1029; // @[Fringe.scala 134:42:@146876.4]
  wire  _T_1030; // @[Fringe.scala 135:27:@146878.4]
  wire [63:0] _T_1040; // @[Fringe.scala 156:22:@146914.4]
  reg  _T_1047; // @[package.scala 152:20:@146917.4]
  reg [31:0] _RAND_0;
  wire  _T_1048; // @[package.scala 153:13:@146919.4]
  wire  _T_1049; // @[package.scala 153:8:@146920.4]
  wire  _T_1052; // @[Fringe.scala 160:55:@146924.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@146925.4]
  wire  _T_1055; // @[Fringe.scala 161:58:@146928.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@146929.4]
  wire [1:0] _T_1059; // @[Fringe.scala 162:57:@146931.4]
  wire [1:0] _T_1061; // @[Fringe.scala 162:34:@146932.4]
  wire [63:0] _T_1063; // @[Fringe.scala 163:30:@146934.4]
  wire [1:0] _T_1064; // @[Fringe.scala 171:37:@146937.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@146916.4 Fringe.scala 163:24:@146935.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@146916.4 Fringe.scala 162:28:@146933.4]
  wire [61:0] _T_1065; // @[Fringe.scala 171:37:@146938.4]
  wire  alloc; // @[Fringe.scala 202:38:@148568.4]
  wire  dealloc; // @[Fringe.scala 203:40:@148569.4]
  wire  _T_1569; // @[Fringe.scala 204:37:@148570.4]
  reg  _T_1572; // @[package.scala 152:20:@148571.4]
  reg [31:0] _RAND_1;
  wire  _T_1573; // @[package.scala 153:13:@148573.4]
  DRAMArbiter dramArbs_0 ( // @[Fringe.scala 91:25:@140955.4]
    .clock(dramArbs_0_clock),
    .reset(dramArbs_0_reset),
    .io_enable(dramArbs_0_io_enable),
    .io_app_stores_0_cmd_ready(dramArbs_0_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_0_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_0_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_0_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_0_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_0_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_0_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_0_io_app_stores_0_data_bits_wstrb),
    .io_app_stores_0_wresp_ready(dramArbs_0_io_app_stores_0_wresp_ready),
    .io_app_stores_0_wresp_valid(dramArbs_0_io_app_stores_0_wresp_valid),
    .io_app_stores_0_wresp_bits(dramArbs_0_io_app_stores_0_wresp_bits),
    .io_dram_cmd_ready(dramArbs_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_0_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_0_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_0_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_0_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_0_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_0_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_0_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_0_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_0_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_0_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_0_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_0_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_0_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_0_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_0_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_0_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_0_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_0_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_0_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_0_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_0_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_0_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_0_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_0_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_0_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_0_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_0_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_0_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_0_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_0_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_0_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_0_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_0_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_0_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_0_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_0_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_0_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_0_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_0_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_0_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_0_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_0_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_0_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_0_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_0_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_0_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_0_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_0_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_0_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_0_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_0_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_0_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_0_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_0_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_0_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_0_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_0_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_0_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_0_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_0_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_0_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_0_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_0_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_0_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_0_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_0_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_0_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_0_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_0_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_0_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_0_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_0_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_0_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_0_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_1 ( // @[Fringe.scala 91:25:@141948.4]
    .clock(dramArbs_1_clock),
    .reset(dramArbs_1_reset),
    .io_enable(dramArbs_1_io_enable),
    .io_dram_cmd_ready(dramArbs_1_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_1_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_1_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_1_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_1_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_1_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_1_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_1_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_1_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_1_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_1_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_1_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_1_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_1_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_1_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_1_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_1_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_1_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_1_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_1_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_1_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_1_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_1_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_1_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_1_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_1_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_1_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_1_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_1_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_1_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_1_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_1_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_1_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_1_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_1_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_1_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_1_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_1_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_1_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_1_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_1_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_1_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_1_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_1_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_1_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_1_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_1_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_1_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_1_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_1_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_1_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_1_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_1_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_1_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_1_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_1_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_1_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_1_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_1_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_1_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_1_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_1_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_1_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_1_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_1_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_1_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_1_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_1_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_1_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_1_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_1_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_1_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_1_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_1_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_1_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_1_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_1_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_1_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_1_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_1_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_1_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_1_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_1_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_1_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_1_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_1_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_1_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_1_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_1_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_1_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_1_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_1_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_1_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_2 ( // @[Fringe.scala 91:25:@142908.4]
    .clock(dramArbs_2_clock),
    .reset(dramArbs_2_reset),
    .io_enable(dramArbs_2_io_enable),
    .io_dram_cmd_ready(dramArbs_2_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_2_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_2_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_2_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_2_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_2_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_2_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_2_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_2_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_2_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_2_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_2_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_2_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_2_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_2_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_2_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_2_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_2_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_2_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_2_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_2_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_2_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_2_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_2_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_2_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_2_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_2_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_2_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_2_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_2_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_2_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_2_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_2_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_2_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_2_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_2_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_2_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_2_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_2_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_2_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_2_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_2_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_2_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_2_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_2_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_2_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_2_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_2_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_2_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_2_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_2_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_2_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_2_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_2_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_2_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_2_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_2_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_2_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_2_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_2_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_2_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_2_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_2_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_2_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_2_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_2_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_2_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_2_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_2_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_2_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_2_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_2_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_2_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_2_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_2_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_2_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_2_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_2_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_2_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_2_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_2_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_2_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_2_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_2_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_2_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_2_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_2_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_2_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_2_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_2_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_2_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_2_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_2_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_3 ( // @[Fringe.scala 91:25:@143868.4]
    .clock(dramArbs_3_clock),
    .reset(dramArbs_3_reset),
    .io_enable(dramArbs_3_io_enable),
    .io_dram_cmd_ready(dramArbs_3_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_3_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_3_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_3_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_3_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_3_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_3_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_3_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_3_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_3_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_3_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_3_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_3_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_3_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_3_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_3_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_3_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_3_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_3_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_3_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_3_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_3_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_3_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_3_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_3_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_3_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_3_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_3_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_3_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_3_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_3_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_3_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_3_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_3_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_3_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_3_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_3_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_3_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_3_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_3_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_3_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_3_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_3_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_3_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_3_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_3_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_3_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_3_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_3_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_3_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_3_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_3_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_3_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_3_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_3_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_3_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_3_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_3_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_3_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_3_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_3_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_3_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_3_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_3_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_3_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_3_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_3_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_3_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_3_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_3_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_3_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_3_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_3_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_3_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_3_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_3_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_3_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_3_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_3_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_3_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_3_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_3_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_3_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_3_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_3_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_3_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_3_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_3_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_3_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_3_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_3_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_3_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_3_io_dram_wresp_bits_tag)
  );
  DRAMHeap heap ( // @[Fringe.scala 107:20:@144828.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@144837.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@146887.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@146906.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_1020 = regs_io_argIns_1; // @[:@146864.4 :@146865.4]
  assign curStatus_done = _T_1020[0]; // @[Fringe.scala 133:45:@146866.4]
  assign curStatus_timeout = _T_1020[1]; // @[Fringe.scala 133:45:@146868.4]
  assign curStatus_allocDealloc = _T_1020[4:2]; // @[Fringe.scala 133:45:@146870.4]
  assign curStatus_sizeAddr = _T_1020[63:5]; // @[Fringe.scala 133:45:@146872.4]
  assign _T_1025 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@146874.4]
  assign _T_1029 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@146876.4]
  assign _T_1030 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@146878.4]
  assign _T_1040 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@146914.4]
  assign _T_1048 = _T_1047 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@146919.4]
  assign _T_1049 = heap_io_host_0_req_valid & _T_1048; // @[package.scala 153:8:@146920.4]
  assign _T_1052 = _T_1025 & depulser_io_out; // @[Fringe.scala 160:55:@146924.4]
  assign status_bits_done = depulser_io_out ? _T_1052 : curStatus_done; // @[Fringe.scala 160:26:@146925.4]
  assign _T_1055 = _T_1025 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@146928.4]
  assign status_bits_timeout = depulser_io_out ? _T_1055 : curStatus_timeout; // @[Fringe.scala 161:29:@146929.4]
  assign _T_1059 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@146931.4]
  assign _T_1061 = heap_io_host_0_req_valid ? _T_1059 : 2'h0; // @[Fringe.scala 162:34:@146932.4]
  assign _T_1063 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@146934.4]
  assign _T_1064 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@146937.4]
  assign status_bits_sizeAddr = _T_1063[58:0]; // @[Fringe.scala 158:20:@146916.4 Fringe.scala 163:24:@146935.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_1061}; // @[Fringe.scala 158:20:@146916.4 Fringe.scala 162:28:@146933.4]
  assign _T_1065 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@146938.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@148568.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@148569.4]
  assign _T_1569 = alloc | dealloc; // @[Fringe.scala 204:37:@148570.4]
  assign _T_1573 = _T_1572 ^ _T_1569; // @[package.scala 153:13:@148573.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@146862.4]
  assign io_enable = _T_1025 & _T_1029; // @[Fringe.scala 136:13:@146882.4]
  assign io_reset = _T_1030 | reset; // @[Fringe.scala 137:12:@146883.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@146904.4]
  assign io_argIns_1 = regs_io_argIns_3; // @[Fringe.scala 151:51:@146905.4]
  assign io_memStreams_stores_0_cmd_ready = dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 101:72:@141874.4]
  assign io_memStreams_stores_0_data_ready = dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 101:72:@141870.4]
  assign io_memStreams_stores_0_wresp_valid = dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 101:72:@141865.4]
  assign io_memStreams_stores_0_wresp_bits = dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 101:72:@141864.4]
  assign io_dram_0_cmd_valid = dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 195:72:@148066.4]
  assign io_dram_0_cmd_bits_addr = dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@148065.4]
  assign io_dram_0_cmd_bits_size = dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@148064.4]
  assign io_dram_0_cmd_bits_isWr = dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@148062.4]
  assign io_dram_0_cmd_bits_tag = dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@148061.4]
  assign io_dram_0_wdata_valid = dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 195:72:@148059.4]
  assign io_dram_0_wdata_bits_wdata_0 = dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@148043.4]
  assign io_dram_0_wdata_bits_wdata_1 = dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@148044.4]
  assign io_dram_0_wdata_bits_wdata_2 = dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@148045.4]
  assign io_dram_0_wdata_bits_wdata_3 = dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@148046.4]
  assign io_dram_0_wdata_bits_wdata_4 = dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@148047.4]
  assign io_dram_0_wdata_bits_wdata_5 = dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@148048.4]
  assign io_dram_0_wdata_bits_wdata_6 = dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@148049.4]
  assign io_dram_0_wdata_bits_wdata_7 = dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@148050.4]
  assign io_dram_0_wdata_bits_wdata_8 = dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@148051.4]
  assign io_dram_0_wdata_bits_wdata_9 = dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@148052.4]
  assign io_dram_0_wdata_bits_wdata_10 = dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@148053.4]
  assign io_dram_0_wdata_bits_wdata_11 = dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@148054.4]
  assign io_dram_0_wdata_bits_wdata_12 = dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@148055.4]
  assign io_dram_0_wdata_bits_wdata_13 = dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@148056.4]
  assign io_dram_0_wdata_bits_wdata_14 = dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@148057.4]
  assign io_dram_0_wdata_bits_wdata_15 = dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@148058.4]
  assign io_dram_0_wdata_bits_wstrb_0 = dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@147979.4]
  assign io_dram_0_wdata_bits_wstrb_1 = dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@147980.4]
  assign io_dram_0_wdata_bits_wstrb_2 = dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@147981.4]
  assign io_dram_0_wdata_bits_wstrb_3 = dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@147982.4]
  assign io_dram_0_wdata_bits_wstrb_4 = dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@147983.4]
  assign io_dram_0_wdata_bits_wstrb_5 = dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@147984.4]
  assign io_dram_0_wdata_bits_wstrb_6 = dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@147985.4]
  assign io_dram_0_wdata_bits_wstrb_7 = dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@147986.4]
  assign io_dram_0_wdata_bits_wstrb_8 = dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@147987.4]
  assign io_dram_0_wdata_bits_wstrb_9 = dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@147988.4]
  assign io_dram_0_wdata_bits_wstrb_10 = dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@147989.4]
  assign io_dram_0_wdata_bits_wstrb_11 = dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@147990.4]
  assign io_dram_0_wdata_bits_wstrb_12 = dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@147991.4]
  assign io_dram_0_wdata_bits_wstrb_13 = dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@147992.4]
  assign io_dram_0_wdata_bits_wstrb_14 = dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@147993.4]
  assign io_dram_0_wdata_bits_wstrb_15 = dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@147994.4]
  assign io_dram_0_wdata_bits_wstrb_16 = dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@147995.4]
  assign io_dram_0_wdata_bits_wstrb_17 = dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@147996.4]
  assign io_dram_0_wdata_bits_wstrb_18 = dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@147997.4]
  assign io_dram_0_wdata_bits_wstrb_19 = dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@147998.4]
  assign io_dram_0_wdata_bits_wstrb_20 = dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@147999.4]
  assign io_dram_0_wdata_bits_wstrb_21 = dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@148000.4]
  assign io_dram_0_wdata_bits_wstrb_22 = dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@148001.4]
  assign io_dram_0_wdata_bits_wstrb_23 = dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@148002.4]
  assign io_dram_0_wdata_bits_wstrb_24 = dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@148003.4]
  assign io_dram_0_wdata_bits_wstrb_25 = dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@148004.4]
  assign io_dram_0_wdata_bits_wstrb_26 = dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@148005.4]
  assign io_dram_0_wdata_bits_wstrb_27 = dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@148006.4]
  assign io_dram_0_wdata_bits_wstrb_28 = dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@148007.4]
  assign io_dram_0_wdata_bits_wstrb_29 = dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@148008.4]
  assign io_dram_0_wdata_bits_wstrb_30 = dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@148009.4]
  assign io_dram_0_wdata_bits_wstrb_31 = dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@148010.4]
  assign io_dram_0_wdata_bits_wstrb_32 = dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@148011.4]
  assign io_dram_0_wdata_bits_wstrb_33 = dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@148012.4]
  assign io_dram_0_wdata_bits_wstrb_34 = dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@148013.4]
  assign io_dram_0_wdata_bits_wstrb_35 = dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@148014.4]
  assign io_dram_0_wdata_bits_wstrb_36 = dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@148015.4]
  assign io_dram_0_wdata_bits_wstrb_37 = dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@148016.4]
  assign io_dram_0_wdata_bits_wstrb_38 = dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@148017.4]
  assign io_dram_0_wdata_bits_wstrb_39 = dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@148018.4]
  assign io_dram_0_wdata_bits_wstrb_40 = dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@148019.4]
  assign io_dram_0_wdata_bits_wstrb_41 = dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@148020.4]
  assign io_dram_0_wdata_bits_wstrb_42 = dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@148021.4]
  assign io_dram_0_wdata_bits_wstrb_43 = dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@148022.4]
  assign io_dram_0_wdata_bits_wstrb_44 = dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@148023.4]
  assign io_dram_0_wdata_bits_wstrb_45 = dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@148024.4]
  assign io_dram_0_wdata_bits_wstrb_46 = dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@148025.4]
  assign io_dram_0_wdata_bits_wstrb_47 = dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@148026.4]
  assign io_dram_0_wdata_bits_wstrb_48 = dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@148027.4]
  assign io_dram_0_wdata_bits_wstrb_49 = dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@148028.4]
  assign io_dram_0_wdata_bits_wstrb_50 = dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@148029.4]
  assign io_dram_0_wdata_bits_wstrb_51 = dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@148030.4]
  assign io_dram_0_wdata_bits_wstrb_52 = dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@148031.4]
  assign io_dram_0_wdata_bits_wstrb_53 = dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@148032.4]
  assign io_dram_0_wdata_bits_wstrb_54 = dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@148033.4]
  assign io_dram_0_wdata_bits_wstrb_55 = dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@148034.4]
  assign io_dram_0_wdata_bits_wstrb_56 = dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@148035.4]
  assign io_dram_0_wdata_bits_wstrb_57 = dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@148036.4]
  assign io_dram_0_wdata_bits_wstrb_58 = dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@148037.4]
  assign io_dram_0_wdata_bits_wstrb_59 = dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@148038.4]
  assign io_dram_0_wdata_bits_wstrb_60 = dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@148039.4]
  assign io_dram_0_wdata_bits_wstrb_61 = dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@148040.4]
  assign io_dram_0_wdata_bits_wstrb_62 = dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@148041.4]
  assign io_dram_0_wdata_bits_wstrb_63 = dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@148042.4]
  assign io_dram_0_wdata_bits_wlast = dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@147978.4]
  assign io_dram_0_rresp_ready = dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 195:72:@147977.4]
  assign io_dram_0_wresp_ready = dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 195:72:@147958.4]
  assign io_dram_1_cmd_valid = dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 195:72:@148178.4]
  assign io_dram_1_cmd_bits_addr = dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@148177.4]
  assign io_dram_1_cmd_bits_size = dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@148176.4]
  assign io_dram_1_cmd_bits_isWr = dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@148174.4]
  assign io_dram_1_cmd_bits_tag = dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@148173.4]
  assign io_dram_1_wdata_valid = dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 195:72:@148171.4]
  assign io_dram_1_wdata_bits_wdata_0 = dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@148155.4]
  assign io_dram_1_wdata_bits_wdata_1 = dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@148156.4]
  assign io_dram_1_wdata_bits_wdata_2 = dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@148157.4]
  assign io_dram_1_wdata_bits_wdata_3 = dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@148158.4]
  assign io_dram_1_wdata_bits_wdata_4 = dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@148159.4]
  assign io_dram_1_wdata_bits_wdata_5 = dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@148160.4]
  assign io_dram_1_wdata_bits_wdata_6 = dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@148161.4]
  assign io_dram_1_wdata_bits_wdata_7 = dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@148162.4]
  assign io_dram_1_wdata_bits_wdata_8 = dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@148163.4]
  assign io_dram_1_wdata_bits_wdata_9 = dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@148164.4]
  assign io_dram_1_wdata_bits_wdata_10 = dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@148165.4]
  assign io_dram_1_wdata_bits_wdata_11 = dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@148166.4]
  assign io_dram_1_wdata_bits_wdata_12 = dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@148167.4]
  assign io_dram_1_wdata_bits_wdata_13 = dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@148168.4]
  assign io_dram_1_wdata_bits_wdata_14 = dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@148169.4]
  assign io_dram_1_wdata_bits_wdata_15 = dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@148170.4]
  assign io_dram_1_wdata_bits_wstrb_0 = dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@148091.4]
  assign io_dram_1_wdata_bits_wstrb_1 = dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@148092.4]
  assign io_dram_1_wdata_bits_wstrb_2 = dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@148093.4]
  assign io_dram_1_wdata_bits_wstrb_3 = dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@148094.4]
  assign io_dram_1_wdata_bits_wstrb_4 = dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@148095.4]
  assign io_dram_1_wdata_bits_wstrb_5 = dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@148096.4]
  assign io_dram_1_wdata_bits_wstrb_6 = dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@148097.4]
  assign io_dram_1_wdata_bits_wstrb_7 = dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@148098.4]
  assign io_dram_1_wdata_bits_wstrb_8 = dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@148099.4]
  assign io_dram_1_wdata_bits_wstrb_9 = dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@148100.4]
  assign io_dram_1_wdata_bits_wstrb_10 = dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@148101.4]
  assign io_dram_1_wdata_bits_wstrb_11 = dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@148102.4]
  assign io_dram_1_wdata_bits_wstrb_12 = dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@148103.4]
  assign io_dram_1_wdata_bits_wstrb_13 = dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@148104.4]
  assign io_dram_1_wdata_bits_wstrb_14 = dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@148105.4]
  assign io_dram_1_wdata_bits_wstrb_15 = dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@148106.4]
  assign io_dram_1_wdata_bits_wstrb_16 = dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@148107.4]
  assign io_dram_1_wdata_bits_wstrb_17 = dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@148108.4]
  assign io_dram_1_wdata_bits_wstrb_18 = dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@148109.4]
  assign io_dram_1_wdata_bits_wstrb_19 = dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@148110.4]
  assign io_dram_1_wdata_bits_wstrb_20 = dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@148111.4]
  assign io_dram_1_wdata_bits_wstrb_21 = dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@148112.4]
  assign io_dram_1_wdata_bits_wstrb_22 = dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@148113.4]
  assign io_dram_1_wdata_bits_wstrb_23 = dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@148114.4]
  assign io_dram_1_wdata_bits_wstrb_24 = dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@148115.4]
  assign io_dram_1_wdata_bits_wstrb_25 = dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@148116.4]
  assign io_dram_1_wdata_bits_wstrb_26 = dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@148117.4]
  assign io_dram_1_wdata_bits_wstrb_27 = dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@148118.4]
  assign io_dram_1_wdata_bits_wstrb_28 = dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@148119.4]
  assign io_dram_1_wdata_bits_wstrb_29 = dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@148120.4]
  assign io_dram_1_wdata_bits_wstrb_30 = dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@148121.4]
  assign io_dram_1_wdata_bits_wstrb_31 = dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@148122.4]
  assign io_dram_1_wdata_bits_wstrb_32 = dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@148123.4]
  assign io_dram_1_wdata_bits_wstrb_33 = dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@148124.4]
  assign io_dram_1_wdata_bits_wstrb_34 = dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@148125.4]
  assign io_dram_1_wdata_bits_wstrb_35 = dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@148126.4]
  assign io_dram_1_wdata_bits_wstrb_36 = dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@148127.4]
  assign io_dram_1_wdata_bits_wstrb_37 = dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@148128.4]
  assign io_dram_1_wdata_bits_wstrb_38 = dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@148129.4]
  assign io_dram_1_wdata_bits_wstrb_39 = dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@148130.4]
  assign io_dram_1_wdata_bits_wstrb_40 = dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@148131.4]
  assign io_dram_1_wdata_bits_wstrb_41 = dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@148132.4]
  assign io_dram_1_wdata_bits_wstrb_42 = dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@148133.4]
  assign io_dram_1_wdata_bits_wstrb_43 = dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@148134.4]
  assign io_dram_1_wdata_bits_wstrb_44 = dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@148135.4]
  assign io_dram_1_wdata_bits_wstrb_45 = dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@148136.4]
  assign io_dram_1_wdata_bits_wstrb_46 = dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@148137.4]
  assign io_dram_1_wdata_bits_wstrb_47 = dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@148138.4]
  assign io_dram_1_wdata_bits_wstrb_48 = dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@148139.4]
  assign io_dram_1_wdata_bits_wstrb_49 = dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@148140.4]
  assign io_dram_1_wdata_bits_wstrb_50 = dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@148141.4]
  assign io_dram_1_wdata_bits_wstrb_51 = dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@148142.4]
  assign io_dram_1_wdata_bits_wstrb_52 = dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@148143.4]
  assign io_dram_1_wdata_bits_wstrb_53 = dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@148144.4]
  assign io_dram_1_wdata_bits_wstrb_54 = dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@148145.4]
  assign io_dram_1_wdata_bits_wstrb_55 = dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@148146.4]
  assign io_dram_1_wdata_bits_wstrb_56 = dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@148147.4]
  assign io_dram_1_wdata_bits_wstrb_57 = dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@148148.4]
  assign io_dram_1_wdata_bits_wstrb_58 = dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@148149.4]
  assign io_dram_1_wdata_bits_wstrb_59 = dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@148150.4]
  assign io_dram_1_wdata_bits_wstrb_60 = dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@148151.4]
  assign io_dram_1_wdata_bits_wstrb_61 = dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@148152.4]
  assign io_dram_1_wdata_bits_wstrb_62 = dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@148153.4]
  assign io_dram_1_wdata_bits_wstrb_63 = dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@148154.4]
  assign io_dram_1_wdata_bits_wlast = dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@148090.4]
  assign io_dram_1_rresp_ready = dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 195:72:@148089.4]
  assign io_dram_1_wresp_ready = dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 195:72:@148070.4]
  assign io_dram_2_cmd_valid = dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 195:72:@148290.4]
  assign io_dram_2_cmd_bits_addr = dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@148289.4]
  assign io_dram_2_cmd_bits_size = dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@148288.4]
  assign io_dram_2_cmd_bits_isWr = dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@148286.4]
  assign io_dram_2_cmd_bits_tag = dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@148285.4]
  assign io_dram_2_wdata_valid = dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 195:72:@148283.4]
  assign io_dram_2_wdata_bits_wdata_0 = dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@148267.4]
  assign io_dram_2_wdata_bits_wdata_1 = dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@148268.4]
  assign io_dram_2_wdata_bits_wdata_2 = dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@148269.4]
  assign io_dram_2_wdata_bits_wdata_3 = dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@148270.4]
  assign io_dram_2_wdata_bits_wdata_4 = dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@148271.4]
  assign io_dram_2_wdata_bits_wdata_5 = dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@148272.4]
  assign io_dram_2_wdata_bits_wdata_6 = dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@148273.4]
  assign io_dram_2_wdata_bits_wdata_7 = dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@148274.4]
  assign io_dram_2_wdata_bits_wdata_8 = dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@148275.4]
  assign io_dram_2_wdata_bits_wdata_9 = dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@148276.4]
  assign io_dram_2_wdata_bits_wdata_10 = dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@148277.4]
  assign io_dram_2_wdata_bits_wdata_11 = dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@148278.4]
  assign io_dram_2_wdata_bits_wdata_12 = dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@148279.4]
  assign io_dram_2_wdata_bits_wdata_13 = dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@148280.4]
  assign io_dram_2_wdata_bits_wdata_14 = dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@148281.4]
  assign io_dram_2_wdata_bits_wdata_15 = dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@148282.4]
  assign io_dram_2_wdata_bits_wstrb_0 = dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@148203.4]
  assign io_dram_2_wdata_bits_wstrb_1 = dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@148204.4]
  assign io_dram_2_wdata_bits_wstrb_2 = dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@148205.4]
  assign io_dram_2_wdata_bits_wstrb_3 = dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@148206.4]
  assign io_dram_2_wdata_bits_wstrb_4 = dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@148207.4]
  assign io_dram_2_wdata_bits_wstrb_5 = dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@148208.4]
  assign io_dram_2_wdata_bits_wstrb_6 = dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@148209.4]
  assign io_dram_2_wdata_bits_wstrb_7 = dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@148210.4]
  assign io_dram_2_wdata_bits_wstrb_8 = dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@148211.4]
  assign io_dram_2_wdata_bits_wstrb_9 = dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@148212.4]
  assign io_dram_2_wdata_bits_wstrb_10 = dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@148213.4]
  assign io_dram_2_wdata_bits_wstrb_11 = dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@148214.4]
  assign io_dram_2_wdata_bits_wstrb_12 = dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@148215.4]
  assign io_dram_2_wdata_bits_wstrb_13 = dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@148216.4]
  assign io_dram_2_wdata_bits_wstrb_14 = dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@148217.4]
  assign io_dram_2_wdata_bits_wstrb_15 = dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@148218.4]
  assign io_dram_2_wdata_bits_wstrb_16 = dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@148219.4]
  assign io_dram_2_wdata_bits_wstrb_17 = dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@148220.4]
  assign io_dram_2_wdata_bits_wstrb_18 = dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@148221.4]
  assign io_dram_2_wdata_bits_wstrb_19 = dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@148222.4]
  assign io_dram_2_wdata_bits_wstrb_20 = dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@148223.4]
  assign io_dram_2_wdata_bits_wstrb_21 = dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@148224.4]
  assign io_dram_2_wdata_bits_wstrb_22 = dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@148225.4]
  assign io_dram_2_wdata_bits_wstrb_23 = dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@148226.4]
  assign io_dram_2_wdata_bits_wstrb_24 = dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@148227.4]
  assign io_dram_2_wdata_bits_wstrb_25 = dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@148228.4]
  assign io_dram_2_wdata_bits_wstrb_26 = dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@148229.4]
  assign io_dram_2_wdata_bits_wstrb_27 = dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@148230.4]
  assign io_dram_2_wdata_bits_wstrb_28 = dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@148231.4]
  assign io_dram_2_wdata_bits_wstrb_29 = dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@148232.4]
  assign io_dram_2_wdata_bits_wstrb_30 = dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@148233.4]
  assign io_dram_2_wdata_bits_wstrb_31 = dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@148234.4]
  assign io_dram_2_wdata_bits_wstrb_32 = dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@148235.4]
  assign io_dram_2_wdata_bits_wstrb_33 = dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@148236.4]
  assign io_dram_2_wdata_bits_wstrb_34 = dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@148237.4]
  assign io_dram_2_wdata_bits_wstrb_35 = dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@148238.4]
  assign io_dram_2_wdata_bits_wstrb_36 = dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@148239.4]
  assign io_dram_2_wdata_bits_wstrb_37 = dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@148240.4]
  assign io_dram_2_wdata_bits_wstrb_38 = dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@148241.4]
  assign io_dram_2_wdata_bits_wstrb_39 = dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@148242.4]
  assign io_dram_2_wdata_bits_wstrb_40 = dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@148243.4]
  assign io_dram_2_wdata_bits_wstrb_41 = dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@148244.4]
  assign io_dram_2_wdata_bits_wstrb_42 = dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@148245.4]
  assign io_dram_2_wdata_bits_wstrb_43 = dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@148246.4]
  assign io_dram_2_wdata_bits_wstrb_44 = dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@148247.4]
  assign io_dram_2_wdata_bits_wstrb_45 = dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@148248.4]
  assign io_dram_2_wdata_bits_wstrb_46 = dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@148249.4]
  assign io_dram_2_wdata_bits_wstrb_47 = dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@148250.4]
  assign io_dram_2_wdata_bits_wstrb_48 = dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@148251.4]
  assign io_dram_2_wdata_bits_wstrb_49 = dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@148252.4]
  assign io_dram_2_wdata_bits_wstrb_50 = dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@148253.4]
  assign io_dram_2_wdata_bits_wstrb_51 = dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@148254.4]
  assign io_dram_2_wdata_bits_wstrb_52 = dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@148255.4]
  assign io_dram_2_wdata_bits_wstrb_53 = dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@148256.4]
  assign io_dram_2_wdata_bits_wstrb_54 = dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@148257.4]
  assign io_dram_2_wdata_bits_wstrb_55 = dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@148258.4]
  assign io_dram_2_wdata_bits_wstrb_56 = dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@148259.4]
  assign io_dram_2_wdata_bits_wstrb_57 = dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@148260.4]
  assign io_dram_2_wdata_bits_wstrb_58 = dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@148261.4]
  assign io_dram_2_wdata_bits_wstrb_59 = dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@148262.4]
  assign io_dram_2_wdata_bits_wstrb_60 = dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@148263.4]
  assign io_dram_2_wdata_bits_wstrb_61 = dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@148264.4]
  assign io_dram_2_wdata_bits_wstrb_62 = dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@148265.4]
  assign io_dram_2_wdata_bits_wstrb_63 = dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@148266.4]
  assign io_dram_2_wdata_bits_wlast = dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@148202.4]
  assign io_dram_2_rresp_ready = dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 195:72:@148201.4]
  assign io_dram_2_wresp_ready = dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 195:72:@148182.4]
  assign io_dram_3_cmd_valid = dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 195:72:@148402.4]
  assign io_dram_3_cmd_bits_addr = dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@148401.4]
  assign io_dram_3_cmd_bits_size = dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@148400.4]
  assign io_dram_3_cmd_bits_isWr = dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@148398.4]
  assign io_dram_3_cmd_bits_tag = dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@148397.4]
  assign io_dram_3_wdata_valid = dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 195:72:@148395.4]
  assign io_dram_3_wdata_bits_wdata_0 = dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@148379.4]
  assign io_dram_3_wdata_bits_wdata_1 = dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@148380.4]
  assign io_dram_3_wdata_bits_wdata_2 = dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@148381.4]
  assign io_dram_3_wdata_bits_wdata_3 = dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@148382.4]
  assign io_dram_3_wdata_bits_wdata_4 = dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@148383.4]
  assign io_dram_3_wdata_bits_wdata_5 = dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@148384.4]
  assign io_dram_3_wdata_bits_wdata_6 = dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@148385.4]
  assign io_dram_3_wdata_bits_wdata_7 = dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@148386.4]
  assign io_dram_3_wdata_bits_wdata_8 = dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@148387.4]
  assign io_dram_3_wdata_bits_wdata_9 = dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@148388.4]
  assign io_dram_3_wdata_bits_wdata_10 = dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@148389.4]
  assign io_dram_3_wdata_bits_wdata_11 = dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@148390.4]
  assign io_dram_3_wdata_bits_wdata_12 = dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@148391.4]
  assign io_dram_3_wdata_bits_wdata_13 = dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@148392.4]
  assign io_dram_3_wdata_bits_wdata_14 = dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@148393.4]
  assign io_dram_3_wdata_bits_wdata_15 = dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@148394.4]
  assign io_dram_3_wdata_bits_wstrb_0 = dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@148315.4]
  assign io_dram_3_wdata_bits_wstrb_1 = dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@148316.4]
  assign io_dram_3_wdata_bits_wstrb_2 = dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@148317.4]
  assign io_dram_3_wdata_bits_wstrb_3 = dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@148318.4]
  assign io_dram_3_wdata_bits_wstrb_4 = dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@148319.4]
  assign io_dram_3_wdata_bits_wstrb_5 = dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@148320.4]
  assign io_dram_3_wdata_bits_wstrb_6 = dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@148321.4]
  assign io_dram_3_wdata_bits_wstrb_7 = dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@148322.4]
  assign io_dram_3_wdata_bits_wstrb_8 = dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@148323.4]
  assign io_dram_3_wdata_bits_wstrb_9 = dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@148324.4]
  assign io_dram_3_wdata_bits_wstrb_10 = dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@148325.4]
  assign io_dram_3_wdata_bits_wstrb_11 = dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@148326.4]
  assign io_dram_3_wdata_bits_wstrb_12 = dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@148327.4]
  assign io_dram_3_wdata_bits_wstrb_13 = dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@148328.4]
  assign io_dram_3_wdata_bits_wstrb_14 = dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@148329.4]
  assign io_dram_3_wdata_bits_wstrb_15 = dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@148330.4]
  assign io_dram_3_wdata_bits_wstrb_16 = dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@148331.4]
  assign io_dram_3_wdata_bits_wstrb_17 = dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@148332.4]
  assign io_dram_3_wdata_bits_wstrb_18 = dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@148333.4]
  assign io_dram_3_wdata_bits_wstrb_19 = dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@148334.4]
  assign io_dram_3_wdata_bits_wstrb_20 = dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@148335.4]
  assign io_dram_3_wdata_bits_wstrb_21 = dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@148336.4]
  assign io_dram_3_wdata_bits_wstrb_22 = dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@148337.4]
  assign io_dram_3_wdata_bits_wstrb_23 = dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@148338.4]
  assign io_dram_3_wdata_bits_wstrb_24 = dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@148339.4]
  assign io_dram_3_wdata_bits_wstrb_25 = dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@148340.4]
  assign io_dram_3_wdata_bits_wstrb_26 = dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@148341.4]
  assign io_dram_3_wdata_bits_wstrb_27 = dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@148342.4]
  assign io_dram_3_wdata_bits_wstrb_28 = dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@148343.4]
  assign io_dram_3_wdata_bits_wstrb_29 = dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@148344.4]
  assign io_dram_3_wdata_bits_wstrb_30 = dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@148345.4]
  assign io_dram_3_wdata_bits_wstrb_31 = dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@148346.4]
  assign io_dram_3_wdata_bits_wstrb_32 = dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@148347.4]
  assign io_dram_3_wdata_bits_wstrb_33 = dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@148348.4]
  assign io_dram_3_wdata_bits_wstrb_34 = dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@148349.4]
  assign io_dram_3_wdata_bits_wstrb_35 = dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@148350.4]
  assign io_dram_3_wdata_bits_wstrb_36 = dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@148351.4]
  assign io_dram_3_wdata_bits_wstrb_37 = dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@148352.4]
  assign io_dram_3_wdata_bits_wstrb_38 = dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@148353.4]
  assign io_dram_3_wdata_bits_wstrb_39 = dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@148354.4]
  assign io_dram_3_wdata_bits_wstrb_40 = dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@148355.4]
  assign io_dram_3_wdata_bits_wstrb_41 = dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@148356.4]
  assign io_dram_3_wdata_bits_wstrb_42 = dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@148357.4]
  assign io_dram_3_wdata_bits_wstrb_43 = dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@148358.4]
  assign io_dram_3_wdata_bits_wstrb_44 = dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@148359.4]
  assign io_dram_3_wdata_bits_wstrb_45 = dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@148360.4]
  assign io_dram_3_wdata_bits_wstrb_46 = dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@148361.4]
  assign io_dram_3_wdata_bits_wstrb_47 = dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@148362.4]
  assign io_dram_3_wdata_bits_wstrb_48 = dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@148363.4]
  assign io_dram_3_wdata_bits_wstrb_49 = dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@148364.4]
  assign io_dram_3_wdata_bits_wstrb_50 = dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@148365.4]
  assign io_dram_3_wdata_bits_wstrb_51 = dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@148366.4]
  assign io_dram_3_wdata_bits_wstrb_52 = dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@148367.4]
  assign io_dram_3_wdata_bits_wstrb_53 = dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@148368.4]
  assign io_dram_3_wdata_bits_wstrb_54 = dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@148369.4]
  assign io_dram_3_wdata_bits_wstrb_55 = dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@148370.4]
  assign io_dram_3_wdata_bits_wstrb_56 = dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@148371.4]
  assign io_dram_3_wdata_bits_wstrb_57 = dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@148372.4]
  assign io_dram_3_wdata_bits_wstrb_58 = dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@148373.4]
  assign io_dram_3_wdata_bits_wstrb_59 = dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@148374.4]
  assign io_dram_3_wdata_bits_wstrb_60 = dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@148375.4]
  assign io_dram_3_wdata_bits_wstrb_61 = dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@148376.4]
  assign io_dram_3_wdata_bits_wstrb_62 = dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@148377.4]
  assign io_dram_3_wdata_bits_wstrb_63 = dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@148378.4]
  assign io_dram_3_wdata_bits_wlast = dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@148314.4]
  assign io_dram_3_rresp_ready = dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 195:72:@148313.4]
  assign io_dram_3_wresp_ready = dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 195:72:@148294.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@144833.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@144832.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@144831.4]
  assign dramArbs_0_clock = clock; // @[:@140956.4]
  assign dramArbs_0_reset = _T_1030 | reset; // @[:@140957.4 Fringe.scala 187:30:@147948.4]
  assign dramArbs_0_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@147952.4]
  assign dramArbs_0_io_app_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[Fringe.scala 101:72:@141873.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[Fringe.scala 101:72:@141872.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[Fringe.scala 101:72:@141871.4]
  assign dramArbs_0_io_app_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[Fringe.scala 101:72:@141869.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[Fringe.scala 101:72:@141868.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[Fringe.scala 101:72:@141867.4]
  assign dramArbs_0_io_app_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[Fringe.scala 101:72:@141866.4]
  assign dramArbs_0_io_dram_cmd_ready = io_dram_0_cmd_ready; // @[Fringe.scala 195:72:@148067.4]
  assign dramArbs_0_io_dram_wdata_ready = io_dram_0_wdata_ready; // @[Fringe.scala 195:72:@148060.4]
  assign dramArbs_0_io_dram_wresp_valid = io_dram_0_wresp_valid; // @[Fringe.scala 195:72:@147957.4]
  assign dramArbs_0_io_dram_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[Fringe.scala 195:72:@147956.4]
  assign dramArbs_1_clock = clock; // @[:@141949.4]
  assign dramArbs_1_reset = _T_1030 | reset; // @[:@141950.4 Fringe.scala 187:30:@147949.4]
  assign dramArbs_1_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@147953.4]
  assign dramArbs_1_io_dram_cmd_ready = io_dram_1_cmd_ready; // @[Fringe.scala 195:72:@148179.4]
  assign dramArbs_1_io_dram_wdata_ready = io_dram_1_wdata_ready; // @[Fringe.scala 195:72:@148172.4]
  assign dramArbs_1_io_dram_wresp_valid = io_dram_1_wresp_valid; // @[Fringe.scala 195:72:@148069.4]
  assign dramArbs_1_io_dram_wresp_bits_tag = io_dram_1_wresp_bits_tag; // @[Fringe.scala 195:72:@148068.4]
  assign dramArbs_2_clock = clock; // @[:@142909.4]
  assign dramArbs_2_reset = _T_1030 | reset; // @[:@142910.4 Fringe.scala 187:30:@147950.4]
  assign dramArbs_2_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@147954.4]
  assign dramArbs_2_io_dram_cmd_ready = io_dram_2_cmd_ready; // @[Fringe.scala 195:72:@148291.4]
  assign dramArbs_2_io_dram_wdata_ready = io_dram_2_wdata_ready; // @[Fringe.scala 195:72:@148284.4]
  assign dramArbs_2_io_dram_wresp_valid = io_dram_2_wresp_valid; // @[Fringe.scala 195:72:@148181.4]
  assign dramArbs_2_io_dram_wresp_bits_tag = io_dram_2_wresp_bits_tag; // @[Fringe.scala 195:72:@148180.4]
  assign dramArbs_3_clock = clock; // @[:@143869.4]
  assign dramArbs_3_reset = _T_1030 | reset; // @[:@143870.4 Fringe.scala 187:30:@147951.4]
  assign dramArbs_3_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@147955.4]
  assign dramArbs_3_io_dram_cmd_ready = io_dram_3_cmd_ready; // @[Fringe.scala 195:72:@148403.4]
  assign dramArbs_3_io_dram_wdata_ready = io_dram_3_wdata_ready; // @[Fringe.scala 195:72:@148396.4]
  assign dramArbs_3_io_dram_wresp_valid = io_dram_3_wresp_valid; // @[Fringe.scala 195:72:@148293.4]
  assign dramArbs_3_io_dram_wresp_bits_tag = io_dram_3_wresp_bits_tag; // @[Fringe.scala 195:72:@148292.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@144836.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@144835.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@144834.4]
  assign heap_io_host_0_resp_valid = _T_1569 & _T_1573; // @[Fringe.scala 204:22:@148575.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@148576.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@148577.4]
  assign regs_clock = clock; // @[:@144838.4]
  assign regs_reset = reset; // @[:@144839.4 Fringe.scala 139:14:@146886.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@146858.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@146860.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@146859.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@146861.4]
  assign regs_io_reset = _T_1030 | reset; // @[Fringe.scala 138:17:@146884.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_1049; // @[Fringe.scala 170:23:@146936.4]
  assign regs_io_argOuts_0_bits = {_T_1065,_T_1064}; // @[Fringe.scala 171:22:@146940.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@146943.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@146942.4]
  assign timeoutCtr_clock = clock; // @[:@146888.4]
  assign timeoutCtr_reset = reset; // @[:@146889.4]
  assign timeoutCtr_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 149:24:@146903.4]
  assign depulser_clock = clock; // @[:@146907.4]
  assign depulser_reset = reset; // @[:@146908.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@146913.4]
  assign depulser_io_rst = _T_1040[0]; // @[Fringe.scala 156:19:@146915.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1047 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1572 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1047 <= 1'h0;
    end else begin
      _T_1047 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1572 <= 1'h0;
    end else begin
      _T_1572 <= _T_1569;
    end
  end
endmodule
module AXI4LiteToRFBridge( // @[:@148592.2]
  input         clock, // @[:@148593.4]
  input         reset, // @[:@148594.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@148595.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@148595.4]
  input         io_S_AXI_AWVALID, // @[:@148595.4]
  output        io_S_AXI_AWREADY, // @[:@148595.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@148595.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@148595.4]
  input         io_S_AXI_ARVALID, // @[:@148595.4]
  output        io_S_AXI_ARREADY, // @[:@148595.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@148595.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@148595.4]
  input         io_S_AXI_WVALID, // @[:@148595.4]
  output        io_S_AXI_WREADY, // @[:@148595.4]
  output [31:0] io_S_AXI_RDATA, // @[:@148595.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@148595.4]
  output        io_S_AXI_RVALID, // @[:@148595.4]
  input         io_S_AXI_RREADY, // @[:@148595.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@148595.4]
  output        io_S_AXI_BVALID, // @[:@148595.4]
  input         io_S_AXI_BREADY, // @[:@148595.4]
  output [31:0] io_raddr, // @[:@148595.4]
  output        io_wen, // @[:@148595.4]
  output [31:0] io_waddr, // @[:@148595.4]
  output [31:0] io_wdata, // @[:@148595.4]
  input  [31:0] io_rdata // @[:@148595.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 36:17:@148597.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 38:14:@148621.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 38:14:@148617.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 38:14:@148613.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 38:14:@148612.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 38:14:@148611.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 38:14:@148610.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 38:14:@148608.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 38:14:@148607.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 42:12:@148629.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 45:12:@148632.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 43:12:@148630.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 44:12:@148631.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 46:17:@148633.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 40:22:@148628.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 39:19:@148625.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 38:14:@148624.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 38:14:@148623.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 38:14:@148622.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 38:14:@148620.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 38:14:@148619.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 38:14:@148618.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 38:14:@148616.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 38:14:@148615.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 38:14:@148614.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 38:14:@148609.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 38:14:@148606.4]
endmodule
module MAGToAXI4Bridge( // @[:@148635.2]
  output         io_in_cmd_ready, // @[:@148638.4]
  input          io_in_cmd_valid, // @[:@148638.4]
  input  [63:0]  io_in_cmd_bits_addr, // @[:@148638.4]
  input  [31:0]  io_in_cmd_bits_size, // @[:@148638.4]
  input          io_in_cmd_bits_isWr, // @[:@148638.4]
  input  [31:0]  io_in_cmd_bits_tag, // @[:@148638.4]
  output         io_in_wdata_ready, // @[:@148638.4]
  input          io_in_wdata_valid, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_0, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_1, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_2, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_3, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_4, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_5, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_6, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_7, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_8, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_9, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_10, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_11, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_12, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_13, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_14, // @[:@148638.4]
  input  [31:0]  io_in_wdata_bits_wdata_15, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_0, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_1, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_2, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_3, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_4, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_5, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_6, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_7, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_8, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_9, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_10, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_11, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_12, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_13, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_14, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_15, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_16, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_17, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_18, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_19, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_20, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_21, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_22, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_23, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_24, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_25, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_26, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_27, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_28, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_29, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_30, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_31, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_32, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_33, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_34, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_35, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_36, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_37, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_38, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_39, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_40, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_41, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_42, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_43, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_44, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_45, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_46, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_47, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_48, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_49, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_50, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_51, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_52, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_53, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_54, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_55, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_56, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_57, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_58, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_59, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_60, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_61, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_62, // @[:@148638.4]
  input          io_in_wdata_bits_wstrb_63, // @[:@148638.4]
  input          io_in_wdata_bits_wlast, // @[:@148638.4]
  input          io_in_rresp_ready, // @[:@148638.4]
  input          io_in_wresp_ready, // @[:@148638.4]
  output         io_in_wresp_valid, // @[:@148638.4]
  output [31:0]  io_in_wresp_bits_tag, // @[:@148638.4]
  output [31:0]  io_M_AXI_AWID, // @[:@148638.4]
  output [31:0]  io_M_AXI_AWADDR, // @[:@148638.4]
  output [7:0]   io_M_AXI_AWLEN, // @[:@148638.4]
  output         io_M_AXI_AWVALID, // @[:@148638.4]
  input          io_M_AXI_AWREADY, // @[:@148638.4]
  output [31:0]  io_M_AXI_ARID, // @[:@148638.4]
  output [31:0]  io_M_AXI_ARADDR, // @[:@148638.4]
  output [7:0]   io_M_AXI_ARLEN, // @[:@148638.4]
  output         io_M_AXI_ARVALID, // @[:@148638.4]
  input          io_M_AXI_ARREADY, // @[:@148638.4]
  output [511:0] io_M_AXI_WDATA, // @[:@148638.4]
  output [63:0]  io_M_AXI_WSTRB, // @[:@148638.4]
  output         io_M_AXI_WLAST, // @[:@148638.4]
  output         io_M_AXI_WVALID, // @[:@148638.4]
  input          io_M_AXI_WREADY, // @[:@148638.4]
  output         io_M_AXI_RREADY, // @[:@148638.4]
  input  [31:0]  io_M_AXI_BID, // @[:@148638.4]
  input          io_M_AXI_BVALID, // @[:@148638.4]
  output         io_M_AXI_BREADY // @[:@148638.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@148795.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@148796.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@148797.4]
  wire  _T_228; // @[MAGToAXI4Bridge.scala 35:42:@148805.4]
  wire [319:0] _T_250; // @[Cat.scala 30:58:@148832.4]
  wire [479:0] _T_255; // @[Cat.scala 30:58:@148837.4]
  wire [9:0] _T_265; // @[Cat.scala 30:58:@148848.4]
  wire [18:0] _T_274; // @[Cat.scala 30:58:@148857.4]
  wire [27:0] _T_283; // @[Cat.scala 30:58:@148866.4]
  wire [36:0] _T_292; // @[Cat.scala 30:58:@148875.4]
  wire [45:0] _T_301; // @[Cat.scala 30:58:@148884.4]
  wire [54:0] _T_310; // @[Cat.scala 30:58:@148893.4]
  wire [62:0] _T_318; // @[Cat.scala 30:58:@148901.4]
  assign _T_218 = io_in_cmd_bits_size - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@148795.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@148796.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@148797.4]
  assign _T_228 = io_in_cmd_bits_isWr == 1'h0; // @[MAGToAXI4Bridge.scala 35:42:@148805.4]
  assign _T_250 = {io_in_wdata_bits_wdata_15,io_in_wdata_bits_wdata_14,io_in_wdata_bits_wdata_13,io_in_wdata_bits_wdata_12,io_in_wdata_bits_wdata_11,io_in_wdata_bits_wdata_10,io_in_wdata_bits_wdata_9,io_in_wdata_bits_wdata_8,io_in_wdata_bits_wdata_7,io_in_wdata_bits_wdata_6}; // @[Cat.scala 30:58:@148832.4]
  assign _T_255 = {_T_250,io_in_wdata_bits_wdata_5,io_in_wdata_bits_wdata_4,io_in_wdata_bits_wdata_3,io_in_wdata_bits_wdata_2,io_in_wdata_bits_wdata_1}; // @[Cat.scala 30:58:@148837.4]
  assign _T_265 = {io_in_wdata_bits_wstrb_63,io_in_wdata_bits_wstrb_62,io_in_wdata_bits_wstrb_61,io_in_wdata_bits_wstrb_60,io_in_wdata_bits_wstrb_59,io_in_wdata_bits_wstrb_58,io_in_wdata_bits_wstrb_57,io_in_wdata_bits_wstrb_56,io_in_wdata_bits_wstrb_55,io_in_wdata_bits_wstrb_54}; // @[Cat.scala 30:58:@148848.4]
  assign _T_274 = {_T_265,io_in_wdata_bits_wstrb_53,io_in_wdata_bits_wstrb_52,io_in_wdata_bits_wstrb_51,io_in_wdata_bits_wstrb_50,io_in_wdata_bits_wstrb_49,io_in_wdata_bits_wstrb_48,io_in_wdata_bits_wstrb_47,io_in_wdata_bits_wstrb_46,io_in_wdata_bits_wstrb_45}; // @[Cat.scala 30:58:@148857.4]
  assign _T_283 = {_T_274,io_in_wdata_bits_wstrb_44,io_in_wdata_bits_wstrb_43,io_in_wdata_bits_wstrb_42,io_in_wdata_bits_wstrb_41,io_in_wdata_bits_wstrb_40,io_in_wdata_bits_wstrb_39,io_in_wdata_bits_wstrb_38,io_in_wdata_bits_wstrb_37,io_in_wdata_bits_wstrb_36}; // @[Cat.scala 30:58:@148866.4]
  assign _T_292 = {_T_283,io_in_wdata_bits_wstrb_35,io_in_wdata_bits_wstrb_34,io_in_wdata_bits_wstrb_33,io_in_wdata_bits_wstrb_32,io_in_wdata_bits_wstrb_31,io_in_wdata_bits_wstrb_30,io_in_wdata_bits_wstrb_29,io_in_wdata_bits_wstrb_28,io_in_wdata_bits_wstrb_27}; // @[Cat.scala 30:58:@148875.4]
  assign _T_301 = {_T_292,io_in_wdata_bits_wstrb_26,io_in_wdata_bits_wstrb_25,io_in_wdata_bits_wstrb_24,io_in_wdata_bits_wstrb_23,io_in_wdata_bits_wstrb_22,io_in_wdata_bits_wstrb_21,io_in_wdata_bits_wstrb_20,io_in_wdata_bits_wstrb_19,io_in_wdata_bits_wstrb_18}; // @[Cat.scala 30:58:@148884.4]
  assign _T_310 = {_T_301,io_in_wdata_bits_wstrb_17,io_in_wdata_bits_wstrb_16,io_in_wdata_bits_wstrb_15,io_in_wdata_bits_wstrb_14,io_in_wdata_bits_wstrb_13,io_in_wdata_bits_wstrb_12,io_in_wdata_bits_wstrb_11,io_in_wdata_bits_wstrb_10,io_in_wdata_bits_wstrb_9}; // @[Cat.scala 30:58:@148893.4]
  assign _T_318 = {_T_310,io_in_wdata_bits_wstrb_8,io_in_wdata_bits_wstrb_7,io_in_wdata_bits_wstrb_6,io_in_wdata_bits_wstrb_5,io_in_wdata_bits_wstrb_4,io_in_wdata_bits_wstrb_3,io_in_wdata_bits_wstrb_2,io_in_wdata_bits_wstrb_1}; // @[Cat.scala 30:58:@148901.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? io_M_AXI_AWREADY : io_M_AXI_ARREADY; // @[MAGToAXI4Bridge.scala 36:21:@148809.4]
  assign io_in_wdata_ready = io_M_AXI_WREADY; // @[MAGToAXI4Bridge.scala 56:21:@148906.4]
  assign io_in_wresp_valid = io_M_AXI_BVALID; // @[MAGToAXI4Bridge.scala 71:21:@148959.4]
  assign io_in_wresp_bits_tag = io_M_AXI_BID; // @[MAGToAXI4Bridge.scala 74:24:@148961.4]
  assign io_M_AXI_AWID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 39:21:@148810.4]
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 40:21:@148811.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@148815.4]
  assign io_M_AXI_AWVALID = io_in_cmd_valid & io_in_cmd_bits_isWr; // @[MAGToAXI4Bridge.scala 49:21:@148823.4]
  assign io_M_AXI_ARID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 25:21:@148793.4]
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 26:21:@148794.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@148798.4]
  assign io_M_AXI_ARVALID = io_in_cmd_valid & _T_228; // @[MAGToAXI4Bridge.scala 35:21:@148807.4]
  assign io_M_AXI_WDATA = {_T_255,io_in_wdata_bits_wdata_0}; // @[MAGToAXI4Bridge.scala 52:21:@148839.4]
  assign io_M_AXI_WSTRB = {_T_318,io_in_wdata_bits_wstrb_0}; // @[MAGToAXI4Bridge.scala 53:21:@148903.4]
  assign io_M_AXI_WLAST = io_in_wdata_bits_wlast; // @[MAGToAXI4Bridge.scala 54:21:@148904.4]
  assign io_M_AXI_WVALID = io_in_wdata_valid; // @[MAGToAXI4Bridge.scala 55:21:@148905.4]
  assign io_M_AXI_RREADY = io_in_rresp_ready; // @[MAGToAXI4Bridge.scala 64:19:@148956.4]
  assign io_M_AXI_BREADY = io_in_wresp_ready; // @[MAGToAXI4Bridge.scala 67:19:@148957.4]
endmodule
module FringeZynq( // @[:@149947.2]
  input          clock, // @[:@149948.4]
  input          reset, // @[:@149949.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@149950.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@149950.4]
  input          io_S_AXI_AWVALID, // @[:@149950.4]
  output         io_S_AXI_AWREADY, // @[:@149950.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@149950.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@149950.4]
  input          io_S_AXI_ARVALID, // @[:@149950.4]
  output         io_S_AXI_ARREADY, // @[:@149950.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@149950.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@149950.4]
  input          io_S_AXI_WVALID, // @[:@149950.4]
  output         io_S_AXI_WREADY, // @[:@149950.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@149950.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@149950.4]
  output         io_S_AXI_RVALID, // @[:@149950.4]
  input          io_S_AXI_RREADY, // @[:@149950.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@149950.4]
  output         io_S_AXI_BVALID, // @[:@149950.4]
  input          io_S_AXI_BREADY, // @[:@149950.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@149950.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@149950.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@149950.4]
  output         io_M_AXI_0_AWVALID, // @[:@149950.4]
  input          io_M_AXI_0_AWREADY, // @[:@149950.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@149950.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@149950.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@149950.4]
  output         io_M_AXI_0_ARVALID, // @[:@149950.4]
  input          io_M_AXI_0_ARREADY, // @[:@149950.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@149950.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@149950.4]
  output         io_M_AXI_0_WLAST, // @[:@149950.4]
  output         io_M_AXI_0_WVALID, // @[:@149950.4]
  input          io_M_AXI_0_WREADY, // @[:@149950.4]
  output         io_M_AXI_0_RREADY, // @[:@149950.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@149950.4]
  input          io_M_AXI_0_BVALID, // @[:@149950.4]
  output         io_M_AXI_0_BREADY, // @[:@149950.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@149950.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@149950.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@149950.4]
  output         io_M_AXI_1_AWVALID, // @[:@149950.4]
  input          io_M_AXI_1_AWREADY, // @[:@149950.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@149950.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@149950.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@149950.4]
  output         io_M_AXI_1_ARVALID, // @[:@149950.4]
  input          io_M_AXI_1_ARREADY, // @[:@149950.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@149950.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@149950.4]
  output         io_M_AXI_1_WLAST, // @[:@149950.4]
  output         io_M_AXI_1_WVALID, // @[:@149950.4]
  input          io_M_AXI_1_WREADY, // @[:@149950.4]
  output         io_M_AXI_1_RREADY, // @[:@149950.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@149950.4]
  input          io_M_AXI_1_BVALID, // @[:@149950.4]
  output         io_M_AXI_1_BREADY, // @[:@149950.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@149950.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@149950.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@149950.4]
  output         io_M_AXI_2_AWVALID, // @[:@149950.4]
  input          io_M_AXI_2_AWREADY, // @[:@149950.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@149950.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@149950.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@149950.4]
  output         io_M_AXI_2_ARVALID, // @[:@149950.4]
  input          io_M_AXI_2_ARREADY, // @[:@149950.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@149950.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@149950.4]
  output         io_M_AXI_2_WLAST, // @[:@149950.4]
  output         io_M_AXI_2_WVALID, // @[:@149950.4]
  input          io_M_AXI_2_WREADY, // @[:@149950.4]
  output         io_M_AXI_2_RREADY, // @[:@149950.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@149950.4]
  input          io_M_AXI_2_BVALID, // @[:@149950.4]
  output         io_M_AXI_2_BREADY, // @[:@149950.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@149950.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@149950.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@149950.4]
  output         io_M_AXI_3_AWVALID, // @[:@149950.4]
  input          io_M_AXI_3_AWREADY, // @[:@149950.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@149950.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@149950.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@149950.4]
  output         io_M_AXI_3_ARVALID, // @[:@149950.4]
  input          io_M_AXI_3_ARREADY, // @[:@149950.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@149950.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@149950.4]
  output         io_M_AXI_3_WLAST, // @[:@149950.4]
  output         io_M_AXI_3_WVALID, // @[:@149950.4]
  input          io_M_AXI_3_WREADY, // @[:@149950.4]
  output         io_M_AXI_3_RREADY, // @[:@149950.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@149950.4]
  input          io_M_AXI_3_BVALID, // @[:@149950.4]
  output         io_M_AXI_3_BREADY, // @[:@149950.4]
  output         io_enable, // @[:@149950.4]
  input          io_done, // @[:@149950.4]
  output         io_reset, // @[:@149950.4]
  output [63:0]  io_argIns_0, // @[:@149950.4]
  output [63:0]  io_argIns_1, // @[:@149950.4]
  input          io_argOuts_0_valid, // @[:@149950.4]
  input  [63:0]  io_argOuts_0_bits, // @[:@149950.4]
  output         io_memStreams_stores_0_cmd_ready, // @[:@149950.4]
  input          io_memStreams_stores_0_cmd_valid, // @[:@149950.4]
  input  [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@149950.4]
  input  [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@149950.4]
  output         io_memStreams_stores_0_data_ready, // @[:@149950.4]
  input          io_memStreams_stores_0_data_valid, // @[:@149950.4]
  input  [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@149950.4]
  input          io_memStreams_stores_0_data_bits_wstrb, // @[:@149950.4]
  input          io_memStreams_stores_0_wresp_ready, // @[:@149950.4]
  output         io_memStreams_stores_0_wresp_valid, // @[:@149950.4]
  output         io_memStreams_stores_0_wresp_bits, // @[:@149950.4]
  input          io_heap_0_req_valid, // @[:@149950.4]
  input          io_heap_0_req_bits_allocDealloc, // @[:@149950.4]
  input  [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@149950.4]
  output         io_heap_0_resp_valid, // @[:@149950.4]
  output         io_heap_0_resp_bits_allocDealloc, // @[:@149950.4]
  output [63:0]  io_heap_0_resp_bits_sizeAddr // @[:@149950.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 69:28:@150421.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 69:28:@150421.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 69:28:@150421.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 69:28:@150421.4]
  wire [63:0] fringeCommon_io_argIns_1; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire [63:0] fringeCommon_io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_cmd_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_0_wresp_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_0_wresp_bits_tag; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_cmd_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire [63:0] fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_1_wresp_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_1_wresp_bits_tag; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_cmd_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire [63:0] fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_2_wresp_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_2_wresp_bits_tag; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_cmd_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire [63:0] fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_dram_3_wresp_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire [31:0] fringeCommon_io_dram_3_wresp_bits_tag; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 69:28:@150421.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 69:28:@150421.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 69:28:@150421.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 69:28:@150421.4]
  wire  AXI4LiteToRFBridge_clock; // @[FringeZynq.scala 90:31:@151327.4]
  wire  AXI4LiteToRFBridge_reset; // @[FringeZynq.scala 90:31:@151327.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_AWADDR; // @[FringeZynq.scala 90:31:@151327.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_AWPROT; // @[FringeZynq.scala 90:31:@151327.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWVALID; // @[FringeZynq.scala 90:31:@151327.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 90:31:@151327.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_ARADDR; // @[FringeZynq.scala 90:31:@151327.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_ARPROT; // @[FringeZynq.scala 90:31:@151327.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARVALID; // @[FringeZynq.scala 90:31:@151327.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 90:31:@151327.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_WDATA; // @[FringeZynq.scala 90:31:@151327.4]
  wire [3:0] AXI4LiteToRFBridge_io_S_AXI_WSTRB; // @[FringeZynq.scala 90:31:@151327.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WVALID; // @[FringeZynq.scala 90:31:@151327.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 90:31:@151327.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 90:31:@151327.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 90:31:@151327.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 90:31:@151327.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RREADY; // @[FringeZynq.scala 90:31:@151327.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 90:31:@151327.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 90:31:@151327.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BREADY; // @[FringeZynq.scala 90:31:@151327.4]
  wire [31:0] AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 90:31:@151327.4]
  wire  AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 90:31:@151327.4]
  wire [31:0] AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 90:31:@151327.4]
  wire [31:0] AXI4LiteToRFBridge_io_wdata; // @[FringeZynq.scala 90:31:@151327.4]
  wire [31:0] AXI4LiteToRFBridge_io_rdata; // @[FringeZynq.scala 90:31:@151327.4]
  wire  MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@151477.4]
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@151477.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@151477.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@151477.4]
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@151477.4]
  wire [63:0] MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@151477.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@151477.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@151633.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@151633.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@151633.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@151633.4]
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@151633.4]
  wire [63:0] MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@151633.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@151633.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@151789.4]
  wire [63:0] MAGToAXI4Bridge_2_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@151789.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@151789.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@151789.4]
  wire [511:0] MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@151789.4]
  wire [63:0] MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@151789.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@151789.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@151945.4]
  wire [63:0] MAGToAXI4Bridge_3_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@151945.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@151945.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@151945.4]
  wire [511:0] MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@151945.4]
  wire [63:0] MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@151945.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@151945.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@151945.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 69:28:@150421.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argIns_1(fringeCommon_io_argIns_1),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(fringeCommon_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(fringeCommon_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(fringeCommon_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(fringeCommon_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(fringeCommon_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(fringeCommon_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(fringeCommon_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(fringeCommon_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(fringeCommon_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(fringeCommon_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(fringeCommon_io_memStreams_stores_0_wresp_bits),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_isWr(fringeCommon_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag(fringeCommon_io_dram_0_cmd_bits_tag),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(fringeCommon_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(fringeCommon_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(fringeCommon_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(fringeCommon_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(fringeCommon_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(fringeCommon_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(fringeCommon_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(fringeCommon_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(fringeCommon_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wdata_8(fringeCommon_io_dram_0_wdata_bits_wdata_8),
    .io_dram_0_wdata_bits_wdata_9(fringeCommon_io_dram_0_wdata_bits_wdata_9),
    .io_dram_0_wdata_bits_wdata_10(fringeCommon_io_dram_0_wdata_bits_wdata_10),
    .io_dram_0_wdata_bits_wdata_11(fringeCommon_io_dram_0_wdata_bits_wdata_11),
    .io_dram_0_wdata_bits_wdata_12(fringeCommon_io_dram_0_wdata_bits_wdata_12),
    .io_dram_0_wdata_bits_wdata_13(fringeCommon_io_dram_0_wdata_bits_wdata_13),
    .io_dram_0_wdata_bits_wdata_14(fringeCommon_io_dram_0_wdata_bits_wdata_14),
    .io_dram_0_wdata_bits_wdata_15(fringeCommon_io_dram_0_wdata_bits_wdata_15),
    .io_dram_0_wdata_bits_wstrb_0(fringeCommon_io_dram_0_wdata_bits_wstrb_0),
    .io_dram_0_wdata_bits_wstrb_1(fringeCommon_io_dram_0_wdata_bits_wstrb_1),
    .io_dram_0_wdata_bits_wstrb_2(fringeCommon_io_dram_0_wdata_bits_wstrb_2),
    .io_dram_0_wdata_bits_wstrb_3(fringeCommon_io_dram_0_wdata_bits_wstrb_3),
    .io_dram_0_wdata_bits_wstrb_4(fringeCommon_io_dram_0_wdata_bits_wstrb_4),
    .io_dram_0_wdata_bits_wstrb_5(fringeCommon_io_dram_0_wdata_bits_wstrb_5),
    .io_dram_0_wdata_bits_wstrb_6(fringeCommon_io_dram_0_wdata_bits_wstrb_6),
    .io_dram_0_wdata_bits_wstrb_7(fringeCommon_io_dram_0_wdata_bits_wstrb_7),
    .io_dram_0_wdata_bits_wstrb_8(fringeCommon_io_dram_0_wdata_bits_wstrb_8),
    .io_dram_0_wdata_bits_wstrb_9(fringeCommon_io_dram_0_wdata_bits_wstrb_9),
    .io_dram_0_wdata_bits_wstrb_10(fringeCommon_io_dram_0_wdata_bits_wstrb_10),
    .io_dram_0_wdata_bits_wstrb_11(fringeCommon_io_dram_0_wdata_bits_wstrb_11),
    .io_dram_0_wdata_bits_wstrb_12(fringeCommon_io_dram_0_wdata_bits_wstrb_12),
    .io_dram_0_wdata_bits_wstrb_13(fringeCommon_io_dram_0_wdata_bits_wstrb_13),
    .io_dram_0_wdata_bits_wstrb_14(fringeCommon_io_dram_0_wdata_bits_wstrb_14),
    .io_dram_0_wdata_bits_wstrb_15(fringeCommon_io_dram_0_wdata_bits_wstrb_15),
    .io_dram_0_wdata_bits_wstrb_16(fringeCommon_io_dram_0_wdata_bits_wstrb_16),
    .io_dram_0_wdata_bits_wstrb_17(fringeCommon_io_dram_0_wdata_bits_wstrb_17),
    .io_dram_0_wdata_bits_wstrb_18(fringeCommon_io_dram_0_wdata_bits_wstrb_18),
    .io_dram_0_wdata_bits_wstrb_19(fringeCommon_io_dram_0_wdata_bits_wstrb_19),
    .io_dram_0_wdata_bits_wstrb_20(fringeCommon_io_dram_0_wdata_bits_wstrb_20),
    .io_dram_0_wdata_bits_wstrb_21(fringeCommon_io_dram_0_wdata_bits_wstrb_21),
    .io_dram_0_wdata_bits_wstrb_22(fringeCommon_io_dram_0_wdata_bits_wstrb_22),
    .io_dram_0_wdata_bits_wstrb_23(fringeCommon_io_dram_0_wdata_bits_wstrb_23),
    .io_dram_0_wdata_bits_wstrb_24(fringeCommon_io_dram_0_wdata_bits_wstrb_24),
    .io_dram_0_wdata_bits_wstrb_25(fringeCommon_io_dram_0_wdata_bits_wstrb_25),
    .io_dram_0_wdata_bits_wstrb_26(fringeCommon_io_dram_0_wdata_bits_wstrb_26),
    .io_dram_0_wdata_bits_wstrb_27(fringeCommon_io_dram_0_wdata_bits_wstrb_27),
    .io_dram_0_wdata_bits_wstrb_28(fringeCommon_io_dram_0_wdata_bits_wstrb_28),
    .io_dram_0_wdata_bits_wstrb_29(fringeCommon_io_dram_0_wdata_bits_wstrb_29),
    .io_dram_0_wdata_bits_wstrb_30(fringeCommon_io_dram_0_wdata_bits_wstrb_30),
    .io_dram_0_wdata_bits_wstrb_31(fringeCommon_io_dram_0_wdata_bits_wstrb_31),
    .io_dram_0_wdata_bits_wstrb_32(fringeCommon_io_dram_0_wdata_bits_wstrb_32),
    .io_dram_0_wdata_bits_wstrb_33(fringeCommon_io_dram_0_wdata_bits_wstrb_33),
    .io_dram_0_wdata_bits_wstrb_34(fringeCommon_io_dram_0_wdata_bits_wstrb_34),
    .io_dram_0_wdata_bits_wstrb_35(fringeCommon_io_dram_0_wdata_bits_wstrb_35),
    .io_dram_0_wdata_bits_wstrb_36(fringeCommon_io_dram_0_wdata_bits_wstrb_36),
    .io_dram_0_wdata_bits_wstrb_37(fringeCommon_io_dram_0_wdata_bits_wstrb_37),
    .io_dram_0_wdata_bits_wstrb_38(fringeCommon_io_dram_0_wdata_bits_wstrb_38),
    .io_dram_0_wdata_bits_wstrb_39(fringeCommon_io_dram_0_wdata_bits_wstrb_39),
    .io_dram_0_wdata_bits_wstrb_40(fringeCommon_io_dram_0_wdata_bits_wstrb_40),
    .io_dram_0_wdata_bits_wstrb_41(fringeCommon_io_dram_0_wdata_bits_wstrb_41),
    .io_dram_0_wdata_bits_wstrb_42(fringeCommon_io_dram_0_wdata_bits_wstrb_42),
    .io_dram_0_wdata_bits_wstrb_43(fringeCommon_io_dram_0_wdata_bits_wstrb_43),
    .io_dram_0_wdata_bits_wstrb_44(fringeCommon_io_dram_0_wdata_bits_wstrb_44),
    .io_dram_0_wdata_bits_wstrb_45(fringeCommon_io_dram_0_wdata_bits_wstrb_45),
    .io_dram_0_wdata_bits_wstrb_46(fringeCommon_io_dram_0_wdata_bits_wstrb_46),
    .io_dram_0_wdata_bits_wstrb_47(fringeCommon_io_dram_0_wdata_bits_wstrb_47),
    .io_dram_0_wdata_bits_wstrb_48(fringeCommon_io_dram_0_wdata_bits_wstrb_48),
    .io_dram_0_wdata_bits_wstrb_49(fringeCommon_io_dram_0_wdata_bits_wstrb_49),
    .io_dram_0_wdata_bits_wstrb_50(fringeCommon_io_dram_0_wdata_bits_wstrb_50),
    .io_dram_0_wdata_bits_wstrb_51(fringeCommon_io_dram_0_wdata_bits_wstrb_51),
    .io_dram_0_wdata_bits_wstrb_52(fringeCommon_io_dram_0_wdata_bits_wstrb_52),
    .io_dram_0_wdata_bits_wstrb_53(fringeCommon_io_dram_0_wdata_bits_wstrb_53),
    .io_dram_0_wdata_bits_wstrb_54(fringeCommon_io_dram_0_wdata_bits_wstrb_54),
    .io_dram_0_wdata_bits_wstrb_55(fringeCommon_io_dram_0_wdata_bits_wstrb_55),
    .io_dram_0_wdata_bits_wstrb_56(fringeCommon_io_dram_0_wdata_bits_wstrb_56),
    .io_dram_0_wdata_bits_wstrb_57(fringeCommon_io_dram_0_wdata_bits_wstrb_57),
    .io_dram_0_wdata_bits_wstrb_58(fringeCommon_io_dram_0_wdata_bits_wstrb_58),
    .io_dram_0_wdata_bits_wstrb_59(fringeCommon_io_dram_0_wdata_bits_wstrb_59),
    .io_dram_0_wdata_bits_wstrb_60(fringeCommon_io_dram_0_wdata_bits_wstrb_60),
    .io_dram_0_wdata_bits_wstrb_61(fringeCommon_io_dram_0_wdata_bits_wstrb_61),
    .io_dram_0_wdata_bits_wstrb_62(fringeCommon_io_dram_0_wdata_bits_wstrb_62),
    .io_dram_0_wdata_bits_wstrb_63(fringeCommon_io_dram_0_wdata_bits_wstrb_63),
    .io_dram_0_wdata_bits_wlast(fringeCommon_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag(fringeCommon_io_dram_0_wresp_bits_tag),
    .io_dram_1_cmd_ready(fringeCommon_io_dram_1_cmd_ready),
    .io_dram_1_cmd_valid(fringeCommon_io_dram_1_cmd_valid),
    .io_dram_1_cmd_bits_addr(fringeCommon_io_dram_1_cmd_bits_addr),
    .io_dram_1_cmd_bits_size(fringeCommon_io_dram_1_cmd_bits_size),
    .io_dram_1_cmd_bits_isWr(fringeCommon_io_dram_1_cmd_bits_isWr),
    .io_dram_1_cmd_bits_tag(fringeCommon_io_dram_1_cmd_bits_tag),
    .io_dram_1_wdata_ready(fringeCommon_io_dram_1_wdata_ready),
    .io_dram_1_wdata_valid(fringeCommon_io_dram_1_wdata_valid),
    .io_dram_1_wdata_bits_wdata_0(fringeCommon_io_dram_1_wdata_bits_wdata_0),
    .io_dram_1_wdata_bits_wdata_1(fringeCommon_io_dram_1_wdata_bits_wdata_1),
    .io_dram_1_wdata_bits_wdata_2(fringeCommon_io_dram_1_wdata_bits_wdata_2),
    .io_dram_1_wdata_bits_wdata_3(fringeCommon_io_dram_1_wdata_bits_wdata_3),
    .io_dram_1_wdata_bits_wdata_4(fringeCommon_io_dram_1_wdata_bits_wdata_4),
    .io_dram_1_wdata_bits_wdata_5(fringeCommon_io_dram_1_wdata_bits_wdata_5),
    .io_dram_1_wdata_bits_wdata_6(fringeCommon_io_dram_1_wdata_bits_wdata_6),
    .io_dram_1_wdata_bits_wdata_7(fringeCommon_io_dram_1_wdata_bits_wdata_7),
    .io_dram_1_wdata_bits_wdata_8(fringeCommon_io_dram_1_wdata_bits_wdata_8),
    .io_dram_1_wdata_bits_wdata_9(fringeCommon_io_dram_1_wdata_bits_wdata_9),
    .io_dram_1_wdata_bits_wdata_10(fringeCommon_io_dram_1_wdata_bits_wdata_10),
    .io_dram_1_wdata_bits_wdata_11(fringeCommon_io_dram_1_wdata_bits_wdata_11),
    .io_dram_1_wdata_bits_wdata_12(fringeCommon_io_dram_1_wdata_bits_wdata_12),
    .io_dram_1_wdata_bits_wdata_13(fringeCommon_io_dram_1_wdata_bits_wdata_13),
    .io_dram_1_wdata_bits_wdata_14(fringeCommon_io_dram_1_wdata_bits_wdata_14),
    .io_dram_1_wdata_bits_wdata_15(fringeCommon_io_dram_1_wdata_bits_wdata_15),
    .io_dram_1_wdata_bits_wstrb_0(fringeCommon_io_dram_1_wdata_bits_wstrb_0),
    .io_dram_1_wdata_bits_wstrb_1(fringeCommon_io_dram_1_wdata_bits_wstrb_1),
    .io_dram_1_wdata_bits_wstrb_2(fringeCommon_io_dram_1_wdata_bits_wstrb_2),
    .io_dram_1_wdata_bits_wstrb_3(fringeCommon_io_dram_1_wdata_bits_wstrb_3),
    .io_dram_1_wdata_bits_wstrb_4(fringeCommon_io_dram_1_wdata_bits_wstrb_4),
    .io_dram_1_wdata_bits_wstrb_5(fringeCommon_io_dram_1_wdata_bits_wstrb_5),
    .io_dram_1_wdata_bits_wstrb_6(fringeCommon_io_dram_1_wdata_bits_wstrb_6),
    .io_dram_1_wdata_bits_wstrb_7(fringeCommon_io_dram_1_wdata_bits_wstrb_7),
    .io_dram_1_wdata_bits_wstrb_8(fringeCommon_io_dram_1_wdata_bits_wstrb_8),
    .io_dram_1_wdata_bits_wstrb_9(fringeCommon_io_dram_1_wdata_bits_wstrb_9),
    .io_dram_1_wdata_bits_wstrb_10(fringeCommon_io_dram_1_wdata_bits_wstrb_10),
    .io_dram_1_wdata_bits_wstrb_11(fringeCommon_io_dram_1_wdata_bits_wstrb_11),
    .io_dram_1_wdata_bits_wstrb_12(fringeCommon_io_dram_1_wdata_bits_wstrb_12),
    .io_dram_1_wdata_bits_wstrb_13(fringeCommon_io_dram_1_wdata_bits_wstrb_13),
    .io_dram_1_wdata_bits_wstrb_14(fringeCommon_io_dram_1_wdata_bits_wstrb_14),
    .io_dram_1_wdata_bits_wstrb_15(fringeCommon_io_dram_1_wdata_bits_wstrb_15),
    .io_dram_1_wdata_bits_wstrb_16(fringeCommon_io_dram_1_wdata_bits_wstrb_16),
    .io_dram_1_wdata_bits_wstrb_17(fringeCommon_io_dram_1_wdata_bits_wstrb_17),
    .io_dram_1_wdata_bits_wstrb_18(fringeCommon_io_dram_1_wdata_bits_wstrb_18),
    .io_dram_1_wdata_bits_wstrb_19(fringeCommon_io_dram_1_wdata_bits_wstrb_19),
    .io_dram_1_wdata_bits_wstrb_20(fringeCommon_io_dram_1_wdata_bits_wstrb_20),
    .io_dram_1_wdata_bits_wstrb_21(fringeCommon_io_dram_1_wdata_bits_wstrb_21),
    .io_dram_1_wdata_bits_wstrb_22(fringeCommon_io_dram_1_wdata_bits_wstrb_22),
    .io_dram_1_wdata_bits_wstrb_23(fringeCommon_io_dram_1_wdata_bits_wstrb_23),
    .io_dram_1_wdata_bits_wstrb_24(fringeCommon_io_dram_1_wdata_bits_wstrb_24),
    .io_dram_1_wdata_bits_wstrb_25(fringeCommon_io_dram_1_wdata_bits_wstrb_25),
    .io_dram_1_wdata_bits_wstrb_26(fringeCommon_io_dram_1_wdata_bits_wstrb_26),
    .io_dram_1_wdata_bits_wstrb_27(fringeCommon_io_dram_1_wdata_bits_wstrb_27),
    .io_dram_1_wdata_bits_wstrb_28(fringeCommon_io_dram_1_wdata_bits_wstrb_28),
    .io_dram_1_wdata_bits_wstrb_29(fringeCommon_io_dram_1_wdata_bits_wstrb_29),
    .io_dram_1_wdata_bits_wstrb_30(fringeCommon_io_dram_1_wdata_bits_wstrb_30),
    .io_dram_1_wdata_bits_wstrb_31(fringeCommon_io_dram_1_wdata_bits_wstrb_31),
    .io_dram_1_wdata_bits_wstrb_32(fringeCommon_io_dram_1_wdata_bits_wstrb_32),
    .io_dram_1_wdata_bits_wstrb_33(fringeCommon_io_dram_1_wdata_bits_wstrb_33),
    .io_dram_1_wdata_bits_wstrb_34(fringeCommon_io_dram_1_wdata_bits_wstrb_34),
    .io_dram_1_wdata_bits_wstrb_35(fringeCommon_io_dram_1_wdata_bits_wstrb_35),
    .io_dram_1_wdata_bits_wstrb_36(fringeCommon_io_dram_1_wdata_bits_wstrb_36),
    .io_dram_1_wdata_bits_wstrb_37(fringeCommon_io_dram_1_wdata_bits_wstrb_37),
    .io_dram_1_wdata_bits_wstrb_38(fringeCommon_io_dram_1_wdata_bits_wstrb_38),
    .io_dram_1_wdata_bits_wstrb_39(fringeCommon_io_dram_1_wdata_bits_wstrb_39),
    .io_dram_1_wdata_bits_wstrb_40(fringeCommon_io_dram_1_wdata_bits_wstrb_40),
    .io_dram_1_wdata_bits_wstrb_41(fringeCommon_io_dram_1_wdata_bits_wstrb_41),
    .io_dram_1_wdata_bits_wstrb_42(fringeCommon_io_dram_1_wdata_bits_wstrb_42),
    .io_dram_1_wdata_bits_wstrb_43(fringeCommon_io_dram_1_wdata_bits_wstrb_43),
    .io_dram_1_wdata_bits_wstrb_44(fringeCommon_io_dram_1_wdata_bits_wstrb_44),
    .io_dram_1_wdata_bits_wstrb_45(fringeCommon_io_dram_1_wdata_bits_wstrb_45),
    .io_dram_1_wdata_bits_wstrb_46(fringeCommon_io_dram_1_wdata_bits_wstrb_46),
    .io_dram_1_wdata_bits_wstrb_47(fringeCommon_io_dram_1_wdata_bits_wstrb_47),
    .io_dram_1_wdata_bits_wstrb_48(fringeCommon_io_dram_1_wdata_bits_wstrb_48),
    .io_dram_1_wdata_bits_wstrb_49(fringeCommon_io_dram_1_wdata_bits_wstrb_49),
    .io_dram_1_wdata_bits_wstrb_50(fringeCommon_io_dram_1_wdata_bits_wstrb_50),
    .io_dram_1_wdata_bits_wstrb_51(fringeCommon_io_dram_1_wdata_bits_wstrb_51),
    .io_dram_1_wdata_bits_wstrb_52(fringeCommon_io_dram_1_wdata_bits_wstrb_52),
    .io_dram_1_wdata_bits_wstrb_53(fringeCommon_io_dram_1_wdata_bits_wstrb_53),
    .io_dram_1_wdata_bits_wstrb_54(fringeCommon_io_dram_1_wdata_bits_wstrb_54),
    .io_dram_1_wdata_bits_wstrb_55(fringeCommon_io_dram_1_wdata_bits_wstrb_55),
    .io_dram_1_wdata_bits_wstrb_56(fringeCommon_io_dram_1_wdata_bits_wstrb_56),
    .io_dram_1_wdata_bits_wstrb_57(fringeCommon_io_dram_1_wdata_bits_wstrb_57),
    .io_dram_1_wdata_bits_wstrb_58(fringeCommon_io_dram_1_wdata_bits_wstrb_58),
    .io_dram_1_wdata_bits_wstrb_59(fringeCommon_io_dram_1_wdata_bits_wstrb_59),
    .io_dram_1_wdata_bits_wstrb_60(fringeCommon_io_dram_1_wdata_bits_wstrb_60),
    .io_dram_1_wdata_bits_wstrb_61(fringeCommon_io_dram_1_wdata_bits_wstrb_61),
    .io_dram_1_wdata_bits_wstrb_62(fringeCommon_io_dram_1_wdata_bits_wstrb_62),
    .io_dram_1_wdata_bits_wstrb_63(fringeCommon_io_dram_1_wdata_bits_wstrb_63),
    .io_dram_1_wdata_bits_wlast(fringeCommon_io_dram_1_wdata_bits_wlast),
    .io_dram_1_rresp_ready(fringeCommon_io_dram_1_rresp_ready),
    .io_dram_1_wresp_ready(fringeCommon_io_dram_1_wresp_ready),
    .io_dram_1_wresp_valid(fringeCommon_io_dram_1_wresp_valid),
    .io_dram_1_wresp_bits_tag(fringeCommon_io_dram_1_wresp_bits_tag),
    .io_dram_2_cmd_ready(fringeCommon_io_dram_2_cmd_ready),
    .io_dram_2_cmd_valid(fringeCommon_io_dram_2_cmd_valid),
    .io_dram_2_cmd_bits_addr(fringeCommon_io_dram_2_cmd_bits_addr),
    .io_dram_2_cmd_bits_size(fringeCommon_io_dram_2_cmd_bits_size),
    .io_dram_2_cmd_bits_isWr(fringeCommon_io_dram_2_cmd_bits_isWr),
    .io_dram_2_cmd_bits_tag(fringeCommon_io_dram_2_cmd_bits_tag),
    .io_dram_2_wdata_ready(fringeCommon_io_dram_2_wdata_ready),
    .io_dram_2_wdata_valid(fringeCommon_io_dram_2_wdata_valid),
    .io_dram_2_wdata_bits_wdata_0(fringeCommon_io_dram_2_wdata_bits_wdata_0),
    .io_dram_2_wdata_bits_wdata_1(fringeCommon_io_dram_2_wdata_bits_wdata_1),
    .io_dram_2_wdata_bits_wdata_2(fringeCommon_io_dram_2_wdata_bits_wdata_2),
    .io_dram_2_wdata_bits_wdata_3(fringeCommon_io_dram_2_wdata_bits_wdata_3),
    .io_dram_2_wdata_bits_wdata_4(fringeCommon_io_dram_2_wdata_bits_wdata_4),
    .io_dram_2_wdata_bits_wdata_5(fringeCommon_io_dram_2_wdata_bits_wdata_5),
    .io_dram_2_wdata_bits_wdata_6(fringeCommon_io_dram_2_wdata_bits_wdata_6),
    .io_dram_2_wdata_bits_wdata_7(fringeCommon_io_dram_2_wdata_bits_wdata_7),
    .io_dram_2_wdata_bits_wdata_8(fringeCommon_io_dram_2_wdata_bits_wdata_8),
    .io_dram_2_wdata_bits_wdata_9(fringeCommon_io_dram_2_wdata_bits_wdata_9),
    .io_dram_2_wdata_bits_wdata_10(fringeCommon_io_dram_2_wdata_bits_wdata_10),
    .io_dram_2_wdata_bits_wdata_11(fringeCommon_io_dram_2_wdata_bits_wdata_11),
    .io_dram_2_wdata_bits_wdata_12(fringeCommon_io_dram_2_wdata_bits_wdata_12),
    .io_dram_2_wdata_bits_wdata_13(fringeCommon_io_dram_2_wdata_bits_wdata_13),
    .io_dram_2_wdata_bits_wdata_14(fringeCommon_io_dram_2_wdata_bits_wdata_14),
    .io_dram_2_wdata_bits_wdata_15(fringeCommon_io_dram_2_wdata_bits_wdata_15),
    .io_dram_2_wdata_bits_wstrb_0(fringeCommon_io_dram_2_wdata_bits_wstrb_0),
    .io_dram_2_wdata_bits_wstrb_1(fringeCommon_io_dram_2_wdata_bits_wstrb_1),
    .io_dram_2_wdata_bits_wstrb_2(fringeCommon_io_dram_2_wdata_bits_wstrb_2),
    .io_dram_2_wdata_bits_wstrb_3(fringeCommon_io_dram_2_wdata_bits_wstrb_3),
    .io_dram_2_wdata_bits_wstrb_4(fringeCommon_io_dram_2_wdata_bits_wstrb_4),
    .io_dram_2_wdata_bits_wstrb_5(fringeCommon_io_dram_2_wdata_bits_wstrb_5),
    .io_dram_2_wdata_bits_wstrb_6(fringeCommon_io_dram_2_wdata_bits_wstrb_6),
    .io_dram_2_wdata_bits_wstrb_7(fringeCommon_io_dram_2_wdata_bits_wstrb_7),
    .io_dram_2_wdata_bits_wstrb_8(fringeCommon_io_dram_2_wdata_bits_wstrb_8),
    .io_dram_2_wdata_bits_wstrb_9(fringeCommon_io_dram_2_wdata_bits_wstrb_9),
    .io_dram_2_wdata_bits_wstrb_10(fringeCommon_io_dram_2_wdata_bits_wstrb_10),
    .io_dram_2_wdata_bits_wstrb_11(fringeCommon_io_dram_2_wdata_bits_wstrb_11),
    .io_dram_2_wdata_bits_wstrb_12(fringeCommon_io_dram_2_wdata_bits_wstrb_12),
    .io_dram_2_wdata_bits_wstrb_13(fringeCommon_io_dram_2_wdata_bits_wstrb_13),
    .io_dram_2_wdata_bits_wstrb_14(fringeCommon_io_dram_2_wdata_bits_wstrb_14),
    .io_dram_2_wdata_bits_wstrb_15(fringeCommon_io_dram_2_wdata_bits_wstrb_15),
    .io_dram_2_wdata_bits_wstrb_16(fringeCommon_io_dram_2_wdata_bits_wstrb_16),
    .io_dram_2_wdata_bits_wstrb_17(fringeCommon_io_dram_2_wdata_bits_wstrb_17),
    .io_dram_2_wdata_bits_wstrb_18(fringeCommon_io_dram_2_wdata_bits_wstrb_18),
    .io_dram_2_wdata_bits_wstrb_19(fringeCommon_io_dram_2_wdata_bits_wstrb_19),
    .io_dram_2_wdata_bits_wstrb_20(fringeCommon_io_dram_2_wdata_bits_wstrb_20),
    .io_dram_2_wdata_bits_wstrb_21(fringeCommon_io_dram_2_wdata_bits_wstrb_21),
    .io_dram_2_wdata_bits_wstrb_22(fringeCommon_io_dram_2_wdata_bits_wstrb_22),
    .io_dram_2_wdata_bits_wstrb_23(fringeCommon_io_dram_2_wdata_bits_wstrb_23),
    .io_dram_2_wdata_bits_wstrb_24(fringeCommon_io_dram_2_wdata_bits_wstrb_24),
    .io_dram_2_wdata_bits_wstrb_25(fringeCommon_io_dram_2_wdata_bits_wstrb_25),
    .io_dram_2_wdata_bits_wstrb_26(fringeCommon_io_dram_2_wdata_bits_wstrb_26),
    .io_dram_2_wdata_bits_wstrb_27(fringeCommon_io_dram_2_wdata_bits_wstrb_27),
    .io_dram_2_wdata_bits_wstrb_28(fringeCommon_io_dram_2_wdata_bits_wstrb_28),
    .io_dram_2_wdata_bits_wstrb_29(fringeCommon_io_dram_2_wdata_bits_wstrb_29),
    .io_dram_2_wdata_bits_wstrb_30(fringeCommon_io_dram_2_wdata_bits_wstrb_30),
    .io_dram_2_wdata_bits_wstrb_31(fringeCommon_io_dram_2_wdata_bits_wstrb_31),
    .io_dram_2_wdata_bits_wstrb_32(fringeCommon_io_dram_2_wdata_bits_wstrb_32),
    .io_dram_2_wdata_bits_wstrb_33(fringeCommon_io_dram_2_wdata_bits_wstrb_33),
    .io_dram_2_wdata_bits_wstrb_34(fringeCommon_io_dram_2_wdata_bits_wstrb_34),
    .io_dram_2_wdata_bits_wstrb_35(fringeCommon_io_dram_2_wdata_bits_wstrb_35),
    .io_dram_2_wdata_bits_wstrb_36(fringeCommon_io_dram_2_wdata_bits_wstrb_36),
    .io_dram_2_wdata_bits_wstrb_37(fringeCommon_io_dram_2_wdata_bits_wstrb_37),
    .io_dram_2_wdata_bits_wstrb_38(fringeCommon_io_dram_2_wdata_bits_wstrb_38),
    .io_dram_2_wdata_bits_wstrb_39(fringeCommon_io_dram_2_wdata_bits_wstrb_39),
    .io_dram_2_wdata_bits_wstrb_40(fringeCommon_io_dram_2_wdata_bits_wstrb_40),
    .io_dram_2_wdata_bits_wstrb_41(fringeCommon_io_dram_2_wdata_bits_wstrb_41),
    .io_dram_2_wdata_bits_wstrb_42(fringeCommon_io_dram_2_wdata_bits_wstrb_42),
    .io_dram_2_wdata_bits_wstrb_43(fringeCommon_io_dram_2_wdata_bits_wstrb_43),
    .io_dram_2_wdata_bits_wstrb_44(fringeCommon_io_dram_2_wdata_bits_wstrb_44),
    .io_dram_2_wdata_bits_wstrb_45(fringeCommon_io_dram_2_wdata_bits_wstrb_45),
    .io_dram_2_wdata_bits_wstrb_46(fringeCommon_io_dram_2_wdata_bits_wstrb_46),
    .io_dram_2_wdata_bits_wstrb_47(fringeCommon_io_dram_2_wdata_bits_wstrb_47),
    .io_dram_2_wdata_bits_wstrb_48(fringeCommon_io_dram_2_wdata_bits_wstrb_48),
    .io_dram_2_wdata_bits_wstrb_49(fringeCommon_io_dram_2_wdata_bits_wstrb_49),
    .io_dram_2_wdata_bits_wstrb_50(fringeCommon_io_dram_2_wdata_bits_wstrb_50),
    .io_dram_2_wdata_bits_wstrb_51(fringeCommon_io_dram_2_wdata_bits_wstrb_51),
    .io_dram_2_wdata_bits_wstrb_52(fringeCommon_io_dram_2_wdata_bits_wstrb_52),
    .io_dram_2_wdata_bits_wstrb_53(fringeCommon_io_dram_2_wdata_bits_wstrb_53),
    .io_dram_2_wdata_bits_wstrb_54(fringeCommon_io_dram_2_wdata_bits_wstrb_54),
    .io_dram_2_wdata_bits_wstrb_55(fringeCommon_io_dram_2_wdata_bits_wstrb_55),
    .io_dram_2_wdata_bits_wstrb_56(fringeCommon_io_dram_2_wdata_bits_wstrb_56),
    .io_dram_2_wdata_bits_wstrb_57(fringeCommon_io_dram_2_wdata_bits_wstrb_57),
    .io_dram_2_wdata_bits_wstrb_58(fringeCommon_io_dram_2_wdata_bits_wstrb_58),
    .io_dram_2_wdata_bits_wstrb_59(fringeCommon_io_dram_2_wdata_bits_wstrb_59),
    .io_dram_2_wdata_bits_wstrb_60(fringeCommon_io_dram_2_wdata_bits_wstrb_60),
    .io_dram_2_wdata_bits_wstrb_61(fringeCommon_io_dram_2_wdata_bits_wstrb_61),
    .io_dram_2_wdata_bits_wstrb_62(fringeCommon_io_dram_2_wdata_bits_wstrb_62),
    .io_dram_2_wdata_bits_wstrb_63(fringeCommon_io_dram_2_wdata_bits_wstrb_63),
    .io_dram_2_wdata_bits_wlast(fringeCommon_io_dram_2_wdata_bits_wlast),
    .io_dram_2_rresp_ready(fringeCommon_io_dram_2_rresp_ready),
    .io_dram_2_wresp_ready(fringeCommon_io_dram_2_wresp_ready),
    .io_dram_2_wresp_valid(fringeCommon_io_dram_2_wresp_valid),
    .io_dram_2_wresp_bits_tag(fringeCommon_io_dram_2_wresp_bits_tag),
    .io_dram_3_cmd_ready(fringeCommon_io_dram_3_cmd_ready),
    .io_dram_3_cmd_valid(fringeCommon_io_dram_3_cmd_valid),
    .io_dram_3_cmd_bits_addr(fringeCommon_io_dram_3_cmd_bits_addr),
    .io_dram_3_cmd_bits_size(fringeCommon_io_dram_3_cmd_bits_size),
    .io_dram_3_cmd_bits_isWr(fringeCommon_io_dram_3_cmd_bits_isWr),
    .io_dram_3_cmd_bits_tag(fringeCommon_io_dram_3_cmd_bits_tag),
    .io_dram_3_wdata_ready(fringeCommon_io_dram_3_wdata_ready),
    .io_dram_3_wdata_valid(fringeCommon_io_dram_3_wdata_valid),
    .io_dram_3_wdata_bits_wdata_0(fringeCommon_io_dram_3_wdata_bits_wdata_0),
    .io_dram_3_wdata_bits_wdata_1(fringeCommon_io_dram_3_wdata_bits_wdata_1),
    .io_dram_3_wdata_bits_wdata_2(fringeCommon_io_dram_3_wdata_bits_wdata_2),
    .io_dram_3_wdata_bits_wdata_3(fringeCommon_io_dram_3_wdata_bits_wdata_3),
    .io_dram_3_wdata_bits_wdata_4(fringeCommon_io_dram_3_wdata_bits_wdata_4),
    .io_dram_3_wdata_bits_wdata_5(fringeCommon_io_dram_3_wdata_bits_wdata_5),
    .io_dram_3_wdata_bits_wdata_6(fringeCommon_io_dram_3_wdata_bits_wdata_6),
    .io_dram_3_wdata_bits_wdata_7(fringeCommon_io_dram_3_wdata_bits_wdata_7),
    .io_dram_3_wdata_bits_wdata_8(fringeCommon_io_dram_3_wdata_bits_wdata_8),
    .io_dram_3_wdata_bits_wdata_9(fringeCommon_io_dram_3_wdata_bits_wdata_9),
    .io_dram_3_wdata_bits_wdata_10(fringeCommon_io_dram_3_wdata_bits_wdata_10),
    .io_dram_3_wdata_bits_wdata_11(fringeCommon_io_dram_3_wdata_bits_wdata_11),
    .io_dram_3_wdata_bits_wdata_12(fringeCommon_io_dram_3_wdata_bits_wdata_12),
    .io_dram_3_wdata_bits_wdata_13(fringeCommon_io_dram_3_wdata_bits_wdata_13),
    .io_dram_3_wdata_bits_wdata_14(fringeCommon_io_dram_3_wdata_bits_wdata_14),
    .io_dram_3_wdata_bits_wdata_15(fringeCommon_io_dram_3_wdata_bits_wdata_15),
    .io_dram_3_wdata_bits_wstrb_0(fringeCommon_io_dram_3_wdata_bits_wstrb_0),
    .io_dram_3_wdata_bits_wstrb_1(fringeCommon_io_dram_3_wdata_bits_wstrb_1),
    .io_dram_3_wdata_bits_wstrb_2(fringeCommon_io_dram_3_wdata_bits_wstrb_2),
    .io_dram_3_wdata_bits_wstrb_3(fringeCommon_io_dram_3_wdata_bits_wstrb_3),
    .io_dram_3_wdata_bits_wstrb_4(fringeCommon_io_dram_3_wdata_bits_wstrb_4),
    .io_dram_3_wdata_bits_wstrb_5(fringeCommon_io_dram_3_wdata_bits_wstrb_5),
    .io_dram_3_wdata_bits_wstrb_6(fringeCommon_io_dram_3_wdata_bits_wstrb_6),
    .io_dram_3_wdata_bits_wstrb_7(fringeCommon_io_dram_3_wdata_bits_wstrb_7),
    .io_dram_3_wdata_bits_wstrb_8(fringeCommon_io_dram_3_wdata_bits_wstrb_8),
    .io_dram_3_wdata_bits_wstrb_9(fringeCommon_io_dram_3_wdata_bits_wstrb_9),
    .io_dram_3_wdata_bits_wstrb_10(fringeCommon_io_dram_3_wdata_bits_wstrb_10),
    .io_dram_3_wdata_bits_wstrb_11(fringeCommon_io_dram_3_wdata_bits_wstrb_11),
    .io_dram_3_wdata_bits_wstrb_12(fringeCommon_io_dram_3_wdata_bits_wstrb_12),
    .io_dram_3_wdata_bits_wstrb_13(fringeCommon_io_dram_3_wdata_bits_wstrb_13),
    .io_dram_3_wdata_bits_wstrb_14(fringeCommon_io_dram_3_wdata_bits_wstrb_14),
    .io_dram_3_wdata_bits_wstrb_15(fringeCommon_io_dram_3_wdata_bits_wstrb_15),
    .io_dram_3_wdata_bits_wstrb_16(fringeCommon_io_dram_3_wdata_bits_wstrb_16),
    .io_dram_3_wdata_bits_wstrb_17(fringeCommon_io_dram_3_wdata_bits_wstrb_17),
    .io_dram_3_wdata_bits_wstrb_18(fringeCommon_io_dram_3_wdata_bits_wstrb_18),
    .io_dram_3_wdata_bits_wstrb_19(fringeCommon_io_dram_3_wdata_bits_wstrb_19),
    .io_dram_3_wdata_bits_wstrb_20(fringeCommon_io_dram_3_wdata_bits_wstrb_20),
    .io_dram_3_wdata_bits_wstrb_21(fringeCommon_io_dram_3_wdata_bits_wstrb_21),
    .io_dram_3_wdata_bits_wstrb_22(fringeCommon_io_dram_3_wdata_bits_wstrb_22),
    .io_dram_3_wdata_bits_wstrb_23(fringeCommon_io_dram_3_wdata_bits_wstrb_23),
    .io_dram_3_wdata_bits_wstrb_24(fringeCommon_io_dram_3_wdata_bits_wstrb_24),
    .io_dram_3_wdata_bits_wstrb_25(fringeCommon_io_dram_3_wdata_bits_wstrb_25),
    .io_dram_3_wdata_bits_wstrb_26(fringeCommon_io_dram_3_wdata_bits_wstrb_26),
    .io_dram_3_wdata_bits_wstrb_27(fringeCommon_io_dram_3_wdata_bits_wstrb_27),
    .io_dram_3_wdata_bits_wstrb_28(fringeCommon_io_dram_3_wdata_bits_wstrb_28),
    .io_dram_3_wdata_bits_wstrb_29(fringeCommon_io_dram_3_wdata_bits_wstrb_29),
    .io_dram_3_wdata_bits_wstrb_30(fringeCommon_io_dram_3_wdata_bits_wstrb_30),
    .io_dram_3_wdata_bits_wstrb_31(fringeCommon_io_dram_3_wdata_bits_wstrb_31),
    .io_dram_3_wdata_bits_wstrb_32(fringeCommon_io_dram_3_wdata_bits_wstrb_32),
    .io_dram_3_wdata_bits_wstrb_33(fringeCommon_io_dram_3_wdata_bits_wstrb_33),
    .io_dram_3_wdata_bits_wstrb_34(fringeCommon_io_dram_3_wdata_bits_wstrb_34),
    .io_dram_3_wdata_bits_wstrb_35(fringeCommon_io_dram_3_wdata_bits_wstrb_35),
    .io_dram_3_wdata_bits_wstrb_36(fringeCommon_io_dram_3_wdata_bits_wstrb_36),
    .io_dram_3_wdata_bits_wstrb_37(fringeCommon_io_dram_3_wdata_bits_wstrb_37),
    .io_dram_3_wdata_bits_wstrb_38(fringeCommon_io_dram_3_wdata_bits_wstrb_38),
    .io_dram_3_wdata_bits_wstrb_39(fringeCommon_io_dram_3_wdata_bits_wstrb_39),
    .io_dram_3_wdata_bits_wstrb_40(fringeCommon_io_dram_3_wdata_bits_wstrb_40),
    .io_dram_3_wdata_bits_wstrb_41(fringeCommon_io_dram_3_wdata_bits_wstrb_41),
    .io_dram_3_wdata_bits_wstrb_42(fringeCommon_io_dram_3_wdata_bits_wstrb_42),
    .io_dram_3_wdata_bits_wstrb_43(fringeCommon_io_dram_3_wdata_bits_wstrb_43),
    .io_dram_3_wdata_bits_wstrb_44(fringeCommon_io_dram_3_wdata_bits_wstrb_44),
    .io_dram_3_wdata_bits_wstrb_45(fringeCommon_io_dram_3_wdata_bits_wstrb_45),
    .io_dram_3_wdata_bits_wstrb_46(fringeCommon_io_dram_3_wdata_bits_wstrb_46),
    .io_dram_3_wdata_bits_wstrb_47(fringeCommon_io_dram_3_wdata_bits_wstrb_47),
    .io_dram_3_wdata_bits_wstrb_48(fringeCommon_io_dram_3_wdata_bits_wstrb_48),
    .io_dram_3_wdata_bits_wstrb_49(fringeCommon_io_dram_3_wdata_bits_wstrb_49),
    .io_dram_3_wdata_bits_wstrb_50(fringeCommon_io_dram_3_wdata_bits_wstrb_50),
    .io_dram_3_wdata_bits_wstrb_51(fringeCommon_io_dram_3_wdata_bits_wstrb_51),
    .io_dram_3_wdata_bits_wstrb_52(fringeCommon_io_dram_3_wdata_bits_wstrb_52),
    .io_dram_3_wdata_bits_wstrb_53(fringeCommon_io_dram_3_wdata_bits_wstrb_53),
    .io_dram_3_wdata_bits_wstrb_54(fringeCommon_io_dram_3_wdata_bits_wstrb_54),
    .io_dram_3_wdata_bits_wstrb_55(fringeCommon_io_dram_3_wdata_bits_wstrb_55),
    .io_dram_3_wdata_bits_wstrb_56(fringeCommon_io_dram_3_wdata_bits_wstrb_56),
    .io_dram_3_wdata_bits_wstrb_57(fringeCommon_io_dram_3_wdata_bits_wstrb_57),
    .io_dram_3_wdata_bits_wstrb_58(fringeCommon_io_dram_3_wdata_bits_wstrb_58),
    .io_dram_3_wdata_bits_wstrb_59(fringeCommon_io_dram_3_wdata_bits_wstrb_59),
    .io_dram_3_wdata_bits_wstrb_60(fringeCommon_io_dram_3_wdata_bits_wstrb_60),
    .io_dram_3_wdata_bits_wstrb_61(fringeCommon_io_dram_3_wdata_bits_wstrb_61),
    .io_dram_3_wdata_bits_wstrb_62(fringeCommon_io_dram_3_wdata_bits_wstrb_62),
    .io_dram_3_wdata_bits_wstrb_63(fringeCommon_io_dram_3_wdata_bits_wstrb_63),
    .io_dram_3_wdata_bits_wlast(fringeCommon_io_dram_3_wdata_bits_wlast),
    .io_dram_3_rresp_ready(fringeCommon_io_dram_3_rresp_ready),
    .io_dram_3_wresp_ready(fringeCommon_io_dram_3_wresp_ready),
    .io_dram_3_wresp_valid(fringeCommon_io_dram_3_wresp_valid),
    .io_dram_3_wresp_bits_tag(fringeCommon_io_dram_3_wresp_bits_tag),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridge AXI4LiteToRFBridge ( // @[FringeZynq.scala 90:31:@151327.4]
    .clock(AXI4LiteToRFBridge_clock),
    .reset(AXI4LiteToRFBridge_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridge_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridge_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridge_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridge_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridge_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridge_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridge_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridge_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridge_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridge_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridge_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridge_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridge_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridge_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridge_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridge_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridge_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridge_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridge_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridge_io_raddr),
    .io_wen(AXI4LiteToRFBridge_io_wen),
    .io_waddr(AXI4LiteToRFBridge_io_waddr),
    .io_wdata(AXI4LiteToRFBridge_io_wdata),
    .io_rdata(AXI4LiteToRFBridge_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 131:27:@151477.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_1 ( // @[FringeZynq.scala 131:27:@151633.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_1_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_1_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_1_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_1_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_1_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_1_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_1_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_1_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_1_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_1_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_1_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_1_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_1_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_1_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_1_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_1_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_1_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_1_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_1_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_1_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_1_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_1_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_1_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_1_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_1_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_1_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_1_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_1_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_1_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_1_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_1_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_1_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_2 ( // @[FringeZynq.scala 131:27:@151789.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_2_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_2_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_2_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_2_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_2_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_2_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_2_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_2_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_2_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_2_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_2_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_2_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_2_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_2_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_2_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_2_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_2_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_2_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_2_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_2_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_2_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_2_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_2_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_2_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_2_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_2_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_2_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_2_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_2_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_2_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_2_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_2_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_3 ( // @[FringeZynq.scala 131:27:@151945.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_3_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_3_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_3_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_3_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_3_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_3_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_3_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_3_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_3_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_3_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_3_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_3_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_3_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_3_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_3_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_3_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_3_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_3_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_3_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_3_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_3_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_3_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_3_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_3_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_3_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_3_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_3_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_3_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_3_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_3_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_3_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_3_io_M_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 91:28:@151345.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 91:28:@151341.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 91:28:@151337.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 91:28:@151336.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 91:28:@151335.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 91:28:@151334.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 91:28:@151332.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 91:28:@151331.4]
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@151632.4]
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@151630.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@151629.4]
  assign io_M_AXI_0_AWVALID = MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@151622.4]
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@151620.4]
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@151618.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@151617.4]
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@151610.4]
  assign io_M_AXI_0_WDATA = MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@151608.4]
  assign io_M_AXI_0_WSTRB = MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@151607.4]
  assign io_M_AXI_0_WLAST = MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@151606.4]
  assign io_M_AXI_0_WVALID = MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@151605.4]
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@151597.4]
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@151592.4]
  assign io_M_AXI_1_AWID = MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@151788.4]
  assign io_M_AXI_1_AWADDR = MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@151786.4]
  assign io_M_AXI_1_AWLEN = MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@151785.4]
  assign io_M_AXI_1_AWVALID = MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@151778.4]
  assign io_M_AXI_1_ARID = MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@151776.4]
  assign io_M_AXI_1_ARADDR = MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@151774.4]
  assign io_M_AXI_1_ARLEN = MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@151773.4]
  assign io_M_AXI_1_ARVALID = MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@151766.4]
  assign io_M_AXI_1_WDATA = MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@151764.4]
  assign io_M_AXI_1_WSTRB = MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@151763.4]
  assign io_M_AXI_1_WLAST = MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@151762.4]
  assign io_M_AXI_1_WVALID = MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@151761.4]
  assign io_M_AXI_1_RREADY = MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@151753.4]
  assign io_M_AXI_1_BREADY = MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@151748.4]
  assign io_M_AXI_2_AWID = MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@151944.4]
  assign io_M_AXI_2_AWADDR = MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@151942.4]
  assign io_M_AXI_2_AWLEN = MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@151941.4]
  assign io_M_AXI_2_AWVALID = MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@151934.4]
  assign io_M_AXI_2_ARID = MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@151932.4]
  assign io_M_AXI_2_ARADDR = MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@151930.4]
  assign io_M_AXI_2_ARLEN = MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@151929.4]
  assign io_M_AXI_2_ARVALID = MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@151922.4]
  assign io_M_AXI_2_WDATA = MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@151920.4]
  assign io_M_AXI_2_WSTRB = MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@151919.4]
  assign io_M_AXI_2_WLAST = MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@151918.4]
  assign io_M_AXI_2_WVALID = MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@151917.4]
  assign io_M_AXI_2_RREADY = MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@151909.4]
  assign io_M_AXI_2_BREADY = MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@151904.4]
  assign io_M_AXI_3_AWID = MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@152100.4]
  assign io_M_AXI_3_AWADDR = MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@152098.4]
  assign io_M_AXI_3_AWLEN = MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@152097.4]
  assign io_M_AXI_3_AWVALID = MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@152090.4]
  assign io_M_AXI_3_ARID = MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@152088.4]
  assign io_M_AXI_3_ARADDR = MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@152086.4]
  assign io_M_AXI_3_ARLEN = MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@152085.4]
  assign io_M_AXI_3_ARVALID = MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@152078.4]
  assign io_M_AXI_3_WDATA = MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@152076.4]
  assign io_M_AXI_3_WSTRB = MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@152075.4]
  assign io_M_AXI_3_WLAST = MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@152074.4]
  assign io_M_AXI_3_WVALID = MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@152073.4]
  assign io_M_AXI_3_RREADY = MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@152065.4]
  assign io_M_AXI_3_BREADY = MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@152060.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 115:13:@151355.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 119:12:@151359.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 121:13:@151360.4]
  assign io_argIns_1 = fringeCommon_io_argIns_1; // @[FringeZynq.scala 121:13:@151361.4]
  assign io_memStreams_stores_0_cmd_ready = fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 126:17:@151448.4]
  assign io_memStreams_stores_0_data_ready = fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 126:17:@151444.4]
  assign io_memStreams_stores_0_wresp_valid = fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 126:17:@151439.4]
  assign io_memStreams_stores_0_wresp_bits = fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 126:17:@151438.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 127:11:@151473.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 127:11:@151472.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 127:11:@151471.4]
  assign fringeCommon_clock = clock; // @[:@150422.4]
  assign fringeCommon_reset = reset; // @[:@150423.4 FringeZynq.scala 117:22:@151358.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 94:27:@151349.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 95:27:@151350.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 96:27:@151351.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridge_io_wdata}; // @[FringeZynq.scala 97:27:@151352.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 116:24:@151356.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 122:27:@151363.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 122:27:@151362.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 126:17:@151447.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 126:17:@151446.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 126:17:@151445.4]
  assign fringeCommon_io_memStreams_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 126:17:@151443.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 126:17:@151442.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 126:17:@151441.4]
  assign fringeCommon_io_memStreams_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 126:17:@151440.4]
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@151591.4]
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@151584.4]
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@151481.4]
  assign fringeCommon_io_dram_0_wresp_bits_tag = MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@151480.4]
  assign fringeCommon_io_dram_1_cmd_ready = MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@151747.4]
  assign fringeCommon_io_dram_1_wdata_ready = MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@151740.4]
  assign fringeCommon_io_dram_1_wresp_valid = MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@151637.4]
  assign fringeCommon_io_dram_1_wresp_bits_tag = MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@151636.4]
  assign fringeCommon_io_dram_2_cmd_ready = MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@151903.4]
  assign fringeCommon_io_dram_2_wdata_ready = MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@151896.4]
  assign fringeCommon_io_dram_2_wresp_valid = MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@151793.4]
  assign fringeCommon_io_dram_2_wresp_bits_tag = MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@151792.4]
  assign fringeCommon_io_dram_3_cmd_ready = MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@152059.4]
  assign fringeCommon_io_dram_3_wdata_ready = MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@152052.4]
  assign fringeCommon_io_dram_3_wresp_valid = MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@151949.4]
  assign fringeCommon_io_dram_3_wresp_bits_tag = MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@151948.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 127:11:@151476.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 127:11:@151475.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 127:11:@151474.4]
  assign AXI4LiteToRFBridge_clock = clock; // @[:@151328.4]
  assign AXI4LiteToRFBridge_reset = reset; // @[:@151329.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 91:28:@151348.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 91:28:@151347.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 91:28:@151346.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 91:28:@151344.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 91:28:@151343.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 91:28:@151342.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 91:28:@151340.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 91:28:@151339.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 91:28:@151338.4]
  assign AXI4LiteToRFBridge_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 91:28:@151333.4]
  assign AXI4LiteToRFBridge_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 91:28:@151330.4]
  assign AXI4LiteToRFBridge_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 98:28:@151353.4]
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 132:21:@151590.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 132:21:@151589.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 132:21:@151588.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_isWr = fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@151586.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag = fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 132:21:@151585.4]
  assign MAGToAXI4Bridge_io_in_wdata_valid = fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 132:21:@151583.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@151567.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@151568.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@151569.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@151570.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@151571.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@151572.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@151573.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@151574.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@151575.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@151576.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@151577.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@151578.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@151579.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@151580.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@151581.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@151582.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@151503.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@151504.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@151505.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@151506.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@151507.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@151508.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@151509.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@151510.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@151511.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@151512.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@151513.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@151514.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@151515.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@151516.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@151517.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@151518.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@151519.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@151520.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@151521.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@151522.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@151523.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@151524.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@151525.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@151526.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@151527.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@151528.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@151529.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@151530.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@151531.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@151532.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@151533.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@151534.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@151535.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@151536.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@151537.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@151538.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@151539.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@151540.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@151541.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@151542.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@151543.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@151544.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@151545.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@151546.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@151547.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@151548.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@151549.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@151550.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@151551.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@151552.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@151553.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@151554.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@151555.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@151556.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@151557.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@151558.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@151559.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@151560.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@151561.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@151562.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@151563.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@151564.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@151565.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@151566.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wlast = fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@151502.4]
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 132:21:@151501.4]
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 132:21:@151482.4]
  assign MAGToAXI4Bridge_io_M_AXI_AWREADY = io_M_AXI_0_AWREADY; // @[FringeZynq.scala 133:10:@151621.4]
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY; // @[FringeZynq.scala 133:10:@151609.4]
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY; // @[FringeZynq.scala 133:10:@151604.4]
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID; // @[FringeZynq.scala 133:10:@151596.4]
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID; // @[FringeZynq.scala 133:10:@151593.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_valid = fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 132:21:@151746.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_addr = fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 132:21:@151745.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_size = fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 132:21:@151744.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_isWr = fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@151742.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_tag = fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 132:21:@151741.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_valid = fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 132:21:@151739.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@151723.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@151724.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@151725.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@151726.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@151727.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@151728.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@151729.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@151730.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@151731.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@151732.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@151733.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@151734.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@151735.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@151736.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@151737.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@151738.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@151659.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@151660.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@151661.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@151662.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@151663.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@151664.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@151665.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@151666.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@151667.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@151668.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@151669.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@151670.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@151671.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@151672.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@151673.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@151674.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@151675.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@151676.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@151677.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@151678.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@151679.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@151680.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@151681.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@151682.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@151683.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@151684.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@151685.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@151686.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@151687.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@151688.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@151689.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@151690.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@151691.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@151692.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@151693.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@151694.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@151695.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@151696.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@151697.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@151698.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@151699.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@151700.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@151701.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@151702.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@151703.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@151704.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@151705.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@151706.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@151707.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@151708.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@151709.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@151710.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@151711.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@151712.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@151713.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@151714.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@151715.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@151716.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@151717.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@151718.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@151719.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@151720.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@151721.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@151722.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wlast = fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@151658.4]
  assign MAGToAXI4Bridge_1_io_in_rresp_ready = fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 132:21:@151657.4]
  assign MAGToAXI4Bridge_1_io_in_wresp_ready = fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 132:21:@151638.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_AWREADY = io_M_AXI_1_AWREADY; // @[FringeZynq.scala 133:10:@151777.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_ARREADY = io_M_AXI_1_ARREADY; // @[FringeZynq.scala 133:10:@151765.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_WREADY = io_M_AXI_1_WREADY; // @[FringeZynq.scala 133:10:@151760.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BID = io_M_AXI_1_BID; // @[FringeZynq.scala 133:10:@151752.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BVALID = io_M_AXI_1_BVALID; // @[FringeZynq.scala 133:10:@151749.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_valid = fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 132:21:@151902.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_addr = fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 132:21:@151901.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_size = fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 132:21:@151900.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_isWr = fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@151898.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_tag = fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 132:21:@151897.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_valid = fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 132:21:@151895.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@151879.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@151880.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@151881.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@151882.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@151883.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@151884.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@151885.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@151886.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@151887.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@151888.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@151889.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@151890.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@151891.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@151892.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@151893.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@151894.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@151815.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@151816.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@151817.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@151818.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@151819.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@151820.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@151821.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@151822.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@151823.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@151824.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@151825.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@151826.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@151827.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@151828.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@151829.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@151830.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@151831.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@151832.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@151833.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@151834.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@151835.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@151836.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@151837.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@151838.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@151839.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@151840.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@151841.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@151842.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@151843.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@151844.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@151845.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@151846.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@151847.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@151848.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@151849.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@151850.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@151851.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@151852.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@151853.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@151854.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@151855.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@151856.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@151857.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@151858.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@151859.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@151860.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@151861.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@151862.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@151863.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@151864.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@151865.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@151866.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@151867.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@151868.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@151869.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@151870.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@151871.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@151872.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@151873.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@151874.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@151875.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@151876.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@151877.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@151878.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wlast = fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@151814.4]
  assign MAGToAXI4Bridge_2_io_in_rresp_ready = fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 132:21:@151813.4]
  assign MAGToAXI4Bridge_2_io_in_wresp_ready = fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 132:21:@151794.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_AWREADY = io_M_AXI_2_AWREADY; // @[FringeZynq.scala 133:10:@151933.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_ARREADY = io_M_AXI_2_ARREADY; // @[FringeZynq.scala 133:10:@151921.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_WREADY = io_M_AXI_2_WREADY; // @[FringeZynq.scala 133:10:@151916.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BID = io_M_AXI_2_BID; // @[FringeZynq.scala 133:10:@151908.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BVALID = io_M_AXI_2_BVALID; // @[FringeZynq.scala 133:10:@151905.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_valid = fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 132:21:@152058.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_addr = fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 132:21:@152057.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_size = fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 132:21:@152056.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_isWr = fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@152054.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_tag = fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 132:21:@152053.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_valid = fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 132:21:@152051.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@152035.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@152036.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@152037.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@152038.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@152039.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@152040.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@152041.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@152042.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@152043.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@152044.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@152045.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@152046.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@152047.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@152048.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@152049.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@152050.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@151971.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@151972.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@151973.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@151974.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@151975.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@151976.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@151977.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@151978.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@151979.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@151980.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@151981.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@151982.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@151983.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@151984.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@151985.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@151986.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@151987.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@151988.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@151989.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@151990.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@151991.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@151992.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@151993.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@151994.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@151995.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@151996.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@151997.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@151998.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@151999.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@152000.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@152001.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@152002.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@152003.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@152004.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@152005.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@152006.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@152007.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@152008.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@152009.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@152010.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@152011.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@152012.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@152013.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@152014.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@152015.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@152016.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@152017.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@152018.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@152019.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@152020.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@152021.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@152022.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@152023.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@152024.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@152025.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@152026.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@152027.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@152028.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@152029.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@152030.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@152031.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@152032.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@152033.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@152034.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wlast = fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@151970.4]
  assign MAGToAXI4Bridge_3_io_in_rresp_ready = fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 132:21:@151969.4]
  assign MAGToAXI4Bridge_3_io_in_wresp_ready = fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 132:21:@151950.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_AWREADY = io_M_AXI_3_AWREADY; // @[FringeZynq.scala 133:10:@152089.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_ARREADY = io_M_AXI_3_ARREADY; // @[FringeZynq.scala 133:10:@152077.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_WREADY = io_M_AXI_3_WREADY; // @[FringeZynq.scala 133:10:@152072.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BID = io_M_AXI_3_BID; // @[FringeZynq.scala 133:10:@152064.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BVALID = io_M_AXI_3_BVALID; // @[FringeZynq.scala 133:10:@152061.4]
endmodule
module SpatialIP( // @[:@152102.2]
  input          clock, // @[:@152103.4]
  input          reset, // @[:@152104.4]
  input          io_raddr, // @[:@152105.4]
  input          io_wen, // @[:@152105.4]
  input          io_waddr, // @[:@152105.4]
  input          io_wdata, // @[:@152105.4]
  output         io_rdata, // @[:@152105.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@152105.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@152105.4]
  input          io_S_AXI_AWVALID, // @[:@152105.4]
  output         io_S_AXI_AWREADY, // @[:@152105.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@152105.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@152105.4]
  input          io_S_AXI_ARVALID, // @[:@152105.4]
  output         io_S_AXI_ARREADY, // @[:@152105.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@152105.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@152105.4]
  input          io_S_AXI_WVALID, // @[:@152105.4]
  output         io_S_AXI_WREADY, // @[:@152105.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@152105.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@152105.4]
  output         io_S_AXI_RVALID, // @[:@152105.4]
  input          io_S_AXI_RREADY, // @[:@152105.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@152105.4]
  output         io_S_AXI_BVALID, // @[:@152105.4]
  input          io_S_AXI_BREADY, // @[:@152105.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@152105.4]
  output [31:0]  io_M_AXI_0_AWUSER, // @[:@152105.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@152105.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@152105.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@152105.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@152105.4]
  output         io_M_AXI_0_AWLOCK, // @[:@152105.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@152105.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@152105.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@152105.4]
  output         io_M_AXI_0_AWVALID, // @[:@152105.4]
  input          io_M_AXI_0_AWREADY, // @[:@152105.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@152105.4]
  output [31:0]  io_M_AXI_0_ARUSER, // @[:@152105.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@152105.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@152105.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@152105.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@152105.4]
  output         io_M_AXI_0_ARLOCK, // @[:@152105.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@152105.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@152105.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@152105.4]
  output         io_M_AXI_0_ARVALID, // @[:@152105.4]
  input          io_M_AXI_0_ARREADY, // @[:@152105.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@152105.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@152105.4]
  output         io_M_AXI_0_WLAST, // @[:@152105.4]
  output         io_M_AXI_0_WVALID, // @[:@152105.4]
  input          io_M_AXI_0_WREADY, // @[:@152105.4]
  input  [31:0]  io_M_AXI_0_RID, // @[:@152105.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@152105.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@152105.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@152105.4]
  input          io_M_AXI_0_RLAST, // @[:@152105.4]
  input          io_M_AXI_0_RVALID, // @[:@152105.4]
  output         io_M_AXI_0_RREADY, // @[:@152105.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@152105.4]
  input  [31:0]  io_M_AXI_0_BUSER, // @[:@152105.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@152105.4]
  input          io_M_AXI_0_BVALID, // @[:@152105.4]
  output         io_M_AXI_0_BREADY, // @[:@152105.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@152105.4]
  output [31:0]  io_M_AXI_1_AWUSER, // @[:@152105.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@152105.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@152105.4]
  output [2:0]   io_M_AXI_1_AWSIZE, // @[:@152105.4]
  output [1:0]   io_M_AXI_1_AWBURST, // @[:@152105.4]
  output         io_M_AXI_1_AWLOCK, // @[:@152105.4]
  output [3:0]   io_M_AXI_1_AWCACHE, // @[:@152105.4]
  output [2:0]   io_M_AXI_1_AWPROT, // @[:@152105.4]
  output [3:0]   io_M_AXI_1_AWQOS, // @[:@152105.4]
  output         io_M_AXI_1_AWVALID, // @[:@152105.4]
  input          io_M_AXI_1_AWREADY, // @[:@152105.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@152105.4]
  output [31:0]  io_M_AXI_1_ARUSER, // @[:@152105.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@152105.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@152105.4]
  output [2:0]   io_M_AXI_1_ARSIZE, // @[:@152105.4]
  output [1:0]   io_M_AXI_1_ARBURST, // @[:@152105.4]
  output         io_M_AXI_1_ARLOCK, // @[:@152105.4]
  output [3:0]   io_M_AXI_1_ARCACHE, // @[:@152105.4]
  output [2:0]   io_M_AXI_1_ARPROT, // @[:@152105.4]
  output [3:0]   io_M_AXI_1_ARQOS, // @[:@152105.4]
  output         io_M_AXI_1_ARVALID, // @[:@152105.4]
  input          io_M_AXI_1_ARREADY, // @[:@152105.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@152105.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@152105.4]
  output         io_M_AXI_1_WLAST, // @[:@152105.4]
  output         io_M_AXI_1_WVALID, // @[:@152105.4]
  input          io_M_AXI_1_WREADY, // @[:@152105.4]
  input  [31:0]  io_M_AXI_1_RID, // @[:@152105.4]
  input  [31:0]  io_M_AXI_1_RUSER, // @[:@152105.4]
  input  [511:0] io_M_AXI_1_RDATA, // @[:@152105.4]
  input  [1:0]   io_M_AXI_1_RRESP, // @[:@152105.4]
  input          io_M_AXI_1_RLAST, // @[:@152105.4]
  input          io_M_AXI_1_RVALID, // @[:@152105.4]
  output         io_M_AXI_1_RREADY, // @[:@152105.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@152105.4]
  input  [31:0]  io_M_AXI_1_BUSER, // @[:@152105.4]
  input  [1:0]   io_M_AXI_1_BRESP, // @[:@152105.4]
  input          io_M_AXI_1_BVALID, // @[:@152105.4]
  output         io_M_AXI_1_BREADY, // @[:@152105.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@152105.4]
  output [31:0]  io_M_AXI_2_AWUSER, // @[:@152105.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@152105.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@152105.4]
  output [2:0]   io_M_AXI_2_AWSIZE, // @[:@152105.4]
  output [1:0]   io_M_AXI_2_AWBURST, // @[:@152105.4]
  output         io_M_AXI_2_AWLOCK, // @[:@152105.4]
  output [3:0]   io_M_AXI_2_AWCACHE, // @[:@152105.4]
  output [2:0]   io_M_AXI_2_AWPROT, // @[:@152105.4]
  output [3:0]   io_M_AXI_2_AWQOS, // @[:@152105.4]
  output         io_M_AXI_2_AWVALID, // @[:@152105.4]
  input          io_M_AXI_2_AWREADY, // @[:@152105.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@152105.4]
  output [31:0]  io_M_AXI_2_ARUSER, // @[:@152105.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@152105.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@152105.4]
  output [2:0]   io_M_AXI_2_ARSIZE, // @[:@152105.4]
  output [1:0]   io_M_AXI_2_ARBURST, // @[:@152105.4]
  output         io_M_AXI_2_ARLOCK, // @[:@152105.4]
  output [3:0]   io_M_AXI_2_ARCACHE, // @[:@152105.4]
  output [2:0]   io_M_AXI_2_ARPROT, // @[:@152105.4]
  output [3:0]   io_M_AXI_2_ARQOS, // @[:@152105.4]
  output         io_M_AXI_2_ARVALID, // @[:@152105.4]
  input          io_M_AXI_2_ARREADY, // @[:@152105.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@152105.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@152105.4]
  output         io_M_AXI_2_WLAST, // @[:@152105.4]
  output         io_M_AXI_2_WVALID, // @[:@152105.4]
  input          io_M_AXI_2_WREADY, // @[:@152105.4]
  input  [31:0]  io_M_AXI_2_RID, // @[:@152105.4]
  input  [31:0]  io_M_AXI_2_RUSER, // @[:@152105.4]
  input  [511:0] io_M_AXI_2_RDATA, // @[:@152105.4]
  input  [1:0]   io_M_AXI_2_RRESP, // @[:@152105.4]
  input          io_M_AXI_2_RLAST, // @[:@152105.4]
  input          io_M_AXI_2_RVALID, // @[:@152105.4]
  output         io_M_AXI_2_RREADY, // @[:@152105.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@152105.4]
  input  [31:0]  io_M_AXI_2_BUSER, // @[:@152105.4]
  input  [1:0]   io_M_AXI_2_BRESP, // @[:@152105.4]
  input          io_M_AXI_2_BVALID, // @[:@152105.4]
  output         io_M_AXI_2_BREADY, // @[:@152105.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@152105.4]
  output [31:0]  io_M_AXI_3_AWUSER, // @[:@152105.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@152105.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@152105.4]
  output [2:0]   io_M_AXI_3_AWSIZE, // @[:@152105.4]
  output [1:0]   io_M_AXI_3_AWBURST, // @[:@152105.4]
  output         io_M_AXI_3_AWLOCK, // @[:@152105.4]
  output [3:0]   io_M_AXI_3_AWCACHE, // @[:@152105.4]
  output [2:0]   io_M_AXI_3_AWPROT, // @[:@152105.4]
  output [3:0]   io_M_AXI_3_AWQOS, // @[:@152105.4]
  output         io_M_AXI_3_AWVALID, // @[:@152105.4]
  input          io_M_AXI_3_AWREADY, // @[:@152105.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@152105.4]
  output [31:0]  io_M_AXI_3_ARUSER, // @[:@152105.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@152105.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@152105.4]
  output [2:0]   io_M_AXI_3_ARSIZE, // @[:@152105.4]
  output [1:0]   io_M_AXI_3_ARBURST, // @[:@152105.4]
  output         io_M_AXI_3_ARLOCK, // @[:@152105.4]
  output [3:0]   io_M_AXI_3_ARCACHE, // @[:@152105.4]
  output [2:0]   io_M_AXI_3_ARPROT, // @[:@152105.4]
  output [3:0]   io_M_AXI_3_ARQOS, // @[:@152105.4]
  output         io_M_AXI_3_ARVALID, // @[:@152105.4]
  input          io_M_AXI_3_ARREADY, // @[:@152105.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@152105.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@152105.4]
  output         io_M_AXI_3_WLAST, // @[:@152105.4]
  output         io_M_AXI_3_WVALID, // @[:@152105.4]
  input          io_M_AXI_3_WREADY, // @[:@152105.4]
  input  [31:0]  io_M_AXI_3_RID, // @[:@152105.4]
  input  [31:0]  io_M_AXI_3_RUSER, // @[:@152105.4]
  input  [511:0] io_M_AXI_3_RDATA, // @[:@152105.4]
  input  [1:0]   io_M_AXI_3_RRESP, // @[:@152105.4]
  input          io_M_AXI_3_RLAST, // @[:@152105.4]
  input          io_M_AXI_3_RVALID, // @[:@152105.4]
  output         io_M_AXI_3_RREADY, // @[:@152105.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@152105.4]
  input  [31:0]  io_M_AXI_3_BUSER, // @[:@152105.4]
  input  [1:0]   io_M_AXI_3_BRESP, // @[:@152105.4]
  input          io_M_AXI_3_BVALID, // @[:@152105.4]
  output         io_M_AXI_3_BREADY, // @[:@152105.4]
  input          io_TOP_AXI_AWID, // @[:@152105.4]
  input          io_TOP_AXI_AWUSER, // @[:@152105.4]
  input  [31:0]  io_TOP_AXI_AWADDR, // @[:@152105.4]
  input  [7:0]   io_TOP_AXI_AWLEN, // @[:@152105.4]
  input  [2:0]   io_TOP_AXI_AWSIZE, // @[:@152105.4]
  input  [1:0]   io_TOP_AXI_AWBURST, // @[:@152105.4]
  input          io_TOP_AXI_AWLOCK, // @[:@152105.4]
  input  [3:0]   io_TOP_AXI_AWCACHE, // @[:@152105.4]
  input  [2:0]   io_TOP_AXI_AWPROT, // @[:@152105.4]
  input  [3:0]   io_TOP_AXI_AWQOS, // @[:@152105.4]
  input          io_TOP_AXI_AWVALID, // @[:@152105.4]
  input          io_TOP_AXI_AWREADY, // @[:@152105.4]
  input          io_TOP_AXI_ARID, // @[:@152105.4]
  input          io_TOP_AXI_ARUSER, // @[:@152105.4]
  input  [31:0]  io_TOP_AXI_ARADDR, // @[:@152105.4]
  input  [7:0]   io_TOP_AXI_ARLEN, // @[:@152105.4]
  input  [2:0]   io_TOP_AXI_ARSIZE, // @[:@152105.4]
  input  [1:0]   io_TOP_AXI_ARBURST, // @[:@152105.4]
  input          io_TOP_AXI_ARLOCK, // @[:@152105.4]
  input  [3:0]   io_TOP_AXI_ARCACHE, // @[:@152105.4]
  input  [2:0]   io_TOP_AXI_ARPROT, // @[:@152105.4]
  input  [3:0]   io_TOP_AXI_ARQOS, // @[:@152105.4]
  input          io_TOP_AXI_ARVALID, // @[:@152105.4]
  input          io_TOP_AXI_ARREADY, // @[:@152105.4]
  input  [31:0]  io_TOP_AXI_WDATA, // @[:@152105.4]
  input  [63:0]  io_TOP_AXI_WSTRB, // @[:@152105.4]
  input          io_TOP_AXI_WLAST, // @[:@152105.4]
  input          io_TOP_AXI_WVALID, // @[:@152105.4]
  input          io_TOP_AXI_WREADY, // @[:@152105.4]
  input          io_TOP_AXI_RID, // @[:@152105.4]
  input          io_TOP_AXI_RUSER, // @[:@152105.4]
  input  [31:0]  io_TOP_AXI_RDATA, // @[:@152105.4]
  input  [1:0]   io_TOP_AXI_RRESP, // @[:@152105.4]
  input          io_TOP_AXI_RLAST, // @[:@152105.4]
  input          io_TOP_AXI_RVALID, // @[:@152105.4]
  input          io_TOP_AXI_RREADY, // @[:@152105.4]
  input          io_TOP_AXI_BID, // @[:@152105.4]
  input          io_TOP_AXI_BUSER, // @[:@152105.4]
  input  [1:0]   io_TOP_AXI_BRESP, // @[:@152105.4]
  input          io_TOP_AXI_BVALID, // @[:@152105.4]
  input          io_TOP_AXI_BREADY, // @[:@152105.4]
  input          io_DWIDTH_AXI_AWID, // @[:@152105.4]
  input          io_DWIDTH_AXI_AWUSER, // @[:@152105.4]
  input  [31:0]  io_DWIDTH_AXI_AWADDR, // @[:@152105.4]
  input  [7:0]   io_DWIDTH_AXI_AWLEN, // @[:@152105.4]
  input  [2:0]   io_DWIDTH_AXI_AWSIZE, // @[:@152105.4]
  input  [1:0]   io_DWIDTH_AXI_AWBURST, // @[:@152105.4]
  input          io_DWIDTH_AXI_AWLOCK, // @[:@152105.4]
  input  [3:0]   io_DWIDTH_AXI_AWCACHE, // @[:@152105.4]
  input  [2:0]   io_DWIDTH_AXI_AWPROT, // @[:@152105.4]
  input  [3:0]   io_DWIDTH_AXI_AWQOS, // @[:@152105.4]
  input          io_DWIDTH_AXI_AWVALID, // @[:@152105.4]
  input          io_DWIDTH_AXI_AWREADY, // @[:@152105.4]
  input          io_DWIDTH_AXI_ARID, // @[:@152105.4]
  input          io_DWIDTH_AXI_ARUSER, // @[:@152105.4]
  input  [31:0]  io_DWIDTH_AXI_ARADDR, // @[:@152105.4]
  input  [7:0]   io_DWIDTH_AXI_ARLEN, // @[:@152105.4]
  input  [2:0]   io_DWIDTH_AXI_ARSIZE, // @[:@152105.4]
  input  [1:0]   io_DWIDTH_AXI_ARBURST, // @[:@152105.4]
  input          io_DWIDTH_AXI_ARLOCK, // @[:@152105.4]
  input  [3:0]   io_DWIDTH_AXI_ARCACHE, // @[:@152105.4]
  input  [2:0]   io_DWIDTH_AXI_ARPROT, // @[:@152105.4]
  input  [3:0]   io_DWIDTH_AXI_ARQOS, // @[:@152105.4]
  input          io_DWIDTH_AXI_ARVALID, // @[:@152105.4]
  input          io_DWIDTH_AXI_ARREADY, // @[:@152105.4]
  input  [31:0]  io_DWIDTH_AXI_WDATA, // @[:@152105.4]
  input  [63:0]  io_DWIDTH_AXI_WSTRB, // @[:@152105.4]
  input          io_DWIDTH_AXI_WLAST, // @[:@152105.4]
  input          io_DWIDTH_AXI_WVALID, // @[:@152105.4]
  input          io_DWIDTH_AXI_WREADY, // @[:@152105.4]
  input          io_DWIDTH_AXI_RID, // @[:@152105.4]
  input          io_DWIDTH_AXI_RUSER, // @[:@152105.4]
  input  [31:0]  io_DWIDTH_AXI_RDATA, // @[:@152105.4]
  input  [1:0]   io_DWIDTH_AXI_RRESP, // @[:@152105.4]
  input          io_DWIDTH_AXI_RLAST, // @[:@152105.4]
  input          io_DWIDTH_AXI_RVALID, // @[:@152105.4]
  input          io_DWIDTH_AXI_RREADY, // @[:@152105.4]
  input          io_DWIDTH_AXI_BID, // @[:@152105.4]
  input          io_DWIDTH_AXI_BUSER, // @[:@152105.4]
  input  [1:0]   io_DWIDTH_AXI_BRESP, // @[:@152105.4]
  input          io_DWIDTH_AXI_BVALID, // @[:@152105.4]
  input          io_DWIDTH_AXI_BREADY, // @[:@152105.4]
  input          io_PROTOCOL_AXI_AWID, // @[:@152105.4]
  input          io_PROTOCOL_AXI_AWUSER, // @[:@152105.4]
  input  [31:0]  io_PROTOCOL_AXI_AWADDR, // @[:@152105.4]
  input  [7:0]   io_PROTOCOL_AXI_AWLEN, // @[:@152105.4]
  input  [2:0]   io_PROTOCOL_AXI_AWSIZE, // @[:@152105.4]
  input  [1:0]   io_PROTOCOL_AXI_AWBURST, // @[:@152105.4]
  input          io_PROTOCOL_AXI_AWLOCK, // @[:@152105.4]
  input  [3:0]   io_PROTOCOL_AXI_AWCACHE, // @[:@152105.4]
  input  [2:0]   io_PROTOCOL_AXI_AWPROT, // @[:@152105.4]
  input  [3:0]   io_PROTOCOL_AXI_AWQOS, // @[:@152105.4]
  input          io_PROTOCOL_AXI_AWVALID, // @[:@152105.4]
  input          io_PROTOCOL_AXI_AWREADY, // @[:@152105.4]
  input          io_PROTOCOL_AXI_ARID, // @[:@152105.4]
  input          io_PROTOCOL_AXI_ARUSER, // @[:@152105.4]
  input  [31:0]  io_PROTOCOL_AXI_ARADDR, // @[:@152105.4]
  input  [7:0]   io_PROTOCOL_AXI_ARLEN, // @[:@152105.4]
  input  [2:0]   io_PROTOCOL_AXI_ARSIZE, // @[:@152105.4]
  input  [1:0]   io_PROTOCOL_AXI_ARBURST, // @[:@152105.4]
  input          io_PROTOCOL_AXI_ARLOCK, // @[:@152105.4]
  input  [3:0]   io_PROTOCOL_AXI_ARCACHE, // @[:@152105.4]
  input  [2:0]   io_PROTOCOL_AXI_ARPROT, // @[:@152105.4]
  input  [3:0]   io_PROTOCOL_AXI_ARQOS, // @[:@152105.4]
  input          io_PROTOCOL_AXI_ARVALID, // @[:@152105.4]
  input          io_PROTOCOL_AXI_ARREADY, // @[:@152105.4]
  input  [31:0]  io_PROTOCOL_AXI_WDATA, // @[:@152105.4]
  input  [63:0]  io_PROTOCOL_AXI_WSTRB, // @[:@152105.4]
  input          io_PROTOCOL_AXI_WLAST, // @[:@152105.4]
  input          io_PROTOCOL_AXI_WVALID, // @[:@152105.4]
  input          io_PROTOCOL_AXI_WREADY, // @[:@152105.4]
  input          io_PROTOCOL_AXI_RID, // @[:@152105.4]
  input          io_PROTOCOL_AXI_RUSER, // @[:@152105.4]
  input  [31:0]  io_PROTOCOL_AXI_RDATA, // @[:@152105.4]
  input  [1:0]   io_PROTOCOL_AXI_RRESP, // @[:@152105.4]
  input          io_PROTOCOL_AXI_RLAST, // @[:@152105.4]
  input          io_PROTOCOL_AXI_RVALID, // @[:@152105.4]
  input          io_PROTOCOL_AXI_RREADY, // @[:@152105.4]
  input          io_PROTOCOL_AXI_BID, // @[:@152105.4]
  input          io_PROTOCOL_AXI_BUSER, // @[:@152105.4]
  input  [1:0]   io_PROTOCOL_AXI_BRESP, // @[:@152105.4]
  input          io_PROTOCOL_AXI_BVALID, // @[:@152105.4]
  input          io_PROTOCOL_AXI_BREADY, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_AWID, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_AWUSER, // @[:@152105.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_AWADDR, // @[:@152105.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_AWLEN, // @[:@152105.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWSIZE, // @[:@152105.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_AWBURST, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_AWLOCK, // @[:@152105.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWCACHE, // @[:@152105.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWPROT, // @[:@152105.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWQOS, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_AWVALID, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_AWREADY, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_ARID, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_ARUSER, // @[:@152105.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_ARADDR, // @[:@152105.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_ARLEN, // @[:@152105.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARSIZE, // @[:@152105.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_ARBURST, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_ARLOCK, // @[:@152105.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARCACHE, // @[:@152105.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARPROT, // @[:@152105.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARQOS, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_ARVALID, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_ARREADY, // @[:@152105.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_WDATA, // @[:@152105.4]
  input  [63:0]  io_CLOCKCONVERT_AXI_WSTRB, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_WLAST, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_WVALID, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_WREADY, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_RID, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_RUSER, // @[:@152105.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_RDATA, // @[:@152105.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_RRESP, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_RLAST, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_RVALID, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_RREADY, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_BID, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_BUSER, // @[:@152105.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_BRESP, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_BVALID, // @[:@152105.4]
  input          io_CLOCKCONVERT_AXI_BREADY // @[:@152105.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@152107.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@152107.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@152107.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@152107.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@152107.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@152107.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@152107.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@152107.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@152107.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@152107.4]
  wire  FringeZynq_clock; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_reset; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[Zynq.scala 18:24:@152249.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[Zynq.scala 18:24:@152249.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[Zynq.scala 18:24:@152249.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 18:24:@152249.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 18:24:@152249.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_0_AWREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 18:24:@152249.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_0_ARREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [511:0] FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 18:24:@152249.4]
  wire [63:0] FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_0_WREADY; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_0_BID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_0_BVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 18:24:@152249.4]
  wire [7:0] FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_1_AWREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 18:24:@152249.4]
  wire [7:0] FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_1_ARREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [511:0] FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 18:24:@152249.4]
  wire [63:0] FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_1_WREADY; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_1_BID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_1_BVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 18:24:@152249.4]
  wire [7:0] FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_2_AWREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 18:24:@152249.4]
  wire [7:0] FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_2_ARREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [511:0] FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 18:24:@152249.4]
  wire [63:0] FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_2_WREADY; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_2_BID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_2_BVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 18:24:@152249.4]
  wire [7:0] FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_3_AWREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 18:24:@152249.4]
  wire [7:0] FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_3_ARREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [511:0] FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 18:24:@152249.4]
  wire [63:0] FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_3_WREADY; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_M_AXI_3_BID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_3_BVALID; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_enable; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_done; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_reset; // @[Zynq.scala 18:24:@152249.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[Zynq.scala 18:24:@152249.4]
  wire [63:0] FringeZynq_io_argIns_1; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[Zynq.scala 18:24:@152249.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 18:24:@152249.4]
  wire [63:0] FringeZynq_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_memStreams_stores_0_data_valid; // @[Zynq.scala 18:24:@152249.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 18:24:@152249.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 18:24:@152249.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 18:24:@152249.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 18:24:@152249.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@152107.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  FringeZynq FringeZynq ( // @[Zynq.scala 18:24:@152249.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWID(FringeZynq_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeZynq_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_AWVALID(FringeZynq_io_M_AXI_0_AWVALID),
    .io_M_AXI_0_AWREADY(FringeZynq_io_M_AXI_0_AWREADY),
    .io_M_AXI_0_ARID(FringeZynq_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeZynq_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeZynq_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeZynq_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WDATA(FringeZynq_io_M_AXI_0_WDATA),
    .io_M_AXI_0_WSTRB(FringeZynq_io_M_AXI_0_WSTRB),
    .io_M_AXI_0_WLAST(FringeZynq_io_M_AXI_0_WLAST),
    .io_M_AXI_0_WVALID(FringeZynq_io_M_AXI_0_WVALID),
    .io_M_AXI_0_WREADY(FringeZynq_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RREADY(FringeZynq_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeZynq_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeZynq_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeZynq_io_M_AXI_0_BREADY),
    .io_M_AXI_1_AWID(FringeZynq_io_M_AXI_1_AWID),
    .io_M_AXI_1_AWADDR(FringeZynq_io_M_AXI_1_AWADDR),
    .io_M_AXI_1_AWLEN(FringeZynq_io_M_AXI_1_AWLEN),
    .io_M_AXI_1_AWVALID(FringeZynq_io_M_AXI_1_AWVALID),
    .io_M_AXI_1_AWREADY(FringeZynq_io_M_AXI_1_AWREADY),
    .io_M_AXI_1_ARID(FringeZynq_io_M_AXI_1_ARID),
    .io_M_AXI_1_ARADDR(FringeZynq_io_M_AXI_1_ARADDR),
    .io_M_AXI_1_ARLEN(FringeZynq_io_M_AXI_1_ARLEN),
    .io_M_AXI_1_ARVALID(FringeZynq_io_M_AXI_1_ARVALID),
    .io_M_AXI_1_ARREADY(FringeZynq_io_M_AXI_1_ARREADY),
    .io_M_AXI_1_WDATA(FringeZynq_io_M_AXI_1_WDATA),
    .io_M_AXI_1_WSTRB(FringeZynq_io_M_AXI_1_WSTRB),
    .io_M_AXI_1_WLAST(FringeZynq_io_M_AXI_1_WLAST),
    .io_M_AXI_1_WVALID(FringeZynq_io_M_AXI_1_WVALID),
    .io_M_AXI_1_WREADY(FringeZynq_io_M_AXI_1_WREADY),
    .io_M_AXI_1_RREADY(FringeZynq_io_M_AXI_1_RREADY),
    .io_M_AXI_1_BID(FringeZynq_io_M_AXI_1_BID),
    .io_M_AXI_1_BVALID(FringeZynq_io_M_AXI_1_BVALID),
    .io_M_AXI_1_BREADY(FringeZynq_io_M_AXI_1_BREADY),
    .io_M_AXI_2_AWID(FringeZynq_io_M_AXI_2_AWID),
    .io_M_AXI_2_AWADDR(FringeZynq_io_M_AXI_2_AWADDR),
    .io_M_AXI_2_AWLEN(FringeZynq_io_M_AXI_2_AWLEN),
    .io_M_AXI_2_AWVALID(FringeZynq_io_M_AXI_2_AWVALID),
    .io_M_AXI_2_AWREADY(FringeZynq_io_M_AXI_2_AWREADY),
    .io_M_AXI_2_ARID(FringeZynq_io_M_AXI_2_ARID),
    .io_M_AXI_2_ARADDR(FringeZynq_io_M_AXI_2_ARADDR),
    .io_M_AXI_2_ARLEN(FringeZynq_io_M_AXI_2_ARLEN),
    .io_M_AXI_2_ARVALID(FringeZynq_io_M_AXI_2_ARVALID),
    .io_M_AXI_2_ARREADY(FringeZynq_io_M_AXI_2_ARREADY),
    .io_M_AXI_2_WDATA(FringeZynq_io_M_AXI_2_WDATA),
    .io_M_AXI_2_WSTRB(FringeZynq_io_M_AXI_2_WSTRB),
    .io_M_AXI_2_WLAST(FringeZynq_io_M_AXI_2_WLAST),
    .io_M_AXI_2_WVALID(FringeZynq_io_M_AXI_2_WVALID),
    .io_M_AXI_2_WREADY(FringeZynq_io_M_AXI_2_WREADY),
    .io_M_AXI_2_RREADY(FringeZynq_io_M_AXI_2_RREADY),
    .io_M_AXI_2_BID(FringeZynq_io_M_AXI_2_BID),
    .io_M_AXI_2_BVALID(FringeZynq_io_M_AXI_2_BVALID),
    .io_M_AXI_2_BREADY(FringeZynq_io_M_AXI_2_BREADY),
    .io_M_AXI_3_AWID(FringeZynq_io_M_AXI_3_AWID),
    .io_M_AXI_3_AWADDR(FringeZynq_io_M_AXI_3_AWADDR),
    .io_M_AXI_3_AWLEN(FringeZynq_io_M_AXI_3_AWLEN),
    .io_M_AXI_3_AWVALID(FringeZynq_io_M_AXI_3_AWVALID),
    .io_M_AXI_3_AWREADY(FringeZynq_io_M_AXI_3_AWREADY),
    .io_M_AXI_3_ARID(FringeZynq_io_M_AXI_3_ARID),
    .io_M_AXI_3_ARADDR(FringeZynq_io_M_AXI_3_ARADDR),
    .io_M_AXI_3_ARLEN(FringeZynq_io_M_AXI_3_ARLEN),
    .io_M_AXI_3_ARVALID(FringeZynq_io_M_AXI_3_ARVALID),
    .io_M_AXI_3_ARREADY(FringeZynq_io_M_AXI_3_ARREADY),
    .io_M_AXI_3_WDATA(FringeZynq_io_M_AXI_3_WDATA),
    .io_M_AXI_3_WSTRB(FringeZynq_io_M_AXI_3_WSTRB),
    .io_M_AXI_3_WLAST(FringeZynq_io_M_AXI_3_WLAST),
    .io_M_AXI_3_WVALID(FringeZynq_io_M_AXI_3_WVALID),
    .io_M_AXI_3_WREADY(FringeZynq_io_M_AXI_3_WREADY),
    .io_M_AXI_3_RREADY(FringeZynq_io_M_AXI_3_RREADY),
    .io_M_AXI_3_BID(FringeZynq_io_M_AXI_3_BID),
    .io_M_AXI_3_BVALID(FringeZynq_io_M_AXI_3_BVALID),
    .io_M_AXI_3_BREADY(FringeZynq_io_M_AXI_3_BREADY),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argIns_1(FringeZynq_io_argIns_1),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(FringeZynq_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(FringeZynq_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(FringeZynq_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(FringeZynq_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(FringeZynq_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(FringeZynq_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(FringeZynq_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(FringeZynq_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(FringeZynq_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(FringeZynq_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(FringeZynq_io_memStreams_stores_0_wresp_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 21:21:@152267.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 21:21:@152263.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 21:21:@152259.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 21:21:@152258.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 21:21:@152257.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 21:21:@152256.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 21:21:@152254.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 21:21:@152253.4]
  assign io_M_AXI_0_AWID = FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 24:14:@152311.4]
  assign io_M_AXI_0_AWUSER = 32'h0; // @[Zynq.scala 24:14:@152310.4]
  assign io_M_AXI_0_AWADDR = FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 24:14:@152309.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 24:14:@152308.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@152307.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[Zynq.scala 24:14:@152306.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@152305.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@152304.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[Zynq.scala 24:14:@152303.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[Zynq.scala 24:14:@152302.4]
  assign io_M_AXI_0_AWVALID = FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 24:14:@152301.4]
  assign io_M_AXI_0_ARID = FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 24:14:@152299.4]
  assign io_M_AXI_0_ARUSER = 32'h0; // @[Zynq.scala 24:14:@152298.4]
  assign io_M_AXI_0_ARADDR = FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 24:14:@152297.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 24:14:@152296.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@152295.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[Zynq.scala 24:14:@152294.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@152293.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@152292.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[Zynq.scala 24:14:@152291.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[Zynq.scala 24:14:@152290.4]
  assign io_M_AXI_0_ARVALID = FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 24:14:@152289.4]
  assign io_M_AXI_0_WDATA = FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 24:14:@152287.4]
  assign io_M_AXI_0_WSTRB = FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 24:14:@152286.4]
  assign io_M_AXI_0_WLAST = FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 24:14:@152285.4]
  assign io_M_AXI_0_WVALID = FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 24:14:@152284.4]
  assign io_M_AXI_0_RREADY = FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 24:14:@152276.4]
  assign io_M_AXI_0_BREADY = FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 24:14:@152271.4]
  assign io_M_AXI_1_AWID = FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 24:14:@152352.4]
  assign io_M_AXI_1_AWUSER = 32'h0; // @[Zynq.scala 24:14:@152351.4]
  assign io_M_AXI_1_AWADDR = FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 24:14:@152350.4]
  assign io_M_AXI_1_AWLEN = FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 24:14:@152349.4]
  assign io_M_AXI_1_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@152348.4]
  assign io_M_AXI_1_AWBURST = 2'h1; // @[Zynq.scala 24:14:@152347.4]
  assign io_M_AXI_1_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@152346.4]
  assign io_M_AXI_1_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@152345.4]
  assign io_M_AXI_1_AWPROT = 3'h0; // @[Zynq.scala 24:14:@152344.4]
  assign io_M_AXI_1_AWQOS = 4'h0; // @[Zynq.scala 24:14:@152343.4]
  assign io_M_AXI_1_AWVALID = FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 24:14:@152342.4]
  assign io_M_AXI_1_ARID = FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 24:14:@152340.4]
  assign io_M_AXI_1_ARUSER = 32'h0; // @[Zynq.scala 24:14:@152339.4]
  assign io_M_AXI_1_ARADDR = FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 24:14:@152338.4]
  assign io_M_AXI_1_ARLEN = FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 24:14:@152337.4]
  assign io_M_AXI_1_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@152336.4]
  assign io_M_AXI_1_ARBURST = 2'h1; // @[Zynq.scala 24:14:@152335.4]
  assign io_M_AXI_1_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@152334.4]
  assign io_M_AXI_1_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@152333.4]
  assign io_M_AXI_1_ARPROT = 3'h0; // @[Zynq.scala 24:14:@152332.4]
  assign io_M_AXI_1_ARQOS = 4'h0; // @[Zynq.scala 24:14:@152331.4]
  assign io_M_AXI_1_ARVALID = FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 24:14:@152330.4]
  assign io_M_AXI_1_WDATA = FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 24:14:@152328.4]
  assign io_M_AXI_1_WSTRB = FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 24:14:@152327.4]
  assign io_M_AXI_1_WLAST = FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 24:14:@152326.4]
  assign io_M_AXI_1_WVALID = FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 24:14:@152325.4]
  assign io_M_AXI_1_RREADY = FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 24:14:@152317.4]
  assign io_M_AXI_1_BREADY = FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 24:14:@152312.4]
  assign io_M_AXI_2_AWID = FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 24:14:@152393.4]
  assign io_M_AXI_2_AWUSER = 32'h0; // @[Zynq.scala 24:14:@152392.4]
  assign io_M_AXI_2_AWADDR = FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 24:14:@152391.4]
  assign io_M_AXI_2_AWLEN = FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 24:14:@152390.4]
  assign io_M_AXI_2_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@152389.4]
  assign io_M_AXI_2_AWBURST = 2'h1; // @[Zynq.scala 24:14:@152388.4]
  assign io_M_AXI_2_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@152387.4]
  assign io_M_AXI_2_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@152386.4]
  assign io_M_AXI_2_AWPROT = 3'h0; // @[Zynq.scala 24:14:@152385.4]
  assign io_M_AXI_2_AWQOS = 4'h0; // @[Zynq.scala 24:14:@152384.4]
  assign io_M_AXI_2_AWVALID = FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 24:14:@152383.4]
  assign io_M_AXI_2_ARID = FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 24:14:@152381.4]
  assign io_M_AXI_2_ARUSER = 32'h0; // @[Zynq.scala 24:14:@152380.4]
  assign io_M_AXI_2_ARADDR = FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 24:14:@152379.4]
  assign io_M_AXI_2_ARLEN = FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 24:14:@152378.4]
  assign io_M_AXI_2_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@152377.4]
  assign io_M_AXI_2_ARBURST = 2'h1; // @[Zynq.scala 24:14:@152376.4]
  assign io_M_AXI_2_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@152375.4]
  assign io_M_AXI_2_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@152374.4]
  assign io_M_AXI_2_ARPROT = 3'h0; // @[Zynq.scala 24:14:@152373.4]
  assign io_M_AXI_2_ARQOS = 4'h0; // @[Zynq.scala 24:14:@152372.4]
  assign io_M_AXI_2_ARVALID = FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 24:14:@152371.4]
  assign io_M_AXI_2_WDATA = FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 24:14:@152369.4]
  assign io_M_AXI_2_WSTRB = FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 24:14:@152368.4]
  assign io_M_AXI_2_WLAST = FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 24:14:@152367.4]
  assign io_M_AXI_2_WVALID = FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 24:14:@152366.4]
  assign io_M_AXI_2_RREADY = FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 24:14:@152358.4]
  assign io_M_AXI_2_BREADY = FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 24:14:@152353.4]
  assign io_M_AXI_3_AWID = FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 24:14:@152434.4]
  assign io_M_AXI_3_AWUSER = 32'h0; // @[Zynq.scala 24:14:@152433.4]
  assign io_M_AXI_3_AWADDR = FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 24:14:@152432.4]
  assign io_M_AXI_3_AWLEN = FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 24:14:@152431.4]
  assign io_M_AXI_3_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@152430.4]
  assign io_M_AXI_3_AWBURST = 2'h1; // @[Zynq.scala 24:14:@152429.4]
  assign io_M_AXI_3_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@152428.4]
  assign io_M_AXI_3_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@152427.4]
  assign io_M_AXI_3_AWPROT = 3'h0; // @[Zynq.scala 24:14:@152426.4]
  assign io_M_AXI_3_AWQOS = 4'h0; // @[Zynq.scala 24:14:@152425.4]
  assign io_M_AXI_3_AWVALID = FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 24:14:@152424.4]
  assign io_M_AXI_3_ARID = FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 24:14:@152422.4]
  assign io_M_AXI_3_ARUSER = 32'h0; // @[Zynq.scala 24:14:@152421.4]
  assign io_M_AXI_3_ARADDR = FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 24:14:@152420.4]
  assign io_M_AXI_3_ARLEN = FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 24:14:@152419.4]
  assign io_M_AXI_3_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@152418.4]
  assign io_M_AXI_3_ARBURST = 2'h1; // @[Zynq.scala 24:14:@152417.4]
  assign io_M_AXI_3_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@152416.4]
  assign io_M_AXI_3_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@152415.4]
  assign io_M_AXI_3_ARPROT = 3'h0; // @[Zynq.scala 24:14:@152414.4]
  assign io_M_AXI_3_ARQOS = 4'h0; // @[Zynq.scala 24:14:@152413.4]
  assign io_M_AXI_3_ARVALID = FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 24:14:@152412.4]
  assign io_M_AXI_3_WDATA = FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 24:14:@152410.4]
  assign io_M_AXI_3_WSTRB = FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 24:14:@152409.4]
  assign io_M_AXI_3_WLAST = FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 24:14:@152408.4]
  assign io_M_AXI_3_WVALID = FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 24:14:@152407.4]
  assign io_M_AXI_3_RREADY = FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 24:14:@152399.4]
  assign io_M_AXI_3_BREADY = FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 24:14:@152394.4]
  assign accel_clock = clock; // @[:@152108.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@152109.4 Zynq.scala 54:17:@152723.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[Zynq.scala 51:21:@152718.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@152711.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@152706.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[Zynq.scala 49:26:@152690.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[Zynq.scala 49:26:@152691.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[Zynq.scala 49:26:@152692.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[Zynq.scala 49:26:@152693.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[Zynq.scala 49:26:@152694.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[Zynq.scala 49:26:@152695.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[Zynq.scala 49:26:@152696.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[Zynq.scala 49:26:@152697.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[Zynq.scala 49:26:@152698.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[Zynq.scala 49:26:@152699.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[Zynq.scala 49:26:@152700.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[Zynq.scala 49:26:@152701.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[Zynq.scala 49:26:@152702.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[Zynq.scala 49:26:@152703.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[Zynq.scala 49:26:@152704.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[Zynq.scala 49:26:@152705.4]
  assign accel_io_memStreams_stores_0_cmd_ready = FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 49:26:@152689.4]
  assign accel_io_memStreams_stores_0_data_ready = FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 49:26:@152685.4]
  assign accel_io_memStreams_stores_0_wresp_valid = FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 49:26:@152680.4]
  assign accel_io_memStreams_stores_0_wresp_bits = FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 49:26:@152679.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@152678.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@152659.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[Zynq.scala 49:26:@152643.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[Zynq.scala 49:26:@152644.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[Zynq.scala 49:26:@152645.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[Zynq.scala 49:26:@152646.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[Zynq.scala 49:26:@152647.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[Zynq.scala 49:26:@152648.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[Zynq.scala 49:26:@152649.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[Zynq.scala 49:26:@152650.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[Zynq.scala 49:26:@152651.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[Zynq.scala 49:26:@152652.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[Zynq.scala 49:26:@152653.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[Zynq.scala 49:26:@152654.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[Zynq.scala 49:26:@152655.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[Zynq.scala 49:26:@152656.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[Zynq.scala 49:26:@152657.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[Zynq.scala 49:26:@152658.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@152642.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[Zynq.scala 49:26:@152607.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[Zynq.scala 49:26:@152606.4]
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 50:20:@152714.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 50:20:@152713.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 50:20:@152712.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[Zynq.scala 34:21:@152600.4]
  assign accel_io_argIns_1 = FringeZynq_io_argIns_1; // @[Zynq.scala 34:21:@152601.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[Zynq.scala 40:24:@152604.4]
  assign FringeZynq_clock = clock; // @[:@152250.4]
  assign FringeZynq_reset = reset == 1'h0; // @[:@152251.4 Zynq.scala 53:18:@152722.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[Zynq.scala 21:21:@152270.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[Zynq.scala 21:21:@152269.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[Zynq.scala 21:21:@152268.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[Zynq.scala 21:21:@152266.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[Zynq.scala 21:21:@152265.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[Zynq.scala 21:21:@152264.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[Zynq.scala 21:21:@152262.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[Zynq.scala 21:21:@152261.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[Zynq.scala 21:21:@152260.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[Zynq.scala 21:21:@152255.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[Zynq.scala 21:21:@152252.4]
  assign FringeZynq_io_M_AXI_0_AWREADY = io_M_AXI_0_AWREADY; // @[Zynq.scala 24:14:@152300.4]
  assign FringeZynq_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY; // @[Zynq.scala 24:14:@152288.4]
  assign FringeZynq_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY; // @[Zynq.scala 24:14:@152283.4]
  assign FringeZynq_io_M_AXI_0_BID = io_M_AXI_0_BID; // @[Zynq.scala 24:14:@152275.4]
  assign FringeZynq_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID; // @[Zynq.scala 24:14:@152272.4]
  assign FringeZynq_io_M_AXI_1_AWREADY = io_M_AXI_1_AWREADY; // @[Zynq.scala 24:14:@152341.4]
  assign FringeZynq_io_M_AXI_1_ARREADY = io_M_AXI_1_ARREADY; // @[Zynq.scala 24:14:@152329.4]
  assign FringeZynq_io_M_AXI_1_WREADY = io_M_AXI_1_WREADY; // @[Zynq.scala 24:14:@152324.4]
  assign FringeZynq_io_M_AXI_1_BID = io_M_AXI_1_BID; // @[Zynq.scala 24:14:@152316.4]
  assign FringeZynq_io_M_AXI_1_BVALID = io_M_AXI_1_BVALID; // @[Zynq.scala 24:14:@152313.4]
  assign FringeZynq_io_M_AXI_2_AWREADY = io_M_AXI_2_AWREADY; // @[Zynq.scala 24:14:@152382.4]
  assign FringeZynq_io_M_AXI_2_ARREADY = io_M_AXI_2_ARREADY; // @[Zynq.scala 24:14:@152370.4]
  assign FringeZynq_io_M_AXI_2_WREADY = io_M_AXI_2_WREADY; // @[Zynq.scala 24:14:@152365.4]
  assign FringeZynq_io_M_AXI_2_BID = io_M_AXI_2_BID; // @[Zynq.scala 24:14:@152357.4]
  assign FringeZynq_io_M_AXI_2_BVALID = io_M_AXI_2_BVALID; // @[Zynq.scala 24:14:@152354.4]
  assign FringeZynq_io_M_AXI_3_AWREADY = io_M_AXI_3_AWREADY; // @[Zynq.scala 24:14:@152423.4]
  assign FringeZynq_io_M_AXI_3_ARREADY = io_M_AXI_3_ARREADY; // @[Zynq.scala 24:14:@152411.4]
  assign FringeZynq_io_M_AXI_3_WREADY = io_M_AXI_3_WREADY; // @[Zynq.scala 24:14:@152406.4]
  assign FringeZynq_io_M_AXI_3_BID = io_M_AXI_3_BID; // @[Zynq.scala 24:14:@152398.4]
  assign FringeZynq_io_M_AXI_3_BVALID = io_M_AXI_3_BVALID; // @[Zynq.scala 24:14:@152395.4]
  assign FringeZynq_io_done = accel_io_done; // @[Zynq.scala 52:20:@152719.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[Zynq.scala 37:26:@152603.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[Zynq.scala 36:25:@152602.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_valid = accel_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 49:26:@152688.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_addr = accel_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 49:26:@152687.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_size = accel_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 49:26:@152686.4]
  assign FringeZynq_io_memStreams_stores_0_data_valid = accel_io_memStreams_stores_0_data_valid; // @[Zynq.scala 49:26:@152684.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wdata_0 = accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 49:26:@152683.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wstrb = accel_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 49:26:@152682.4]
  assign FringeZynq_io_memStreams_stores_0_wresp_ready = accel_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 49:26:@152681.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[Zynq.scala 50:20:@152717.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 50:20:@152716.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 50:20:@152715.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module SRAMVerilogDualRead
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr0,
    input [AWIDTH-1:0] raddr1,
    input [AWIDTH-1:0] waddr,
    input raddrEn0,
    input raddrEn1,
    input waddrEn,
    input wen,
    input backpressure0,
    input backpressure1,
    input [DWIDTH-1:0] wdata,
    output reg [DWIDTH-1:0] rdata0,
    output reg [DWIDTH-1:0] rdata1
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk)
    begin
            if (wen)
            begin
                mem[waddr] <= wdata;
            end
            if (backpressure0) rdata0 <= mem[raddr0];
    end


    always @(posedge clk)
    begin
        if (backpressure1) rdata1 <= mem[raddr1];
    end
endmodule




