module FIFO(
  input        clock,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_1_0_0,
  input  [7:0] I_2_0_0,
  input  [7:0] I_3_0_0,
  input  [7:0] I_4_0_0,
  input  [7:0] I_5_0_0,
  input  [7:0] I_6_0_0,
  input  [7:0] I_7_0_0,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0
);
  reg [7:0] _T__0_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [7:0] _T__1_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg [7:0] _T__2_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg [7:0] _T__3_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg [7:0] _T__4_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_4;
  reg [7:0] _T__5_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_5;
  reg [7:0] _T__6_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_6;
  reg [7:0] _T__7_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_7;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_8;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0_0_0 = _T__0_0_0; // @[FIFO.scala 14:7]
  assign O_1_0_0 = _T__1_0_0; // @[FIFO.scala 14:7]
  assign O_2_0_0 = _T__2_0_0; // @[FIFO.scala 14:7]
  assign O_3_0_0 = _T__3_0_0; // @[FIFO.scala 14:7]
  assign O_4_0_0 = _T__4_0_0; // @[FIFO.scala 14:7]
  assign O_5_0_0 = _T__5_0_0; // @[FIFO.scala 14:7]
  assign O_6_0_0 = _T__6_0_0; // @[FIFO.scala 14:7]
  assign O_7_0_0 = _T__7_0_0; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0_0_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__1_0_0 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__2_0_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__3_0_0 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T__4_0_0 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T__5_0_0 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__6_0_0 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__7_0_0 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0_0_0 <= I_0_0_0;
    _T__1_0_0 <= I_1_0_0;
    _T__2_0_0 <= I_2_0_0;
    _T__3_0_0 <= I_3_0_0;
    _T__4_0_0 <= I_4_0_0;
    _T__5_0_0 <= I_5_0_0;
    _T__6_0_0 <= I_6_0_0;
    _T__7_0_0 <= I_7_0_0;
    _T_1 <= valid_up;
  end
endmodule
module NestedCounters(
  input   CE,
  output  valid
);
  assign valid = CE; // @[NestedCounters.scala 65:13]
endmodule
module NestedCounters_1(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 53:31]
  wire  NestedCounters_valid; // @[NestedCounters.scala 53:31]
  NestedCounters NestedCounters ( // @[NestedCounters.scala 53:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 56:11]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 57:22]
endmodule
module NestedCounters_2(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 53:31]
  wire  NestedCounters_valid; // @[NestedCounters.scala 53:31]
  NestedCounters_1 NestedCounters ( // @[NestedCounters.scala 53:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 56:11]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 57:22]
endmodule
module NestedCountersWithNumValid(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 20:44]
  wire  NestedCounters_valid; // @[NestedCounters.scala 20:44]
  NestedCounters_2 NestedCounters ( // @[NestedCounters.scala 20:44]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 22:9]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 21:27]
endmodule
module RAM_ST(
  input        clock,
  input        RE,
  input  [7:0] RADDR,
  output [7:0] RDATA_0_0,
  input        WE,
  input  [7:0] WADDR,
  input  [7:0] WDATA_0_0
);
  wire  write_elem_counter_CE; // @[RAM_ST.scala 20:34]
  wire  write_elem_counter_valid; // @[RAM_ST.scala 20:34]
  wire  read_elem_counter_CE; // @[RAM_ST.scala 21:33]
  wire  read_elem_counter_valid; // @[RAM_ST.scala 21:33]
  reg [7:0] ram_0_0 [0:239]; // @[RAM_ST.scala 29:24]
  reg [31:0] _RAND_0;
  wire [7:0] ram_0_0__T_8_data; // @[RAM_ST.scala 29:24]
  wire [7:0] ram_0_0__T_8_addr; // @[RAM_ST.scala 29:24]
  reg [31:0] _RAND_1;
  wire [7:0] ram_0_0__T_2_data; // @[RAM_ST.scala 29:24]
  wire [7:0] ram_0_0__T_2_addr; // @[RAM_ST.scala 29:24]
  wire  ram_0_0__T_2_mask; // @[RAM_ST.scala 29:24]
  wire  ram_0_0__T_2_en; // @[RAM_ST.scala 29:24]
  reg  ram_0_0__T_8_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [7:0] ram_0_0__T_8_addr_pipe_0;
  reg [31:0] _RAND_3;
  wire [7:0] _GEN_1; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_2; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_3; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_4; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_5; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_6; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_7; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_8; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_9; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_10; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_11; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_12; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_13; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_14; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_15; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_16; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_17; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_18; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_19; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_20; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_21; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_22; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_23; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_24; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_25; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_26; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_27; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_28; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_29; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_30; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_31; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_32; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_33; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_34; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_35; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_36; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_37; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_38; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_39; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_40; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_41; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_42; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_43; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_44; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_45; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_46; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_47; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_48; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_49; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_50; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_51; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_52; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_53; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_54; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_55; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_56; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_57; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_58; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_59; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_60; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_61; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_62; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_63; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_64; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_65; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_66; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_67; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_68; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_69; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_70; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_71; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_72; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_73; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_74; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_75; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_76; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_77; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_78; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_79; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_80; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_81; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_82; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_83; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_84; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_85; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_86; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_87; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_88; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_89; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_90; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_91; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_92; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_93; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_94; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_95; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_96; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_97; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_98; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_99; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_100; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_101; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_102; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_103; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_104; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_105; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_106; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_107; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_108; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_109; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_110; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_111; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_112; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_113; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_114; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_115; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_116; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_117; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_118; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_119; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_120; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_121; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_122; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_123; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_124; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_125; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_126; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_127; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_128; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_129; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_130; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_131; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_132; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_133; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_134; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_135; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_136; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_137; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_138; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_139; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_140; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_141; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_142; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_143; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_144; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_145; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_146; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_147; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_148; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_149; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_150; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_151; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_152; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_153; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_154; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_155; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_156; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_157; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_158; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_159; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_160; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_161; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_162; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_163; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_164; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_165; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_166; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_167; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_168; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_169; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_170; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_171; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_172; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_173; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_174; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_175; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_176; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_177; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_178; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_179; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_180; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_181; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_182; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_183; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_184; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_185; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_186; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_187; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_188; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_189; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_190; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_191; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_192; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_193; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_194; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_195; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_196; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_197; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_198; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_199; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_200; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_201; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_202; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_203; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_204; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_205; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_206; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_207; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_208; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_209; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_210; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_211; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_212; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_213; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_214; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_215; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_216; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_217; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_218; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_219; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_220; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_221; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_222; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_223; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_224; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_225; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_226; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_227; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_228; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_229; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_230; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_231; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_232; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_233; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_234; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_235; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_236; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_237; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_238; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_239; // @[RAM_ST.scala 31:71]
  wire [8:0] _T; // @[RAM_ST.scala 31:71]
  wire [7:0] _GEN_246; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_247; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_248; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_249; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_250; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_251; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_252; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_253; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_254; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_255; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_256; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_257; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_258; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_259; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_260; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_261; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_262; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_263; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_264; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_265; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_266; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_267; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_268; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_269; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_270; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_271; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_272; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_273; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_274; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_275; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_276; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_277; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_278; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_279; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_280; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_281; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_282; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_283; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_284; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_285; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_286; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_287; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_288; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_289; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_290; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_291; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_292; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_293; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_294; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_295; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_296; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_297; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_298; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_299; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_300; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_301; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_302; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_303; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_304; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_305; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_306; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_307; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_308; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_309; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_310; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_311; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_312; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_313; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_314; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_315; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_316; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_317; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_318; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_319; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_320; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_321; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_322; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_323; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_324; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_325; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_326; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_327; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_328; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_329; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_330; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_331; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_332; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_333; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_334; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_335; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_336; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_337; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_338; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_339; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_340; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_341; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_342; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_343; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_344; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_345; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_346; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_347; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_348; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_349; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_350; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_351; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_352; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_353; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_354; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_355; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_356; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_357; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_358; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_359; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_360; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_361; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_362; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_363; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_364; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_365; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_366; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_367; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_368; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_369; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_370; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_371; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_372; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_373; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_374; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_375; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_376; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_377; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_378; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_379; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_380; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_381; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_382; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_383; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_384; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_385; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_386; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_387; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_388; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_389; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_390; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_391; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_392; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_393; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_394; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_395; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_396; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_397; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_398; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_399; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_400; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_401; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_402; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_403; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_404; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_405; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_406; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_407; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_408; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_409; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_410; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_411; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_412; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_413; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_414; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_415; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_416; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_417; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_418; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_419; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_420; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_421; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_422; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_423; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_424; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_425; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_426; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_427; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_428; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_429; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_430; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_431; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_432; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_433; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_434; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_435; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_436; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_437; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_438; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_439; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_440; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_441; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_442; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_443; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_444; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_445; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_446; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_447; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_448; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_449; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_450; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_451; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_452; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_453; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_454; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_455; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_456; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_457; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_458; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_459; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_460; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_461; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_462; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_463; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_464; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_465; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_466; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_467; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_468; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_469; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_470; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_471; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_472; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_473; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_474; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_475; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_476; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_477; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_478; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_479; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_480; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_481; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_482; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_483; // @[RAM_ST.scala 32:46]
  wire [7:0] _GEN_484; // @[RAM_ST.scala 32:46]
  wire [8:0] _T_3; // @[RAM_ST.scala 32:46]
  NestedCountersWithNumValid write_elem_counter ( // @[RAM_ST.scala 20:34]
    .CE(write_elem_counter_CE),
    .valid(write_elem_counter_valid)
  );
  NestedCountersWithNumValid read_elem_counter ( // @[RAM_ST.scala 21:33]
    .CE(read_elem_counter_CE),
    .valid(read_elem_counter_valid)
  );
  assign ram_0_0__T_8_addr = ram_0_0__T_8_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_0_0__T_8_data = ram_0_0[ram_0_0__T_8_addr]; // @[RAM_ST.scala 29:24]
  `else
  assign ram_0_0__T_8_data = ram_0_0__T_8_addr >= 8'hf0 ? _RAND_1[7:0] : ram_0_0[ram_0_0__T_8_addr]; // @[RAM_ST.scala 29:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_0_0__T_2_data = WDATA_0_0;
  assign ram_0_0__T_2_addr = _T[7:0];
  assign ram_0_0__T_2_mask = 1'h1;
  assign ram_0_0__T_2_en = write_elem_counter_valid;
  assign _GEN_1 = 8'h1 == WADDR ? 8'h1 : 8'h0; // @[RAM_ST.scala 31:71]
  assign _GEN_2 = 8'h2 == WADDR ? 8'h2 : _GEN_1; // @[RAM_ST.scala 31:71]
  assign _GEN_3 = 8'h3 == WADDR ? 8'h3 : _GEN_2; // @[RAM_ST.scala 31:71]
  assign _GEN_4 = 8'h4 == WADDR ? 8'h4 : _GEN_3; // @[RAM_ST.scala 31:71]
  assign _GEN_5 = 8'h5 == WADDR ? 8'h5 : _GEN_4; // @[RAM_ST.scala 31:71]
  assign _GEN_6 = 8'h6 == WADDR ? 8'h6 : _GEN_5; // @[RAM_ST.scala 31:71]
  assign _GEN_7 = 8'h7 == WADDR ? 8'h7 : _GEN_6; // @[RAM_ST.scala 31:71]
  assign _GEN_8 = 8'h8 == WADDR ? 8'h8 : _GEN_7; // @[RAM_ST.scala 31:71]
  assign _GEN_9 = 8'h9 == WADDR ? 8'h9 : _GEN_8; // @[RAM_ST.scala 31:71]
  assign _GEN_10 = 8'ha == WADDR ? 8'ha : _GEN_9; // @[RAM_ST.scala 31:71]
  assign _GEN_11 = 8'hb == WADDR ? 8'hb : _GEN_10; // @[RAM_ST.scala 31:71]
  assign _GEN_12 = 8'hc == WADDR ? 8'hc : _GEN_11; // @[RAM_ST.scala 31:71]
  assign _GEN_13 = 8'hd == WADDR ? 8'hd : _GEN_12; // @[RAM_ST.scala 31:71]
  assign _GEN_14 = 8'he == WADDR ? 8'he : _GEN_13; // @[RAM_ST.scala 31:71]
  assign _GEN_15 = 8'hf == WADDR ? 8'hf : _GEN_14; // @[RAM_ST.scala 31:71]
  assign _GEN_16 = 8'h10 == WADDR ? 8'h10 : _GEN_15; // @[RAM_ST.scala 31:71]
  assign _GEN_17 = 8'h11 == WADDR ? 8'h11 : _GEN_16; // @[RAM_ST.scala 31:71]
  assign _GEN_18 = 8'h12 == WADDR ? 8'h12 : _GEN_17; // @[RAM_ST.scala 31:71]
  assign _GEN_19 = 8'h13 == WADDR ? 8'h13 : _GEN_18; // @[RAM_ST.scala 31:71]
  assign _GEN_20 = 8'h14 == WADDR ? 8'h14 : _GEN_19; // @[RAM_ST.scala 31:71]
  assign _GEN_21 = 8'h15 == WADDR ? 8'h15 : _GEN_20; // @[RAM_ST.scala 31:71]
  assign _GEN_22 = 8'h16 == WADDR ? 8'h16 : _GEN_21; // @[RAM_ST.scala 31:71]
  assign _GEN_23 = 8'h17 == WADDR ? 8'h17 : _GEN_22; // @[RAM_ST.scala 31:71]
  assign _GEN_24 = 8'h18 == WADDR ? 8'h18 : _GEN_23; // @[RAM_ST.scala 31:71]
  assign _GEN_25 = 8'h19 == WADDR ? 8'h19 : _GEN_24; // @[RAM_ST.scala 31:71]
  assign _GEN_26 = 8'h1a == WADDR ? 8'h1a : _GEN_25; // @[RAM_ST.scala 31:71]
  assign _GEN_27 = 8'h1b == WADDR ? 8'h1b : _GEN_26; // @[RAM_ST.scala 31:71]
  assign _GEN_28 = 8'h1c == WADDR ? 8'h1c : _GEN_27; // @[RAM_ST.scala 31:71]
  assign _GEN_29 = 8'h1d == WADDR ? 8'h1d : _GEN_28; // @[RAM_ST.scala 31:71]
  assign _GEN_30 = 8'h1e == WADDR ? 8'h1e : _GEN_29; // @[RAM_ST.scala 31:71]
  assign _GEN_31 = 8'h1f == WADDR ? 8'h1f : _GEN_30; // @[RAM_ST.scala 31:71]
  assign _GEN_32 = 8'h20 == WADDR ? 8'h20 : _GEN_31; // @[RAM_ST.scala 31:71]
  assign _GEN_33 = 8'h21 == WADDR ? 8'h21 : _GEN_32; // @[RAM_ST.scala 31:71]
  assign _GEN_34 = 8'h22 == WADDR ? 8'h22 : _GEN_33; // @[RAM_ST.scala 31:71]
  assign _GEN_35 = 8'h23 == WADDR ? 8'h23 : _GEN_34; // @[RAM_ST.scala 31:71]
  assign _GEN_36 = 8'h24 == WADDR ? 8'h24 : _GEN_35; // @[RAM_ST.scala 31:71]
  assign _GEN_37 = 8'h25 == WADDR ? 8'h25 : _GEN_36; // @[RAM_ST.scala 31:71]
  assign _GEN_38 = 8'h26 == WADDR ? 8'h26 : _GEN_37; // @[RAM_ST.scala 31:71]
  assign _GEN_39 = 8'h27 == WADDR ? 8'h27 : _GEN_38; // @[RAM_ST.scala 31:71]
  assign _GEN_40 = 8'h28 == WADDR ? 8'h28 : _GEN_39; // @[RAM_ST.scala 31:71]
  assign _GEN_41 = 8'h29 == WADDR ? 8'h29 : _GEN_40; // @[RAM_ST.scala 31:71]
  assign _GEN_42 = 8'h2a == WADDR ? 8'h2a : _GEN_41; // @[RAM_ST.scala 31:71]
  assign _GEN_43 = 8'h2b == WADDR ? 8'h2b : _GEN_42; // @[RAM_ST.scala 31:71]
  assign _GEN_44 = 8'h2c == WADDR ? 8'h2c : _GEN_43; // @[RAM_ST.scala 31:71]
  assign _GEN_45 = 8'h2d == WADDR ? 8'h2d : _GEN_44; // @[RAM_ST.scala 31:71]
  assign _GEN_46 = 8'h2e == WADDR ? 8'h2e : _GEN_45; // @[RAM_ST.scala 31:71]
  assign _GEN_47 = 8'h2f == WADDR ? 8'h2f : _GEN_46; // @[RAM_ST.scala 31:71]
  assign _GEN_48 = 8'h30 == WADDR ? 8'h30 : _GEN_47; // @[RAM_ST.scala 31:71]
  assign _GEN_49 = 8'h31 == WADDR ? 8'h31 : _GEN_48; // @[RAM_ST.scala 31:71]
  assign _GEN_50 = 8'h32 == WADDR ? 8'h32 : _GEN_49; // @[RAM_ST.scala 31:71]
  assign _GEN_51 = 8'h33 == WADDR ? 8'h33 : _GEN_50; // @[RAM_ST.scala 31:71]
  assign _GEN_52 = 8'h34 == WADDR ? 8'h34 : _GEN_51; // @[RAM_ST.scala 31:71]
  assign _GEN_53 = 8'h35 == WADDR ? 8'h35 : _GEN_52; // @[RAM_ST.scala 31:71]
  assign _GEN_54 = 8'h36 == WADDR ? 8'h36 : _GEN_53; // @[RAM_ST.scala 31:71]
  assign _GEN_55 = 8'h37 == WADDR ? 8'h37 : _GEN_54; // @[RAM_ST.scala 31:71]
  assign _GEN_56 = 8'h38 == WADDR ? 8'h38 : _GEN_55; // @[RAM_ST.scala 31:71]
  assign _GEN_57 = 8'h39 == WADDR ? 8'h39 : _GEN_56; // @[RAM_ST.scala 31:71]
  assign _GEN_58 = 8'h3a == WADDR ? 8'h3a : _GEN_57; // @[RAM_ST.scala 31:71]
  assign _GEN_59 = 8'h3b == WADDR ? 8'h3b : _GEN_58; // @[RAM_ST.scala 31:71]
  assign _GEN_60 = 8'h3c == WADDR ? 8'h3c : _GEN_59; // @[RAM_ST.scala 31:71]
  assign _GEN_61 = 8'h3d == WADDR ? 8'h3d : _GEN_60; // @[RAM_ST.scala 31:71]
  assign _GEN_62 = 8'h3e == WADDR ? 8'h3e : _GEN_61; // @[RAM_ST.scala 31:71]
  assign _GEN_63 = 8'h3f == WADDR ? 8'h3f : _GEN_62; // @[RAM_ST.scala 31:71]
  assign _GEN_64 = 8'h40 == WADDR ? 8'h40 : _GEN_63; // @[RAM_ST.scala 31:71]
  assign _GEN_65 = 8'h41 == WADDR ? 8'h41 : _GEN_64; // @[RAM_ST.scala 31:71]
  assign _GEN_66 = 8'h42 == WADDR ? 8'h42 : _GEN_65; // @[RAM_ST.scala 31:71]
  assign _GEN_67 = 8'h43 == WADDR ? 8'h43 : _GEN_66; // @[RAM_ST.scala 31:71]
  assign _GEN_68 = 8'h44 == WADDR ? 8'h44 : _GEN_67; // @[RAM_ST.scala 31:71]
  assign _GEN_69 = 8'h45 == WADDR ? 8'h45 : _GEN_68; // @[RAM_ST.scala 31:71]
  assign _GEN_70 = 8'h46 == WADDR ? 8'h46 : _GEN_69; // @[RAM_ST.scala 31:71]
  assign _GEN_71 = 8'h47 == WADDR ? 8'h47 : _GEN_70; // @[RAM_ST.scala 31:71]
  assign _GEN_72 = 8'h48 == WADDR ? 8'h48 : _GEN_71; // @[RAM_ST.scala 31:71]
  assign _GEN_73 = 8'h49 == WADDR ? 8'h49 : _GEN_72; // @[RAM_ST.scala 31:71]
  assign _GEN_74 = 8'h4a == WADDR ? 8'h4a : _GEN_73; // @[RAM_ST.scala 31:71]
  assign _GEN_75 = 8'h4b == WADDR ? 8'h4b : _GEN_74; // @[RAM_ST.scala 31:71]
  assign _GEN_76 = 8'h4c == WADDR ? 8'h4c : _GEN_75; // @[RAM_ST.scala 31:71]
  assign _GEN_77 = 8'h4d == WADDR ? 8'h4d : _GEN_76; // @[RAM_ST.scala 31:71]
  assign _GEN_78 = 8'h4e == WADDR ? 8'h4e : _GEN_77; // @[RAM_ST.scala 31:71]
  assign _GEN_79 = 8'h4f == WADDR ? 8'h4f : _GEN_78; // @[RAM_ST.scala 31:71]
  assign _GEN_80 = 8'h50 == WADDR ? 8'h50 : _GEN_79; // @[RAM_ST.scala 31:71]
  assign _GEN_81 = 8'h51 == WADDR ? 8'h51 : _GEN_80; // @[RAM_ST.scala 31:71]
  assign _GEN_82 = 8'h52 == WADDR ? 8'h52 : _GEN_81; // @[RAM_ST.scala 31:71]
  assign _GEN_83 = 8'h53 == WADDR ? 8'h53 : _GEN_82; // @[RAM_ST.scala 31:71]
  assign _GEN_84 = 8'h54 == WADDR ? 8'h54 : _GEN_83; // @[RAM_ST.scala 31:71]
  assign _GEN_85 = 8'h55 == WADDR ? 8'h55 : _GEN_84; // @[RAM_ST.scala 31:71]
  assign _GEN_86 = 8'h56 == WADDR ? 8'h56 : _GEN_85; // @[RAM_ST.scala 31:71]
  assign _GEN_87 = 8'h57 == WADDR ? 8'h57 : _GEN_86; // @[RAM_ST.scala 31:71]
  assign _GEN_88 = 8'h58 == WADDR ? 8'h58 : _GEN_87; // @[RAM_ST.scala 31:71]
  assign _GEN_89 = 8'h59 == WADDR ? 8'h59 : _GEN_88; // @[RAM_ST.scala 31:71]
  assign _GEN_90 = 8'h5a == WADDR ? 8'h5a : _GEN_89; // @[RAM_ST.scala 31:71]
  assign _GEN_91 = 8'h5b == WADDR ? 8'h5b : _GEN_90; // @[RAM_ST.scala 31:71]
  assign _GEN_92 = 8'h5c == WADDR ? 8'h5c : _GEN_91; // @[RAM_ST.scala 31:71]
  assign _GEN_93 = 8'h5d == WADDR ? 8'h5d : _GEN_92; // @[RAM_ST.scala 31:71]
  assign _GEN_94 = 8'h5e == WADDR ? 8'h5e : _GEN_93; // @[RAM_ST.scala 31:71]
  assign _GEN_95 = 8'h5f == WADDR ? 8'h5f : _GEN_94; // @[RAM_ST.scala 31:71]
  assign _GEN_96 = 8'h60 == WADDR ? 8'h60 : _GEN_95; // @[RAM_ST.scala 31:71]
  assign _GEN_97 = 8'h61 == WADDR ? 8'h61 : _GEN_96; // @[RAM_ST.scala 31:71]
  assign _GEN_98 = 8'h62 == WADDR ? 8'h62 : _GEN_97; // @[RAM_ST.scala 31:71]
  assign _GEN_99 = 8'h63 == WADDR ? 8'h63 : _GEN_98; // @[RAM_ST.scala 31:71]
  assign _GEN_100 = 8'h64 == WADDR ? 8'h64 : _GEN_99; // @[RAM_ST.scala 31:71]
  assign _GEN_101 = 8'h65 == WADDR ? 8'h65 : _GEN_100; // @[RAM_ST.scala 31:71]
  assign _GEN_102 = 8'h66 == WADDR ? 8'h66 : _GEN_101; // @[RAM_ST.scala 31:71]
  assign _GEN_103 = 8'h67 == WADDR ? 8'h67 : _GEN_102; // @[RAM_ST.scala 31:71]
  assign _GEN_104 = 8'h68 == WADDR ? 8'h68 : _GEN_103; // @[RAM_ST.scala 31:71]
  assign _GEN_105 = 8'h69 == WADDR ? 8'h69 : _GEN_104; // @[RAM_ST.scala 31:71]
  assign _GEN_106 = 8'h6a == WADDR ? 8'h6a : _GEN_105; // @[RAM_ST.scala 31:71]
  assign _GEN_107 = 8'h6b == WADDR ? 8'h6b : _GEN_106; // @[RAM_ST.scala 31:71]
  assign _GEN_108 = 8'h6c == WADDR ? 8'h6c : _GEN_107; // @[RAM_ST.scala 31:71]
  assign _GEN_109 = 8'h6d == WADDR ? 8'h6d : _GEN_108; // @[RAM_ST.scala 31:71]
  assign _GEN_110 = 8'h6e == WADDR ? 8'h6e : _GEN_109; // @[RAM_ST.scala 31:71]
  assign _GEN_111 = 8'h6f == WADDR ? 8'h6f : _GEN_110; // @[RAM_ST.scala 31:71]
  assign _GEN_112 = 8'h70 == WADDR ? 8'h70 : _GEN_111; // @[RAM_ST.scala 31:71]
  assign _GEN_113 = 8'h71 == WADDR ? 8'h71 : _GEN_112; // @[RAM_ST.scala 31:71]
  assign _GEN_114 = 8'h72 == WADDR ? 8'h72 : _GEN_113; // @[RAM_ST.scala 31:71]
  assign _GEN_115 = 8'h73 == WADDR ? 8'h73 : _GEN_114; // @[RAM_ST.scala 31:71]
  assign _GEN_116 = 8'h74 == WADDR ? 8'h74 : _GEN_115; // @[RAM_ST.scala 31:71]
  assign _GEN_117 = 8'h75 == WADDR ? 8'h75 : _GEN_116; // @[RAM_ST.scala 31:71]
  assign _GEN_118 = 8'h76 == WADDR ? 8'h76 : _GEN_117; // @[RAM_ST.scala 31:71]
  assign _GEN_119 = 8'h77 == WADDR ? 8'h77 : _GEN_118; // @[RAM_ST.scala 31:71]
  assign _GEN_120 = 8'h78 == WADDR ? 8'h78 : _GEN_119; // @[RAM_ST.scala 31:71]
  assign _GEN_121 = 8'h79 == WADDR ? 8'h79 : _GEN_120; // @[RAM_ST.scala 31:71]
  assign _GEN_122 = 8'h7a == WADDR ? 8'h7a : _GEN_121; // @[RAM_ST.scala 31:71]
  assign _GEN_123 = 8'h7b == WADDR ? 8'h7b : _GEN_122; // @[RAM_ST.scala 31:71]
  assign _GEN_124 = 8'h7c == WADDR ? 8'h7c : _GEN_123; // @[RAM_ST.scala 31:71]
  assign _GEN_125 = 8'h7d == WADDR ? 8'h7d : _GEN_124; // @[RAM_ST.scala 31:71]
  assign _GEN_126 = 8'h7e == WADDR ? 8'h7e : _GEN_125; // @[RAM_ST.scala 31:71]
  assign _GEN_127 = 8'h7f == WADDR ? 8'h7f : _GEN_126; // @[RAM_ST.scala 31:71]
  assign _GEN_128 = 8'h80 == WADDR ? 8'h80 : _GEN_127; // @[RAM_ST.scala 31:71]
  assign _GEN_129 = 8'h81 == WADDR ? 8'h81 : _GEN_128; // @[RAM_ST.scala 31:71]
  assign _GEN_130 = 8'h82 == WADDR ? 8'h82 : _GEN_129; // @[RAM_ST.scala 31:71]
  assign _GEN_131 = 8'h83 == WADDR ? 8'h83 : _GEN_130; // @[RAM_ST.scala 31:71]
  assign _GEN_132 = 8'h84 == WADDR ? 8'h84 : _GEN_131; // @[RAM_ST.scala 31:71]
  assign _GEN_133 = 8'h85 == WADDR ? 8'h85 : _GEN_132; // @[RAM_ST.scala 31:71]
  assign _GEN_134 = 8'h86 == WADDR ? 8'h86 : _GEN_133; // @[RAM_ST.scala 31:71]
  assign _GEN_135 = 8'h87 == WADDR ? 8'h87 : _GEN_134; // @[RAM_ST.scala 31:71]
  assign _GEN_136 = 8'h88 == WADDR ? 8'h88 : _GEN_135; // @[RAM_ST.scala 31:71]
  assign _GEN_137 = 8'h89 == WADDR ? 8'h89 : _GEN_136; // @[RAM_ST.scala 31:71]
  assign _GEN_138 = 8'h8a == WADDR ? 8'h8a : _GEN_137; // @[RAM_ST.scala 31:71]
  assign _GEN_139 = 8'h8b == WADDR ? 8'h8b : _GEN_138; // @[RAM_ST.scala 31:71]
  assign _GEN_140 = 8'h8c == WADDR ? 8'h8c : _GEN_139; // @[RAM_ST.scala 31:71]
  assign _GEN_141 = 8'h8d == WADDR ? 8'h8d : _GEN_140; // @[RAM_ST.scala 31:71]
  assign _GEN_142 = 8'h8e == WADDR ? 8'h8e : _GEN_141; // @[RAM_ST.scala 31:71]
  assign _GEN_143 = 8'h8f == WADDR ? 8'h8f : _GEN_142; // @[RAM_ST.scala 31:71]
  assign _GEN_144 = 8'h90 == WADDR ? 8'h90 : _GEN_143; // @[RAM_ST.scala 31:71]
  assign _GEN_145 = 8'h91 == WADDR ? 8'h91 : _GEN_144; // @[RAM_ST.scala 31:71]
  assign _GEN_146 = 8'h92 == WADDR ? 8'h92 : _GEN_145; // @[RAM_ST.scala 31:71]
  assign _GEN_147 = 8'h93 == WADDR ? 8'h93 : _GEN_146; // @[RAM_ST.scala 31:71]
  assign _GEN_148 = 8'h94 == WADDR ? 8'h94 : _GEN_147; // @[RAM_ST.scala 31:71]
  assign _GEN_149 = 8'h95 == WADDR ? 8'h95 : _GEN_148; // @[RAM_ST.scala 31:71]
  assign _GEN_150 = 8'h96 == WADDR ? 8'h96 : _GEN_149; // @[RAM_ST.scala 31:71]
  assign _GEN_151 = 8'h97 == WADDR ? 8'h97 : _GEN_150; // @[RAM_ST.scala 31:71]
  assign _GEN_152 = 8'h98 == WADDR ? 8'h98 : _GEN_151; // @[RAM_ST.scala 31:71]
  assign _GEN_153 = 8'h99 == WADDR ? 8'h99 : _GEN_152; // @[RAM_ST.scala 31:71]
  assign _GEN_154 = 8'h9a == WADDR ? 8'h9a : _GEN_153; // @[RAM_ST.scala 31:71]
  assign _GEN_155 = 8'h9b == WADDR ? 8'h9b : _GEN_154; // @[RAM_ST.scala 31:71]
  assign _GEN_156 = 8'h9c == WADDR ? 8'h9c : _GEN_155; // @[RAM_ST.scala 31:71]
  assign _GEN_157 = 8'h9d == WADDR ? 8'h9d : _GEN_156; // @[RAM_ST.scala 31:71]
  assign _GEN_158 = 8'h9e == WADDR ? 8'h9e : _GEN_157; // @[RAM_ST.scala 31:71]
  assign _GEN_159 = 8'h9f == WADDR ? 8'h9f : _GEN_158; // @[RAM_ST.scala 31:71]
  assign _GEN_160 = 8'ha0 == WADDR ? 8'ha0 : _GEN_159; // @[RAM_ST.scala 31:71]
  assign _GEN_161 = 8'ha1 == WADDR ? 8'ha1 : _GEN_160; // @[RAM_ST.scala 31:71]
  assign _GEN_162 = 8'ha2 == WADDR ? 8'ha2 : _GEN_161; // @[RAM_ST.scala 31:71]
  assign _GEN_163 = 8'ha3 == WADDR ? 8'ha3 : _GEN_162; // @[RAM_ST.scala 31:71]
  assign _GEN_164 = 8'ha4 == WADDR ? 8'ha4 : _GEN_163; // @[RAM_ST.scala 31:71]
  assign _GEN_165 = 8'ha5 == WADDR ? 8'ha5 : _GEN_164; // @[RAM_ST.scala 31:71]
  assign _GEN_166 = 8'ha6 == WADDR ? 8'ha6 : _GEN_165; // @[RAM_ST.scala 31:71]
  assign _GEN_167 = 8'ha7 == WADDR ? 8'ha7 : _GEN_166; // @[RAM_ST.scala 31:71]
  assign _GEN_168 = 8'ha8 == WADDR ? 8'ha8 : _GEN_167; // @[RAM_ST.scala 31:71]
  assign _GEN_169 = 8'ha9 == WADDR ? 8'ha9 : _GEN_168; // @[RAM_ST.scala 31:71]
  assign _GEN_170 = 8'haa == WADDR ? 8'haa : _GEN_169; // @[RAM_ST.scala 31:71]
  assign _GEN_171 = 8'hab == WADDR ? 8'hab : _GEN_170; // @[RAM_ST.scala 31:71]
  assign _GEN_172 = 8'hac == WADDR ? 8'hac : _GEN_171; // @[RAM_ST.scala 31:71]
  assign _GEN_173 = 8'had == WADDR ? 8'had : _GEN_172; // @[RAM_ST.scala 31:71]
  assign _GEN_174 = 8'hae == WADDR ? 8'hae : _GEN_173; // @[RAM_ST.scala 31:71]
  assign _GEN_175 = 8'haf == WADDR ? 8'haf : _GEN_174; // @[RAM_ST.scala 31:71]
  assign _GEN_176 = 8'hb0 == WADDR ? 8'hb0 : _GEN_175; // @[RAM_ST.scala 31:71]
  assign _GEN_177 = 8'hb1 == WADDR ? 8'hb1 : _GEN_176; // @[RAM_ST.scala 31:71]
  assign _GEN_178 = 8'hb2 == WADDR ? 8'hb2 : _GEN_177; // @[RAM_ST.scala 31:71]
  assign _GEN_179 = 8'hb3 == WADDR ? 8'hb3 : _GEN_178; // @[RAM_ST.scala 31:71]
  assign _GEN_180 = 8'hb4 == WADDR ? 8'hb4 : _GEN_179; // @[RAM_ST.scala 31:71]
  assign _GEN_181 = 8'hb5 == WADDR ? 8'hb5 : _GEN_180; // @[RAM_ST.scala 31:71]
  assign _GEN_182 = 8'hb6 == WADDR ? 8'hb6 : _GEN_181; // @[RAM_ST.scala 31:71]
  assign _GEN_183 = 8'hb7 == WADDR ? 8'hb7 : _GEN_182; // @[RAM_ST.scala 31:71]
  assign _GEN_184 = 8'hb8 == WADDR ? 8'hb8 : _GEN_183; // @[RAM_ST.scala 31:71]
  assign _GEN_185 = 8'hb9 == WADDR ? 8'hb9 : _GEN_184; // @[RAM_ST.scala 31:71]
  assign _GEN_186 = 8'hba == WADDR ? 8'hba : _GEN_185; // @[RAM_ST.scala 31:71]
  assign _GEN_187 = 8'hbb == WADDR ? 8'hbb : _GEN_186; // @[RAM_ST.scala 31:71]
  assign _GEN_188 = 8'hbc == WADDR ? 8'hbc : _GEN_187; // @[RAM_ST.scala 31:71]
  assign _GEN_189 = 8'hbd == WADDR ? 8'hbd : _GEN_188; // @[RAM_ST.scala 31:71]
  assign _GEN_190 = 8'hbe == WADDR ? 8'hbe : _GEN_189; // @[RAM_ST.scala 31:71]
  assign _GEN_191 = 8'hbf == WADDR ? 8'hbf : _GEN_190; // @[RAM_ST.scala 31:71]
  assign _GEN_192 = 8'hc0 == WADDR ? 8'hc0 : _GEN_191; // @[RAM_ST.scala 31:71]
  assign _GEN_193 = 8'hc1 == WADDR ? 8'hc1 : _GEN_192; // @[RAM_ST.scala 31:71]
  assign _GEN_194 = 8'hc2 == WADDR ? 8'hc2 : _GEN_193; // @[RAM_ST.scala 31:71]
  assign _GEN_195 = 8'hc3 == WADDR ? 8'hc3 : _GEN_194; // @[RAM_ST.scala 31:71]
  assign _GEN_196 = 8'hc4 == WADDR ? 8'hc4 : _GEN_195; // @[RAM_ST.scala 31:71]
  assign _GEN_197 = 8'hc5 == WADDR ? 8'hc5 : _GEN_196; // @[RAM_ST.scala 31:71]
  assign _GEN_198 = 8'hc6 == WADDR ? 8'hc6 : _GEN_197; // @[RAM_ST.scala 31:71]
  assign _GEN_199 = 8'hc7 == WADDR ? 8'hc7 : _GEN_198; // @[RAM_ST.scala 31:71]
  assign _GEN_200 = 8'hc8 == WADDR ? 8'hc8 : _GEN_199; // @[RAM_ST.scala 31:71]
  assign _GEN_201 = 8'hc9 == WADDR ? 8'hc9 : _GEN_200; // @[RAM_ST.scala 31:71]
  assign _GEN_202 = 8'hca == WADDR ? 8'hca : _GEN_201; // @[RAM_ST.scala 31:71]
  assign _GEN_203 = 8'hcb == WADDR ? 8'hcb : _GEN_202; // @[RAM_ST.scala 31:71]
  assign _GEN_204 = 8'hcc == WADDR ? 8'hcc : _GEN_203; // @[RAM_ST.scala 31:71]
  assign _GEN_205 = 8'hcd == WADDR ? 8'hcd : _GEN_204; // @[RAM_ST.scala 31:71]
  assign _GEN_206 = 8'hce == WADDR ? 8'hce : _GEN_205; // @[RAM_ST.scala 31:71]
  assign _GEN_207 = 8'hcf == WADDR ? 8'hcf : _GEN_206; // @[RAM_ST.scala 31:71]
  assign _GEN_208 = 8'hd0 == WADDR ? 8'hd0 : _GEN_207; // @[RAM_ST.scala 31:71]
  assign _GEN_209 = 8'hd1 == WADDR ? 8'hd1 : _GEN_208; // @[RAM_ST.scala 31:71]
  assign _GEN_210 = 8'hd2 == WADDR ? 8'hd2 : _GEN_209; // @[RAM_ST.scala 31:71]
  assign _GEN_211 = 8'hd3 == WADDR ? 8'hd3 : _GEN_210; // @[RAM_ST.scala 31:71]
  assign _GEN_212 = 8'hd4 == WADDR ? 8'hd4 : _GEN_211; // @[RAM_ST.scala 31:71]
  assign _GEN_213 = 8'hd5 == WADDR ? 8'hd5 : _GEN_212; // @[RAM_ST.scala 31:71]
  assign _GEN_214 = 8'hd6 == WADDR ? 8'hd6 : _GEN_213; // @[RAM_ST.scala 31:71]
  assign _GEN_215 = 8'hd7 == WADDR ? 8'hd7 : _GEN_214; // @[RAM_ST.scala 31:71]
  assign _GEN_216 = 8'hd8 == WADDR ? 8'hd8 : _GEN_215; // @[RAM_ST.scala 31:71]
  assign _GEN_217 = 8'hd9 == WADDR ? 8'hd9 : _GEN_216; // @[RAM_ST.scala 31:71]
  assign _GEN_218 = 8'hda == WADDR ? 8'hda : _GEN_217; // @[RAM_ST.scala 31:71]
  assign _GEN_219 = 8'hdb == WADDR ? 8'hdb : _GEN_218; // @[RAM_ST.scala 31:71]
  assign _GEN_220 = 8'hdc == WADDR ? 8'hdc : _GEN_219; // @[RAM_ST.scala 31:71]
  assign _GEN_221 = 8'hdd == WADDR ? 8'hdd : _GEN_220; // @[RAM_ST.scala 31:71]
  assign _GEN_222 = 8'hde == WADDR ? 8'hde : _GEN_221; // @[RAM_ST.scala 31:71]
  assign _GEN_223 = 8'hdf == WADDR ? 8'hdf : _GEN_222; // @[RAM_ST.scala 31:71]
  assign _GEN_224 = 8'he0 == WADDR ? 8'he0 : _GEN_223; // @[RAM_ST.scala 31:71]
  assign _GEN_225 = 8'he1 == WADDR ? 8'he1 : _GEN_224; // @[RAM_ST.scala 31:71]
  assign _GEN_226 = 8'he2 == WADDR ? 8'he2 : _GEN_225; // @[RAM_ST.scala 31:71]
  assign _GEN_227 = 8'he3 == WADDR ? 8'he3 : _GEN_226; // @[RAM_ST.scala 31:71]
  assign _GEN_228 = 8'he4 == WADDR ? 8'he4 : _GEN_227; // @[RAM_ST.scala 31:71]
  assign _GEN_229 = 8'he5 == WADDR ? 8'he5 : _GEN_228; // @[RAM_ST.scala 31:71]
  assign _GEN_230 = 8'he6 == WADDR ? 8'he6 : _GEN_229; // @[RAM_ST.scala 31:71]
  assign _GEN_231 = 8'he7 == WADDR ? 8'he7 : _GEN_230; // @[RAM_ST.scala 31:71]
  assign _GEN_232 = 8'he8 == WADDR ? 8'he8 : _GEN_231; // @[RAM_ST.scala 31:71]
  assign _GEN_233 = 8'he9 == WADDR ? 8'he9 : _GEN_232; // @[RAM_ST.scala 31:71]
  assign _GEN_234 = 8'hea == WADDR ? 8'hea : _GEN_233; // @[RAM_ST.scala 31:71]
  assign _GEN_235 = 8'heb == WADDR ? 8'heb : _GEN_234; // @[RAM_ST.scala 31:71]
  assign _GEN_236 = 8'hec == WADDR ? 8'hec : _GEN_235; // @[RAM_ST.scala 31:71]
  assign _GEN_237 = 8'hed == WADDR ? 8'hed : _GEN_236; // @[RAM_ST.scala 31:71]
  assign _GEN_238 = 8'hee == WADDR ? 8'hee : _GEN_237; // @[RAM_ST.scala 31:71]
  assign _GEN_239 = 8'hef == WADDR ? 8'hef : _GEN_238; // @[RAM_ST.scala 31:71]
  assign _T = {{1'd0}, _GEN_239}; // @[RAM_ST.scala 31:71]
  assign _GEN_246 = 8'h1 == RADDR ? 8'h1 : 8'h0; // @[RAM_ST.scala 32:46]
  assign _GEN_247 = 8'h2 == RADDR ? 8'h2 : _GEN_246; // @[RAM_ST.scala 32:46]
  assign _GEN_248 = 8'h3 == RADDR ? 8'h3 : _GEN_247; // @[RAM_ST.scala 32:46]
  assign _GEN_249 = 8'h4 == RADDR ? 8'h4 : _GEN_248; // @[RAM_ST.scala 32:46]
  assign _GEN_250 = 8'h5 == RADDR ? 8'h5 : _GEN_249; // @[RAM_ST.scala 32:46]
  assign _GEN_251 = 8'h6 == RADDR ? 8'h6 : _GEN_250; // @[RAM_ST.scala 32:46]
  assign _GEN_252 = 8'h7 == RADDR ? 8'h7 : _GEN_251; // @[RAM_ST.scala 32:46]
  assign _GEN_253 = 8'h8 == RADDR ? 8'h8 : _GEN_252; // @[RAM_ST.scala 32:46]
  assign _GEN_254 = 8'h9 == RADDR ? 8'h9 : _GEN_253; // @[RAM_ST.scala 32:46]
  assign _GEN_255 = 8'ha == RADDR ? 8'ha : _GEN_254; // @[RAM_ST.scala 32:46]
  assign _GEN_256 = 8'hb == RADDR ? 8'hb : _GEN_255; // @[RAM_ST.scala 32:46]
  assign _GEN_257 = 8'hc == RADDR ? 8'hc : _GEN_256; // @[RAM_ST.scala 32:46]
  assign _GEN_258 = 8'hd == RADDR ? 8'hd : _GEN_257; // @[RAM_ST.scala 32:46]
  assign _GEN_259 = 8'he == RADDR ? 8'he : _GEN_258; // @[RAM_ST.scala 32:46]
  assign _GEN_260 = 8'hf == RADDR ? 8'hf : _GEN_259; // @[RAM_ST.scala 32:46]
  assign _GEN_261 = 8'h10 == RADDR ? 8'h10 : _GEN_260; // @[RAM_ST.scala 32:46]
  assign _GEN_262 = 8'h11 == RADDR ? 8'h11 : _GEN_261; // @[RAM_ST.scala 32:46]
  assign _GEN_263 = 8'h12 == RADDR ? 8'h12 : _GEN_262; // @[RAM_ST.scala 32:46]
  assign _GEN_264 = 8'h13 == RADDR ? 8'h13 : _GEN_263; // @[RAM_ST.scala 32:46]
  assign _GEN_265 = 8'h14 == RADDR ? 8'h14 : _GEN_264; // @[RAM_ST.scala 32:46]
  assign _GEN_266 = 8'h15 == RADDR ? 8'h15 : _GEN_265; // @[RAM_ST.scala 32:46]
  assign _GEN_267 = 8'h16 == RADDR ? 8'h16 : _GEN_266; // @[RAM_ST.scala 32:46]
  assign _GEN_268 = 8'h17 == RADDR ? 8'h17 : _GEN_267; // @[RAM_ST.scala 32:46]
  assign _GEN_269 = 8'h18 == RADDR ? 8'h18 : _GEN_268; // @[RAM_ST.scala 32:46]
  assign _GEN_270 = 8'h19 == RADDR ? 8'h19 : _GEN_269; // @[RAM_ST.scala 32:46]
  assign _GEN_271 = 8'h1a == RADDR ? 8'h1a : _GEN_270; // @[RAM_ST.scala 32:46]
  assign _GEN_272 = 8'h1b == RADDR ? 8'h1b : _GEN_271; // @[RAM_ST.scala 32:46]
  assign _GEN_273 = 8'h1c == RADDR ? 8'h1c : _GEN_272; // @[RAM_ST.scala 32:46]
  assign _GEN_274 = 8'h1d == RADDR ? 8'h1d : _GEN_273; // @[RAM_ST.scala 32:46]
  assign _GEN_275 = 8'h1e == RADDR ? 8'h1e : _GEN_274; // @[RAM_ST.scala 32:46]
  assign _GEN_276 = 8'h1f == RADDR ? 8'h1f : _GEN_275; // @[RAM_ST.scala 32:46]
  assign _GEN_277 = 8'h20 == RADDR ? 8'h20 : _GEN_276; // @[RAM_ST.scala 32:46]
  assign _GEN_278 = 8'h21 == RADDR ? 8'h21 : _GEN_277; // @[RAM_ST.scala 32:46]
  assign _GEN_279 = 8'h22 == RADDR ? 8'h22 : _GEN_278; // @[RAM_ST.scala 32:46]
  assign _GEN_280 = 8'h23 == RADDR ? 8'h23 : _GEN_279; // @[RAM_ST.scala 32:46]
  assign _GEN_281 = 8'h24 == RADDR ? 8'h24 : _GEN_280; // @[RAM_ST.scala 32:46]
  assign _GEN_282 = 8'h25 == RADDR ? 8'h25 : _GEN_281; // @[RAM_ST.scala 32:46]
  assign _GEN_283 = 8'h26 == RADDR ? 8'h26 : _GEN_282; // @[RAM_ST.scala 32:46]
  assign _GEN_284 = 8'h27 == RADDR ? 8'h27 : _GEN_283; // @[RAM_ST.scala 32:46]
  assign _GEN_285 = 8'h28 == RADDR ? 8'h28 : _GEN_284; // @[RAM_ST.scala 32:46]
  assign _GEN_286 = 8'h29 == RADDR ? 8'h29 : _GEN_285; // @[RAM_ST.scala 32:46]
  assign _GEN_287 = 8'h2a == RADDR ? 8'h2a : _GEN_286; // @[RAM_ST.scala 32:46]
  assign _GEN_288 = 8'h2b == RADDR ? 8'h2b : _GEN_287; // @[RAM_ST.scala 32:46]
  assign _GEN_289 = 8'h2c == RADDR ? 8'h2c : _GEN_288; // @[RAM_ST.scala 32:46]
  assign _GEN_290 = 8'h2d == RADDR ? 8'h2d : _GEN_289; // @[RAM_ST.scala 32:46]
  assign _GEN_291 = 8'h2e == RADDR ? 8'h2e : _GEN_290; // @[RAM_ST.scala 32:46]
  assign _GEN_292 = 8'h2f == RADDR ? 8'h2f : _GEN_291; // @[RAM_ST.scala 32:46]
  assign _GEN_293 = 8'h30 == RADDR ? 8'h30 : _GEN_292; // @[RAM_ST.scala 32:46]
  assign _GEN_294 = 8'h31 == RADDR ? 8'h31 : _GEN_293; // @[RAM_ST.scala 32:46]
  assign _GEN_295 = 8'h32 == RADDR ? 8'h32 : _GEN_294; // @[RAM_ST.scala 32:46]
  assign _GEN_296 = 8'h33 == RADDR ? 8'h33 : _GEN_295; // @[RAM_ST.scala 32:46]
  assign _GEN_297 = 8'h34 == RADDR ? 8'h34 : _GEN_296; // @[RAM_ST.scala 32:46]
  assign _GEN_298 = 8'h35 == RADDR ? 8'h35 : _GEN_297; // @[RAM_ST.scala 32:46]
  assign _GEN_299 = 8'h36 == RADDR ? 8'h36 : _GEN_298; // @[RAM_ST.scala 32:46]
  assign _GEN_300 = 8'h37 == RADDR ? 8'h37 : _GEN_299; // @[RAM_ST.scala 32:46]
  assign _GEN_301 = 8'h38 == RADDR ? 8'h38 : _GEN_300; // @[RAM_ST.scala 32:46]
  assign _GEN_302 = 8'h39 == RADDR ? 8'h39 : _GEN_301; // @[RAM_ST.scala 32:46]
  assign _GEN_303 = 8'h3a == RADDR ? 8'h3a : _GEN_302; // @[RAM_ST.scala 32:46]
  assign _GEN_304 = 8'h3b == RADDR ? 8'h3b : _GEN_303; // @[RAM_ST.scala 32:46]
  assign _GEN_305 = 8'h3c == RADDR ? 8'h3c : _GEN_304; // @[RAM_ST.scala 32:46]
  assign _GEN_306 = 8'h3d == RADDR ? 8'h3d : _GEN_305; // @[RAM_ST.scala 32:46]
  assign _GEN_307 = 8'h3e == RADDR ? 8'h3e : _GEN_306; // @[RAM_ST.scala 32:46]
  assign _GEN_308 = 8'h3f == RADDR ? 8'h3f : _GEN_307; // @[RAM_ST.scala 32:46]
  assign _GEN_309 = 8'h40 == RADDR ? 8'h40 : _GEN_308; // @[RAM_ST.scala 32:46]
  assign _GEN_310 = 8'h41 == RADDR ? 8'h41 : _GEN_309; // @[RAM_ST.scala 32:46]
  assign _GEN_311 = 8'h42 == RADDR ? 8'h42 : _GEN_310; // @[RAM_ST.scala 32:46]
  assign _GEN_312 = 8'h43 == RADDR ? 8'h43 : _GEN_311; // @[RAM_ST.scala 32:46]
  assign _GEN_313 = 8'h44 == RADDR ? 8'h44 : _GEN_312; // @[RAM_ST.scala 32:46]
  assign _GEN_314 = 8'h45 == RADDR ? 8'h45 : _GEN_313; // @[RAM_ST.scala 32:46]
  assign _GEN_315 = 8'h46 == RADDR ? 8'h46 : _GEN_314; // @[RAM_ST.scala 32:46]
  assign _GEN_316 = 8'h47 == RADDR ? 8'h47 : _GEN_315; // @[RAM_ST.scala 32:46]
  assign _GEN_317 = 8'h48 == RADDR ? 8'h48 : _GEN_316; // @[RAM_ST.scala 32:46]
  assign _GEN_318 = 8'h49 == RADDR ? 8'h49 : _GEN_317; // @[RAM_ST.scala 32:46]
  assign _GEN_319 = 8'h4a == RADDR ? 8'h4a : _GEN_318; // @[RAM_ST.scala 32:46]
  assign _GEN_320 = 8'h4b == RADDR ? 8'h4b : _GEN_319; // @[RAM_ST.scala 32:46]
  assign _GEN_321 = 8'h4c == RADDR ? 8'h4c : _GEN_320; // @[RAM_ST.scala 32:46]
  assign _GEN_322 = 8'h4d == RADDR ? 8'h4d : _GEN_321; // @[RAM_ST.scala 32:46]
  assign _GEN_323 = 8'h4e == RADDR ? 8'h4e : _GEN_322; // @[RAM_ST.scala 32:46]
  assign _GEN_324 = 8'h4f == RADDR ? 8'h4f : _GEN_323; // @[RAM_ST.scala 32:46]
  assign _GEN_325 = 8'h50 == RADDR ? 8'h50 : _GEN_324; // @[RAM_ST.scala 32:46]
  assign _GEN_326 = 8'h51 == RADDR ? 8'h51 : _GEN_325; // @[RAM_ST.scala 32:46]
  assign _GEN_327 = 8'h52 == RADDR ? 8'h52 : _GEN_326; // @[RAM_ST.scala 32:46]
  assign _GEN_328 = 8'h53 == RADDR ? 8'h53 : _GEN_327; // @[RAM_ST.scala 32:46]
  assign _GEN_329 = 8'h54 == RADDR ? 8'h54 : _GEN_328; // @[RAM_ST.scala 32:46]
  assign _GEN_330 = 8'h55 == RADDR ? 8'h55 : _GEN_329; // @[RAM_ST.scala 32:46]
  assign _GEN_331 = 8'h56 == RADDR ? 8'h56 : _GEN_330; // @[RAM_ST.scala 32:46]
  assign _GEN_332 = 8'h57 == RADDR ? 8'h57 : _GEN_331; // @[RAM_ST.scala 32:46]
  assign _GEN_333 = 8'h58 == RADDR ? 8'h58 : _GEN_332; // @[RAM_ST.scala 32:46]
  assign _GEN_334 = 8'h59 == RADDR ? 8'h59 : _GEN_333; // @[RAM_ST.scala 32:46]
  assign _GEN_335 = 8'h5a == RADDR ? 8'h5a : _GEN_334; // @[RAM_ST.scala 32:46]
  assign _GEN_336 = 8'h5b == RADDR ? 8'h5b : _GEN_335; // @[RAM_ST.scala 32:46]
  assign _GEN_337 = 8'h5c == RADDR ? 8'h5c : _GEN_336; // @[RAM_ST.scala 32:46]
  assign _GEN_338 = 8'h5d == RADDR ? 8'h5d : _GEN_337; // @[RAM_ST.scala 32:46]
  assign _GEN_339 = 8'h5e == RADDR ? 8'h5e : _GEN_338; // @[RAM_ST.scala 32:46]
  assign _GEN_340 = 8'h5f == RADDR ? 8'h5f : _GEN_339; // @[RAM_ST.scala 32:46]
  assign _GEN_341 = 8'h60 == RADDR ? 8'h60 : _GEN_340; // @[RAM_ST.scala 32:46]
  assign _GEN_342 = 8'h61 == RADDR ? 8'h61 : _GEN_341; // @[RAM_ST.scala 32:46]
  assign _GEN_343 = 8'h62 == RADDR ? 8'h62 : _GEN_342; // @[RAM_ST.scala 32:46]
  assign _GEN_344 = 8'h63 == RADDR ? 8'h63 : _GEN_343; // @[RAM_ST.scala 32:46]
  assign _GEN_345 = 8'h64 == RADDR ? 8'h64 : _GEN_344; // @[RAM_ST.scala 32:46]
  assign _GEN_346 = 8'h65 == RADDR ? 8'h65 : _GEN_345; // @[RAM_ST.scala 32:46]
  assign _GEN_347 = 8'h66 == RADDR ? 8'h66 : _GEN_346; // @[RAM_ST.scala 32:46]
  assign _GEN_348 = 8'h67 == RADDR ? 8'h67 : _GEN_347; // @[RAM_ST.scala 32:46]
  assign _GEN_349 = 8'h68 == RADDR ? 8'h68 : _GEN_348; // @[RAM_ST.scala 32:46]
  assign _GEN_350 = 8'h69 == RADDR ? 8'h69 : _GEN_349; // @[RAM_ST.scala 32:46]
  assign _GEN_351 = 8'h6a == RADDR ? 8'h6a : _GEN_350; // @[RAM_ST.scala 32:46]
  assign _GEN_352 = 8'h6b == RADDR ? 8'h6b : _GEN_351; // @[RAM_ST.scala 32:46]
  assign _GEN_353 = 8'h6c == RADDR ? 8'h6c : _GEN_352; // @[RAM_ST.scala 32:46]
  assign _GEN_354 = 8'h6d == RADDR ? 8'h6d : _GEN_353; // @[RAM_ST.scala 32:46]
  assign _GEN_355 = 8'h6e == RADDR ? 8'h6e : _GEN_354; // @[RAM_ST.scala 32:46]
  assign _GEN_356 = 8'h6f == RADDR ? 8'h6f : _GEN_355; // @[RAM_ST.scala 32:46]
  assign _GEN_357 = 8'h70 == RADDR ? 8'h70 : _GEN_356; // @[RAM_ST.scala 32:46]
  assign _GEN_358 = 8'h71 == RADDR ? 8'h71 : _GEN_357; // @[RAM_ST.scala 32:46]
  assign _GEN_359 = 8'h72 == RADDR ? 8'h72 : _GEN_358; // @[RAM_ST.scala 32:46]
  assign _GEN_360 = 8'h73 == RADDR ? 8'h73 : _GEN_359; // @[RAM_ST.scala 32:46]
  assign _GEN_361 = 8'h74 == RADDR ? 8'h74 : _GEN_360; // @[RAM_ST.scala 32:46]
  assign _GEN_362 = 8'h75 == RADDR ? 8'h75 : _GEN_361; // @[RAM_ST.scala 32:46]
  assign _GEN_363 = 8'h76 == RADDR ? 8'h76 : _GEN_362; // @[RAM_ST.scala 32:46]
  assign _GEN_364 = 8'h77 == RADDR ? 8'h77 : _GEN_363; // @[RAM_ST.scala 32:46]
  assign _GEN_365 = 8'h78 == RADDR ? 8'h78 : _GEN_364; // @[RAM_ST.scala 32:46]
  assign _GEN_366 = 8'h79 == RADDR ? 8'h79 : _GEN_365; // @[RAM_ST.scala 32:46]
  assign _GEN_367 = 8'h7a == RADDR ? 8'h7a : _GEN_366; // @[RAM_ST.scala 32:46]
  assign _GEN_368 = 8'h7b == RADDR ? 8'h7b : _GEN_367; // @[RAM_ST.scala 32:46]
  assign _GEN_369 = 8'h7c == RADDR ? 8'h7c : _GEN_368; // @[RAM_ST.scala 32:46]
  assign _GEN_370 = 8'h7d == RADDR ? 8'h7d : _GEN_369; // @[RAM_ST.scala 32:46]
  assign _GEN_371 = 8'h7e == RADDR ? 8'h7e : _GEN_370; // @[RAM_ST.scala 32:46]
  assign _GEN_372 = 8'h7f == RADDR ? 8'h7f : _GEN_371; // @[RAM_ST.scala 32:46]
  assign _GEN_373 = 8'h80 == RADDR ? 8'h80 : _GEN_372; // @[RAM_ST.scala 32:46]
  assign _GEN_374 = 8'h81 == RADDR ? 8'h81 : _GEN_373; // @[RAM_ST.scala 32:46]
  assign _GEN_375 = 8'h82 == RADDR ? 8'h82 : _GEN_374; // @[RAM_ST.scala 32:46]
  assign _GEN_376 = 8'h83 == RADDR ? 8'h83 : _GEN_375; // @[RAM_ST.scala 32:46]
  assign _GEN_377 = 8'h84 == RADDR ? 8'h84 : _GEN_376; // @[RAM_ST.scala 32:46]
  assign _GEN_378 = 8'h85 == RADDR ? 8'h85 : _GEN_377; // @[RAM_ST.scala 32:46]
  assign _GEN_379 = 8'h86 == RADDR ? 8'h86 : _GEN_378; // @[RAM_ST.scala 32:46]
  assign _GEN_380 = 8'h87 == RADDR ? 8'h87 : _GEN_379; // @[RAM_ST.scala 32:46]
  assign _GEN_381 = 8'h88 == RADDR ? 8'h88 : _GEN_380; // @[RAM_ST.scala 32:46]
  assign _GEN_382 = 8'h89 == RADDR ? 8'h89 : _GEN_381; // @[RAM_ST.scala 32:46]
  assign _GEN_383 = 8'h8a == RADDR ? 8'h8a : _GEN_382; // @[RAM_ST.scala 32:46]
  assign _GEN_384 = 8'h8b == RADDR ? 8'h8b : _GEN_383; // @[RAM_ST.scala 32:46]
  assign _GEN_385 = 8'h8c == RADDR ? 8'h8c : _GEN_384; // @[RAM_ST.scala 32:46]
  assign _GEN_386 = 8'h8d == RADDR ? 8'h8d : _GEN_385; // @[RAM_ST.scala 32:46]
  assign _GEN_387 = 8'h8e == RADDR ? 8'h8e : _GEN_386; // @[RAM_ST.scala 32:46]
  assign _GEN_388 = 8'h8f == RADDR ? 8'h8f : _GEN_387; // @[RAM_ST.scala 32:46]
  assign _GEN_389 = 8'h90 == RADDR ? 8'h90 : _GEN_388; // @[RAM_ST.scala 32:46]
  assign _GEN_390 = 8'h91 == RADDR ? 8'h91 : _GEN_389; // @[RAM_ST.scala 32:46]
  assign _GEN_391 = 8'h92 == RADDR ? 8'h92 : _GEN_390; // @[RAM_ST.scala 32:46]
  assign _GEN_392 = 8'h93 == RADDR ? 8'h93 : _GEN_391; // @[RAM_ST.scala 32:46]
  assign _GEN_393 = 8'h94 == RADDR ? 8'h94 : _GEN_392; // @[RAM_ST.scala 32:46]
  assign _GEN_394 = 8'h95 == RADDR ? 8'h95 : _GEN_393; // @[RAM_ST.scala 32:46]
  assign _GEN_395 = 8'h96 == RADDR ? 8'h96 : _GEN_394; // @[RAM_ST.scala 32:46]
  assign _GEN_396 = 8'h97 == RADDR ? 8'h97 : _GEN_395; // @[RAM_ST.scala 32:46]
  assign _GEN_397 = 8'h98 == RADDR ? 8'h98 : _GEN_396; // @[RAM_ST.scala 32:46]
  assign _GEN_398 = 8'h99 == RADDR ? 8'h99 : _GEN_397; // @[RAM_ST.scala 32:46]
  assign _GEN_399 = 8'h9a == RADDR ? 8'h9a : _GEN_398; // @[RAM_ST.scala 32:46]
  assign _GEN_400 = 8'h9b == RADDR ? 8'h9b : _GEN_399; // @[RAM_ST.scala 32:46]
  assign _GEN_401 = 8'h9c == RADDR ? 8'h9c : _GEN_400; // @[RAM_ST.scala 32:46]
  assign _GEN_402 = 8'h9d == RADDR ? 8'h9d : _GEN_401; // @[RAM_ST.scala 32:46]
  assign _GEN_403 = 8'h9e == RADDR ? 8'h9e : _GEN_402; // @[RAM_ST.scala 32:46]
  assign _GEN_404 = 8'h9f == RADDR ? 8'h9f : _GEN_403; // @[RAM_ST.scala 32:46]
  assign _GEN_405 = 8'ha0 == RADDR ? 8'ha0 : _GEN_404; // @[RAM_ST.scala 32:46]
  assign _GEN_406 = 8'ha1 == RADDR ? 8'ha1 : _GEN_405; // @[RAM_ST.scala 32:46]
  assign _GEN_407 = 8'ha2 == RADDR ? 8'ha2 : _GEN_406; // @[RAM_ST.scala 32:46]
  assign _GEN_408 = 8'ha3 == RADDR ? 8'ha3 : _GEN_407; // @[RAM_ST.scala 32:46]
  assign _GEN_409 = 8'ha4 == RADDR ? 8'ha4 : _GEN_408; // @[RAM_ST.scala 32:46]
  assign _GEN_410 = 8'ha5 == RADDR ? 8'ha5 : _GEN_409; // @[RAM_ST.scala 32:46]
  assign _GEN_411 = 8'ha6 == RADDR ? 8'ha6 : _GEN_410; // @[RAM_ST.scala 32:46]
  assign _GEN_412 = 8'ha7 == RADDR ? 8'ha7 : _GEN_411; // @[RAM_ST.scala 32:46]
  assign _GEN_413 = 8'ha8 == RADDR ? 8'ha8 : _GEN_412; // @[RAM_ST.scala 32:46]
  assign _GEN_414 = 8'ha9 == RADDR ? 8'ha9 : _GEN_413; // @[RAM_ST.scala 32:46]
  assign _GEN_415 = 8'haa == RADDR ? 8'haa : _GEN_414; // @[RAM_ST.scala 32:46]
  assign _GEN_416 = 8'hab == RADDR ? 8'hab : _GEN_415; // @[RAM_ST.scala 32:46]
  assign _GEN_417 = 8'hac == RADDR ? 8'hac : _GEN_416; // @[RAM_ST.scala 32:46]
  assign _GEN_418 = 8'had == RADDR ? 8'had : _GEN_417; // @[RAM_ST.scala 32:46]
  assign _GEN_419 = 8'hae == RADDR ? 8'hae : _GEN_418; // @[RAM_ST.scala 32:46]
  assign _GEN_420 = 8'haf == RADDR ? 8'haf : _GEN_419; // @[RAM_ST.scala 32:46]
  assign _GEN_421 = 8'hb0 == RADDR ? 8'hb0 : _GEN_420; // @[RAM_ST.scala 32:46]
  assign _GEN_422 = 8'hb1 == RADDR ? 8'hb1 : _GEN_421; // @[RAM_ST.scala 32:46]
  assign _GEN_423 = 8'hb2 == RADDR ? 8'hb2 : _GEN_422; // @[RAM_ST.scala 32:46]
  assign _GEN_424 = 8'hb3 == RADDR ? 8'hb3 : _GEN_423; // @[RAM_ST.scala 32:46]
  assign _GEN_425 = 8'hb4 == RADDR ? 8'hb4 : _GEN_424; // @[RAM_ST.scala 32:46]
  assign _GEN_426 = 8'hb5 == RADDR ? 8'hb5 : _GEN_425; // @[RAM_ST.scala 32:46]
  assign _GEN_427 = 8'hb6 == RADDR ? 8'hb6 : _GEN_426; // @[RAM_ST.scala 32:46]
  assign _GEN_428 = 8'hb7 == RADDR ? 8'hb7 : _GEN_427; // @[RAM_ST.scala 32:46]
  assign _GEN_429 = 8'hb8 == RADDR ? 8'hb8 : _GEN_428; // @[RAM_ST.scala 32:46]
  assign _GEN_430 = 8'hb9 == RADDR ? 8'hb9 : _GEN_429; // @[RAM_ST.scala 32:46]
  assign _GEN_431 = 8'hba == RADDR ? 8'hba : _GEN_430; // @[RAM_ST.scala 32:46]
  assign _GEN_432 = 8'hbb == RADDR ? 8'hbb : _GEN_431; // @[RAM_ST.scala 32:46]
  assign _GEN_433 = 8'hbc == RADDR ? 8'hbc : _GEN_432; // @[RAM_ST.scala 32:46]
  assign _GEN_434 = 8'hbd == RADDR ? 8'hbd : _GEN_433; // @[RAM_ST.scala 32:46]
  assign _GEN_435 = 8'hbe == RADDR ? 8'hbe : _GEN_434; // @[RAM_ST.scala 32:46]
  assign _GEN_436 = 8'hbf == RADDR ? 8'hbf : _GEN_435; // @[RAM_ST.scala 32:46]
  assign _GEN_437 = 8'hc0 == RADDR ? 8'hc0 : _GEN_436; // @[RAM_ST.scala 32:46]
  assign _GEN_438 = 8'hc1 == RADDR ? 8'hc1 : _GEN_437; // @[RAM_ST.scala 32:46]
  assign _GEN_439 = 8'hc2 == RADDR ? 8'hc2 : _GEN_438; // @[RAM_ST.scala 32:46]
  assign _GEN_440 = 8'hc3 == RADDR ? 8'hc3 : _GEN_439; // @[RAM_ST.scala 32:46]
  assign _GEN_441 = 8'hc4 == RADDR ? 8'hc4 : _GEN_440; // @[RAM_ST.scala 32:46]
  assign _GEN_442 = 8'hc5 == RADDR ? 8'hc5 : _GEN_441; // @[RAM_ST.scala 32:46]
  assign _GEN_443 = 8'hc6 == RADDR ? 8'hc6 : _GEN_442; // @[RAM_ST.scala 32:46]
  assign _GEN_444 = 8'hc7 == RADDR ? 8'hc7 : _GEN_443; // @[RAM_ST.scala 32:46]
  assign _GEN_445 = 8'hc8 == RADDR ? 8'hc8 : _GEN_444; // @[RAM_ST.scala 32:46]
  assign _GEN_446 = 8'hc9 == RADDR ? 8'hc9 : _GEN_445; // @[RAM_ST.scala 32:46]
  assign _GEN_447 = 8'hca == RADDR ? 8'hca : _GEN_446; // @[RAM_ST.scala 32:46]
  assign _GEN_448 = 8'hcb == RADDR ? 8'hcb : _GEN_447; // @[RAM_ST.scala 32:46]
  assign _GEN_449 = 8'hcc == RADDR ? 8'hcc : _GEN_448; // @[RAM_ST.scala 32:46]
  assign _GEN_450 = 8'hcd == RADDR ? 8'hcd : _GEN_449; // @[RAM_ST.scala 32:46]
  assign _GEN_451 = 8'hce == RADDR ? 8'hce : _GEN_450; // @[RAM_ST.scala 32:46]
  assign _GEN_452 = 8'hcf == RADDR ? 8'hcf : _GEN_451; // @[RAM_ST.scala 32:46]
  assign _GEN_453 = 8'hd0 == RADDR ? 8'hd0 : _GEN_452; // @[RAM_ST.scala 32:46]
  assign _GEN_454 = 8'hd1 == RADDR ? 8'hd1 : _GEN_453; // @[RAM_ST.scala 32:46]
  assign _GEN_455 = 8'hd2 == RADDR ? 8'hd2 : _GEN_454; // @[RAM_ST.scala 32:46]
  assign _GEN_456 = 8'hd3 == RADDR ? 8'hd3 : _GEN_455; // @[RAM_ST.scala 32:46]
  assign _GEN_457 = 8'hd4 == RADDR ? 8'hd4 : _GEN_456; // @[RAM_ST.scala 32:46]
  assign _GEN_458 = 8'hd5 == RADDR ? 8'hd5 : _GEN_457; // @[RAM_ST.scala 32:46]
  assign _GEN_459 = 8'hd6 == RADDR ? 8'hd6 : _GEN_458; // @[RAM_ST.scala 32:46]
  assign _GEN_460 = 8'hd7 == RADDR ? 8'hd7 : _GEN_459; // @[RAM_ST.scala 32:46]
  assign _GEN_461 = 8'hd8 == RADDR ? 8'hd8 : _GEN_460; // @[RAM_ST.scala 32:46]
  assign _GEN_462 = 8'hd9 == RADDR ? 8'hd9 : _GEN_461; // @[RAM_ST.scala 32:46]
  assign _GEN_463 = 8'hda == RADDR ? 8'hda : _GEN_462; // @[RAM_ST.scala 32:46]
  assign _GEN_464 = 8'hdb == RADDR ? 8'hdb : _GEN_463; // @[RAM_ST.scala 32:46]
  assign _GEN_465 = 8'hdc == RADDR ? 8'hdc : _GEN_464; // @[RAM_ST.scala 32:46]
  assign _GEN_466 = 8'hdd == RADDR ? 8'hdd : _GEN_465; // @[RAM_ST.scala 32:46]
  assign _GEN_467 = 8'hde == RADDR ? 8'hde : _GEN_466; // @[RAM_ST.scala 32:46]
  assign _GEN_468 = 8'hdf == RADDR ? 8'hdf : _GEN_467; // @[RAM_ST.scala 32:46]
  assign _GEN_469 = 8'he0 == RADDR ? 8'he0 : _GEN_468; // @[RAM_ST.scala 32:46]
  assign _GEN_470 = 8'he1 == RADDR ? 8'he1 : _GEN_469; // @[RAM_ST.scala 32:46]
  assign _GEN_471 = 8'he2 == RADDR ? 8'he2 : _GEN_470; // @[RAM_ST.scala 32:46]
  assign _GEN_472 = 8'he3 == RADDR ? 8'he3 : _GEN_471; // @[RAM_ST.scala 32:46]
  assign _GEN_473 = 8'he4 == RADDR ? 8'he4 : _GEN_472; // @[RAM_ST.scala 32:46]
  assign _GEN_474 = 8'he5 == RADDR ? 8'he5 : _GEN_473; // @[RAM_ST.scala 32:46]
  assign _GEN_475 = 8'he6 == RADDR ? 8'he6 : _GEN_474; // @[RAM_ST.scala 32:46]
  assign _GEN_476 = 8'he7 == RADDR ? 8'he7 : _GEN_475; // @[RAM_ST.scala 32:46]
  assign _GEN_477 = 8'he8 == RADDR ? 8'he8 : _GEN_476; // @[RAM_ST.scala 32:46]
  assign _GEN_478 = 8'he9 == RADDR ? 8'he9 : _GEN_477; // @[RAM_ST.scala 32:46]
  assign _GEN_479 = 8'hea == RADDR ? 8'hea : _GEN_478; // @[RAM_ST.scala 32:46]
  assign _GEN_480 = 8'heb == RADDR ? 8'heb : _GEN_479; // @[RAM_ST.scala 32:46]
  assign _GEN_481 = 8'hec == RADDR ? 8'hec : _GEN_480; // @[RAM_ST.scala 32:46]
  assign _GEN_482 = 8'hed == RADDR ? 8'hed : _GEN_481; // @[RAM_ST.scala 32:46]
  assign _GEN_483 = 8'hee == RADDR ? 8'hee : _GEN_482; // @[RAM_ST.scala 32:46]
  assign _GEN_484 = 8'hef == RADDR ? 8'hef : _GEN_483; // @[RAM_ST.scala 32:46]
  assign _T_3 = {{1'd0}, _GEN_484}; // @[RAM_ST.scala 32:46]
  assign RDATA_0_0 = ram_0_0__T_8_data; // @[RAM_ST.scala 32:9]
  assign write_elem_counter_CE = WE; // @[RAM_ST.scala 23:25]
  assign read_elem_counter_CE = RE; // @[RAM_ST.scala 24:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 240; initvar = initvar+1)
    ram_0_0[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_0_0__T_8_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ram_0_0__T_8_addr_pipe_0 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_0_0__T_2_en & ram_0_0__T_2_mask) begin
      ram_0_0[ram_0_0__T_2_addr] <= ram_0_0__T_2_data; // @[RAM_ST.scala 29:24]
    end
    ram_0_0__T_8_en_pipe_0 <= read_elem_counter_valid;
    if (read_elem_counter_valid) begin
      ram_0_0__T_8_addr_pipe_0 <= _T_3[7:0];
    end
  end
endmodule
module ShiftT(
  input        clock,
  input        reset,
  input        valid_up,
  input  [7:0] I_0_0,
  output [7:0] O_0_0
);
  wire  RAM_ST_clock; // @[ShiftT.scala 39:29]
  wire  RAM_ST_RE; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_RADDR; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_RDATA_0_0; // @[ShiftT.scala 39:29]
  wire  RAM_ST_WE; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_WADDR; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_WDATA_0_0; // @[ShiftT.scala 39:29]
  wire  NestedCounters_CE; // @[ShiftT.scala 41:31]
  wire  NestedCounters_valid; // @[ShiftT.scala 41:31]
  reg [7:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[Counter.scala 37:24]
  wire [7:0] _T_3; // @[Counter.scala 38:22]
  RAM_ST RAM_ST ( // @[ShiftT.scala 39:29]
    .clock(RAM_ST_clock),
    .RE(RAM_ST_RE),
    .RADDR(RAM_ST_RADDR),
    .RDATA_0_0(RAM_ST_RDATA_0_0),
    .WE(RAM_ST_WE),
    .WADDR(RAM_ST_WADDR),
    .WDATA_0_0(RAM_ST_WDATA_0_0)
  );
  NestedCounters_2 NestedCounters ( // @[ShiftT.scala 41:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign _T_1 = value == 8'hef; // @[Counter.scala 37:24]
  assign _T_3 = value + 8'h1; // @[Counter.scala 38:22]
  assign O_0_0 = RAM_ST_RDATA_0_0; // @[ShiftT.scala 51:7]
  assign RAM_ST_clock = clock;
  assign RAM_ST_RE = valid_up; // @[ShiftT.scala 49:20]
  assign RAM_ST_RADDR = _T_1 ? 8'h0 : _T_3; // @[ShiftT.scala 46:76 ShiftT.scala 47:38]
  assign RAM_ST_WE = valid_up; // @[ShiftT.scala 48:20]
  assign RAM_ST_WADDR = value; // @[ShiftT.scala 45:23]
  assign RAM_ST_WDATA_0_0 = I_0_0; // @[ShiftT.scala 50:23]
  assign NestedCounters_CE = valid_up; // @[ShiftT.scala 42:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 8'h0;
    end else if (valid_up) begin
      if (_T_1) begin
        value <= 8'h0;
      end else begin
        value <= _T_3;
      end
    end
  end
endmodule
module ShiftTS(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_1_0_0,
  input  [7:0] I_2_0_0,
  input  [7:0] I_3_0_0,
  input  [7:0] I_4_0_0,
  input  [7:0] I_5_0_0,
  input  [7:0] I_6_0_0,
  input  [7:0] I_7_0_0,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_1_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_1_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_1_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_1_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_1_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_2_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_2_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_2_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_2_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_2_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_3_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_3_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_3_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_3_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_3_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_4_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_4_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_4_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_4_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_4_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_5_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_5_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_5_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_5_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_5_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_6_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_6_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_6_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_6_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_6_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_7_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_7_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_7_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_7_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_7_O_0_0; // @[ShiftTS.scala 32:34]
  ShiftT ShiftT ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_clock),
    .reset(ShiftT_reset),
    .valid_up(ShiftT_valid_up),
    .I_0_0(ShiftT_I_0_0),
    .O_0_0(ShiftT_O_0_0)
  );
  ShiftT ShiftT_1 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_1_clock),
    .reset(ShiftT_1_reset),
    .valid_up(ShiftT_1_valid_up),
    .I_0_0(ShiftT_1_I_0_0),
    .O_0_0(ShiftT_1_O_0_0)
  );
  ShiftT ShiftT_2 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_2_clock),
    .reset(ShiftT_2_reset),
    .valid_up(ShiftT_2_valid_up),
    .I_0_0(ShiftT_2_I_0_0),
    .O_0_0(ShiftT_2_O_0_0)
  );
  ShiftT ShiftT_3 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_3_clock),
    .reset(ShiftT_3_reset),
    .valid_up(ShiftT_3_valid_up),
    .I_0_0(ShiftT_3_I_0_0),
    .O_0_0(ShiftT_3_O_0_0)
  );
  ShiftT ShiftT_4 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_4_clock),
    .reset(ShiftT_4_reset),
    .valid_up(ShiftT_4_valid_up),
    .I_0_0(ShiftT_4_I_0_0),
    .O_0_0(ShiftT_4_O_0_0)
  );
  ShiftT ShiftT_5 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_5_clock),
    .reset(ShiftT_5_reset),
    .valid_up(ShiftT_5_valid_up),
    .I_0_0(ShiftT_5_I_0_0),
    .O_0_0(ShiftT_5_O_0_0)
  );
  ShiftT ShiftT_6 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_6_clock),
    .reset(ShiftT_6_reset),
    .valid_up(ShiftT_6_valid_up),
    .I_0_0(ShiftT_6_I_0_0),
    .O_0_0(ShiftT_6_O_0_0)
  );
  ShiftT ShiftT_7 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_7_clock),
    .reset(ShiftT_7_reset),
    .valid_up(ShiftT_7_valid_up),
    .I_0_0(ShiftT_7_I_0_0),
    .O_0_0(ShiftT_7_O_0_0)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 39:14]
  assign O_0_0_0 = ShiftT_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_1_0_0 = ShiftT_1_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_2_0_0 = ShiftT_2_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_3_0_0 = ShiftT_3_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_4_0_0 = ShiftT_4_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_5_0_0 = ShiftT_5_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_6_0_0 = ShiftT_6_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_7_0_0 = ShiftT_7_O_0_0; // @[ShiftTS.scala 34:36]
  assign ShiftT_clock = clock;
  assign ShiftT_reset = reset;
  assign ShiftT_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_I_0_0 = I_0_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_1_clock = clock;
  assign ShiftT_1_reset = reset;
  assign ShiftT_1_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_1_I_0_0 = I_1_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_2_clock = clock;
  assign ShiftT_2_reset = reset;
  assign ShiftT_2_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_2_I_0_0 = I_2_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_3_clock = clock;
  assign ShiftT_3_reset = reset;
  assign ShiftT_3_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_3_I_0_0 = I_3_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_4_clock = clock;
  assign ShiftT_4_reset = reset;
  assign ShiftT_4_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_4_I_0_0 = I_4_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_5_clock = clock;
  assign ShiftT_5_reset = reset;
  assign ShiftT_5_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_5_I_0_0 = I_5_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_6_clock = clock;
  assign ShiftT_6_reset = reset;
  assign ShiftT_6_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_6_I_0_0 = I_6_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_7_clock = clock;
  assign ShiftT_7_reset = reset;
  assign ShiftT_7_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_7_I_0_0 = I_7_0_0; // @[ShiftTS.scala 33:24]
endmodule
module ShiftT_16(
  input        clock,
  input  [7:0] I_0_0,
  output [7:0] O_0_0
);
  reg [7:0] _T_0_0; // @[ShiftT.scala 24:82]
  reg [31:0] _RAND_0;
  assign O_0_0 = _T_0_0; // @[ShiftT.scala 24:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0_0 <= I_0_0;
  end
endmodule
module ShiftTS_2(
  input        clock,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_1_0_0,
  input  [7:0] I_2_0_0,
  input  [7:0] I_3_0_0,
  input  [7:0] I_4_0_0,
  input  [7:0] I_5_0_0,
  input  [7:0] I_6_0_0,
  input  [7:0] I_7_0_0,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_O_0_0; // @[ShiftTS.scala 32:34]
  ShiftT_16 ShiftT ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_clock),
    .I_0_0(ShiftT_I_0_0),
    .O_0_0(ShiftT_O_0_0)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 39:14]
  assign O_0_0_0 = ShiftT_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_1_0_0 = I_0_0_0; // @[ShiftTS.scala 29:36]
  assign O_2_0_0 = I_1_0_0; // @[ShiftTS.scala 29:36]
  assign O_3_0_0 = I_2_0_0; // @[ShiftTS.scala 29:36]
  assign O_4_0_0 = I_3_0_0; // @[ShiftTS.scala 29:36]
  assign O_5_0_0 = I_4_0_0; // @[ShiftTS.scala 29:36]
  assign O_6_0_0 = I_5_0_0; // @[ShiftTS.scala 29:36]
  assign O_7_0_0 = I_6_0_0; // @[ShiftTS.scala 29:36]
  assign ShiftT_clock = clock;
  assign ShiftT_I_0_0 = I_7_0_0; // @[ShiftTS.scala 33:24]
endmodule
module SSeqTupleCreator(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0 = I0; // @[Tuple.scala 12:32]
  assign O_1 = I1; // @[Tuple.scala 13:32]
endmodule
module Map2S(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I1_0,
  output [7:0] O_0_0,
  output [7:0] O_0_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1; // @[Map2S.scala 9:22]
  SSeqTupleCreator fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I1_0_0,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  Map2S fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I1_0(fst_op_I1_0),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_2(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_1_0_0,
  input  [7:0] I0_2_0_0,
  input  [7:0] I0_3_0_0,
  input  [7:0] I0_4_0_0,
  input  [7:0] I0_5_0_0,
  input  [7:0] I0_6_0_0,
  input  [7:0] I0_7_0_0,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_7_0_0,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_1; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_1; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  Map2S_1 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I1_0_0(fst_op_I1_0_0),
    .O_0_0_0(fst_op_O_0_0_0),
    .O_0_0_1(fst_op_O_0_0_1)
  );
  Map2S_1 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0(other_ops_0_I0_0_0),
    .I1_0_0(other_ops_0_I1_0_0),
    .O_0_0_0(other_ops_0_O_0_0_0),
    .O_0_0_1(other_ops_0_O_0_0_1)
  );
  Map2S_1 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0(other_ops_1_I0_0_0),
    .I1_0_0(other_ops_1_I1_0_0),
    .O_0_0_0(other_ops_1_O_0_0_0),
    .O_0_0_1(other_ops_1_O_0_0_1)
  );
  Map2S_1 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0(other_ops_2_I0_0_0),
    .I1_0_0(other_ops_2_I1_0_0),
    .O_0_0_0(other_ops_2_O_0_0_0),
    .O_0_0_1(other_ops_2_O_0_0_1)
  );
  Map2S_1 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0(other_ops_3_I0_0_0),
    .I1_0_0(other_ops_3_I1_0_0),
    .O_0_0_0(other_ops_3_O_0_0_0),
    .O_0_0_1(other_ops_3_O_0_0_1)
  );
  Map2S_1 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0(other_ops_4_I0_0_0),
    .I1_0_0(other_ops_4_I1_0_0),
    .O_0_0_0(other_ops_4_O_0_0_0),
    .O_0_0_1(other_ops_4_O_0_0_1)
  );
  Map2S_1 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0(other_ops_5_I0_0_0),
    .I1_0_0(other_ops_5_I1_0_0),
    .O_0_0_0(other_ops_5_O_0_0_0),
    .O_0_0_1(other_ops_5_O_0_0_1)
  );
  Map2S_1 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0(other_ops_6_I0_0_0),
    .I1_0_0(other_ops_6_I1_0_0),
    .O_0_0_0(other_ops_6_O_0_0_0),
    .O_0_0_1(other_ops_6_O_0_0_1)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0_0 = fst_op_O_0_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_0_1 = fst_op_O_0_0_1; // @[Map2S.scala 19:8]
  assign O_1_0_0_0 = other_ops_0_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_0_1 = other_ops_0_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_0_0 = other_ops_1_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_0_1 = other_ops_1_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_0_0 = other_ops_2_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_0_1 = other_ops_2_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_0_0 = other_ops_3_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_0_1 = other_ops_3_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_0_0 = other_ops_4_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_0_1 = other_ops_4_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_0_0 = other_ops_5_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_0_1 = other_ops_5_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_0_0 = other_ops_6_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_0_1 = other_ops_6_O_0_0_1; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_0 = I1_0_0_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0 = I0_1_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0_0 = I1_1_0_0; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0 = I0_2_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0_0 = I1_2_0_0; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0 = I0_3_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0_0 = I1_3_0_0; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0 = I0_4_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0_0 = I1_4_0_0; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0 = I0_5_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0_0 = I1_5_0_0; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0 = I0_6_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0_0 = I1_6_0_0; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0 = I0_7_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0_0 = I1_7_0_0; // @[Map2S.scala 23:43]
endmodule
module Map2T(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_1_0_0,
  input  [7:0] I0_2_0_0,
  input  [7:0] I0_3_0_0,
  input  [7:0] I0_4_0_0,
  input  [7:0] I0_5_0_0,
  input  [7:0] I0_6_0_0,
  input  [7:0] I0_7_0_0,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_7_0_0,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_1; // @[Map2T.scala 8:20]
  Map2S_2 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0(op_I0_0_0_0),
    .I0_1_0_0(op_I0_1_0_0),
    .I0_2_0_0(op_I0_2_0_0),
    .I0_3_0_0(op_I0_3_0_0),
    .I0_4_0_0(op_I0_4_0_0),
    .I0_5_0_0(op_I0_5_0_0),
    .I0_6_0_0(op_I0_6_0_0),
    .I0_7_0_0(op_I0_7_0_0),
    .I1_0_0_0(op_I1_0_0_0),
    .I1_1_0_0(op_I1_1_0_0),
    .I1_2_0_0(op_I1_2_0_0),
    .I1_3_0_0(op_I1_3_0_0),
    .I1_4_0_0(op_I1_4_0_0),
    .I1_5_0_0(op_I1_5_0_0),
    .I1_6_0_0(op_I1_6_0_0),
    .I1_7_0_0(op_I1_7_0_0),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_4_0_0_0(op_O_4_0_0_0),
    .O_4_0_0_1(op_O_4_0_0_1),
    .O_5_0_0_0(op_O_5_0_0_0),
    .O_5_0_0_1(op_O_5_0_0_1),
    .O_6_0_0_0(op_O_6_0_0_0),
    .O_6_0_0_1(op_O_6_0_0_1),
    .O_7_0_0_0(op_O_7_0_0_0),
    .O_7_0_0_1(op_O_7_0_0_1)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_0_0 = op_O_4_0_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_0_1 = op_O_4_0_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_0_0 = op_O_5_0_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_0_1 = op_O_5_0_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_0_0 = op_O_6_0_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_0_1 = op_O_6_0_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_0_0 = op_O_7_0_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_0_1 = op_O_7_0_0_1; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0 = I0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0 = I0_1_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0 = I0_2_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0 = I0_3_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0 = I0_4_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0 = I0_5_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0 = I0_6_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0 = I0_7_0_0; // @[Map2T.scala 15:11]
  assign op_I1_0_0_0 = I1_0_0_0; // @[Map2T.scala 16:11]
  assign op_I1_1_0_0 = I1_1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_2_0_0 = I1_2_0_0; // @[Map2T.scala 16:11]
  assign op_I1_3_0_0 = I1_3_0_0; // @[Map2T.scala 16:11]
  assign op_I1_4_0_0 = I1_4_0_0; // @[Map2T.scala 16:11]
  assign op_I1_5_0_0 = I1_5_0_0; // @[Map2T.scala 16:11]
  assign op_I1_6_0_0 = I1_6_0_0; // @[Map2T.scala 16:11]
  assign op_I1_7_0_0 = I1_7_0_0; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0 = I0_0; // @[Tuple.scala 24:34]
  assign O_1 = I0_1; // @[Tuple.scala 24:34]
  assign O_2 = I1; // @[Tuple.scala 26:32]
endmodule
module Map2S_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I1_0,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2; // @[Map2S.scala 9:22]
  SSeqTupleAppender fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_0_2 = fst_op_O_2; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_0_0_1,
  input  [7:0] I1_0_0,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  Map2S_3 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I1_0(fst_op_I1_0),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_5(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0_0,
  input  [7:0] I0_0_0_0_1,
  input  [7:0] I0_1_0_0_0,
  input  [7:0] I0_1_0_0_1,
  input  [7:0] I0_2_0_0_0,
  input  [7:0] I0_2_0_0_1,
  input  [7:0] I0_3_0_0_0,
  input  [7:0] I0_3_0_0_1,
  input  [7:0] I0_4_0_0_0,
  input  [7:0] I0_4_0_0_1,
  input  [7:0] I0_5_0_0_0,
  input  [7:0] I0_5_0_0_1,
  input  [7:0] I0_6_0_0_0,
  input  [7:0] I0_6_0_0_1,
  input  [7:0] I0_7_0_0_0,
  input  [7:0] I0_7_0_0_1,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_7_0_0,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_0_2,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_0_2,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_0_2,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_0_2,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_0_2,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_0_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  Map2S_4 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0_0(fst_op_I0_0_0_0),
    .I0_0_0_1(fst_op_I0_0_0_1),
    .I1_0_0(fst_op_I1_0_0),
    .O_0_0_0(fst_op_O_0_0_0),
    .O_0_0_1(fst_op_O_0_0_1),
    .O_0_0_2(fst_op_O_0_0_2)
  );
  Map2S_4 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0_0(other_ops_0_I0_0_0_0),
    .I0_0_0_1(other_ops_0_I0_0_0_1),
    .I1_0_0(other_ops_0_I1_0_0),
    .O_0_0_0(other_ops_0_O_0_0_0),
    .O_0_0_1(other_ops_0_O_0_0_1),
    .O_0_0_2(other_ops_0_O_0_0_2)
  );
  Map2S_4 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0_0(other_ops_1_I0_0_0_0),
    .I0_0_0_1(other_ops_1_I0_0_0_1),
    .I1_0_0(other_ops_1_I1_0_0),
    .O_0_0_0(other_ops_1_O_0_0_0),
    .O_0_0_1(other_ops_1_O_0_0_1),
    .O_0_0_2(other_ops_1_O_0_0_2)
  );
  Map2S_4 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0_0(other_ops_2_I0_0_0_0),
    .I0_0_0_1(other_ops_2_I0_0_0_1),
    .I1_0_0(other_ops_2_I1_0_0),
    .O_0_0_0(other_ops_2_O_0_0_0),
    .O_0_0_1(other_ops_2_O_0_0_1),
    .O_0_0_2(other_ops_2_O_0_0_2)
  );
  Map2S_4 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0_0(other_ops_3_I0_0_0_0),
    .I0_0_0_1(other_ops_3_I0_0_0_1),
    .I1_0_0(other_ops_3_I1_0_0),
    .O_0_0_0(other_ops_3_O_0_0_0),
    .O_0_0_1(other_ops_3_O_0_0_1),
    .O_0_0_2(other_ops_3_O_0_0_2)
  );
  Map2S_4 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0_0(other_ops_4_I0_0_0_0),
    .I0_0_0_1(other_ops_4_I0_0_0_1),
    .I1_0_0(other_ops_4_I1_0_0),
    .O_0_0_0(other_ops_4_O_0_0_0),
    .O_0_0_1(other_ops_4_O_0_0_1),
    .O_0_0_2(other_ops_4_O_0_0_2)
  );
  Map2S_4 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0_0(other_ops_5_I0_0_0_0),
    .I0_0_0_1(other_ops_5_I0_0_0_1),
    .I1_0_0(other_ops_5_I1_0_0),
    .O_0_0_0(other_ops_5_O_0_0_0),
    .O_0_0_1(other_ops_5_O_0_0_1),
    .O_0_0_2(other_ops_5_O_0_0_2)
  );
  Map2S_4 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0_0(other_ops_6_I0_0_0_0),
    .I0_0_0_1(other_ops_6_I0_0_0_1),
    .I1_0_0(other_ops_6_I1_0_0),
    .O_0_0_0(other_ops_6_O_0_0_0),
    .O_0_0_1(other_ops_6_O_0_0_1),
    .O_0_0_2(other_ops_6_O_0_0_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0_0 = fst_op_O_0_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_0_1 = fst_op_O_0_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_0_2 = fst_op_O_0_0_2; // @[Map2S.scala 19:8]
  assign O_1_0_0_0 = other_ops_0_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_0_1 = other_ops_0_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_0_2 = other_ops_0_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_2_0_0_0 = other_ops_1_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_0_1 = other_ops_1_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_0_2 = other_ops_1_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_3_0_0_0 = other_ops_2_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_0_1 = other_ops_2_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_0_2 = other_ops_2_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_4_0_0_0 = other_ops_3_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_0_1 = other_ops_3_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_0_2 = other_ops_3_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_5_0_0_0 = other_ops_4_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_0_1 = other_ops_4_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_0_2 = other_ops_4_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_6_0_0_0 = other_ops_5_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_0_1 = other_ops_5_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_0_2 = other_ops_5_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_7_0_0_0 = other_ops_6_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_0_1 = other_ops_6_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_0_2 = other_ops_6_O_0_0_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0_0 = I0_0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_0_1 = I0_0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_0 = I1_0_0_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0_0 = I0_1_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_0_1 = I0_1_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0_0 = I1_1_0_0; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0_0 = I0_2_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_0_1 = I0_2_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0_0 = I1_2_0_0; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0_0 = I0_3_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_0_1 = I0_3_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0_0 = I1_3_0_0; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0_0 = I0_4_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_0_1 = I0_4_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0_0 = I1_4_0_0; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0_0 = I0_5_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_0_1 = I0_5_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0_0 = I1_5_0_0; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0_0 = I0_6_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_0_1 = I0_6_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0_0 = I1_6_0_0; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0_0 = I0_7_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_0_1 = I0_7_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0_0 = I1_7_0_0; // @[Map2S.scala 23:43]
endmodule
module Map2T_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0_0,
  input  [7:0] I0_0_0_0_1,
  input  [7:0] I0_1_0_0_0,
  input  [7:0] I0_1_0_0_1,
  input  [7:0] I0_2_0_0_0,
  input  [7:0] I0_2_0_0_1,
  input  [7:0] I0_3_0_0_0,
  input  [7:0] I0_3_0_0_1,
  input  [7:0] I0_4_0_0_0,
  input  [7:0] I0_4_0_0_1,
  input  [7:0] I0_5_0_0_0,
  input  [7:0] I0_5_0_0_1,
  input  [7:0] I0_6_0_0_0,
  input  [7:0] I0_6_0_0_1,
  input  [7:0] I0_7_0_0_0,
  input  [7:0] I0_7_0_0_1,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_7_0_0,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_0_2,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_0_2,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_0_2,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_0_2,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_0_2,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_0_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_2; // @[Map2T.scala 8:20]
  Map2S_5 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0_0(op_I0_0_0_0_0),
    .I0_0_0_0_1(op_I0_0_0_0_1),
    .I0_1_0_0_0(op_I0_1_0_0_0),
    .I0_1_0_0_1(op_I0_1_0_0_1),
    .I0_2_0_0_0(op_I0_2_0_0_0),
    .I0_2_0_0_1(op_I0_2_0_0_1),
    .I0_3_0_0_0(op_I0_3_0_0_0),
    .I0_3_0_0_1(op_I0_3_0_0_1),
    .I0_4_0_0_0(op_I0_4_0_0_0),
    .I0_4_0_0_1(op_I0_4_0_0_1),
    .I0_5_0_0_0(op_I0_5_0_0_0),
    .I0_5_0_0_1(op_I0_5_0_0_1),
    .I0_6_0_0_0(op_I0_6_0_0_0),
    .I0_6_0_0_1(op_I0_6_0_0_1),
    .I0_7_0_0_0(op_I0_7_0_0_0),
    .I0_7_0_0_1(op_I0_7_0_0_1),
    .I1_0_0_0(op_I1_0_0_0),
    .I1_1_0_0(op_I1_1_0_0),
    .I1_2_0_0(op_I1_2_0_0),
    .I1_3_0_0(op_I1_3_0_0),
    .I1_4_0_0(op_I1_4_0_0),
    .I1_5_0_0(op_I1_5_0_0),
    .I1_6_0_0(op_I1_6_0_0),
    .I1_7_0_0(op_I1_7_0_0),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_0_0_0_2(op_O_0_0_0_2),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_1_0_0_2(op_O_1_0_0_2),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_2_0_0_2(op_O_2_0_0_2),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_3_0_0_2(op_O_3_0_0_2),
    .O_4_0_0_0(op_O_4_0_0_0),
    .O_4_0_0_1(op_O_4_0_0_1),
    .O_4_0_0_2(op_O_4_0_0_2),
    .O_5_0_0_0(op_O_5_0_0_0),
    .O_5_0_0_1(op_O_5_0_0_1),
    .O_5_0_0_2(op_O_5_0_0_2),
    .O_6_0_0_0(op_O_6_0_0_0),
    .O_6_0_0_1(op_O_6_0_0_1),
    .O_6_0_0_2(op_O_6_0_0_2),
    .O_7_0_0_0(op_O_7_0_0_0),
    .O_7_0_0_1(op_O_7_0_0_1),
    .O_7_0_0_2(op_O_7_0_0_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_0_2 = op_O_0_0_0_2; // @[Map2T.scala 17:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_0_2 = op_O_1_0_0_2; // @[Map2T.scala 17:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_0_2 = op_O_2_0_0_2; // @[Map2T.scala 17:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_0_2 = op_O_3_0_0_2; // @[Map2T.scala 17:7]
  assign O_4_0_0_0 = op_O_4_0_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_0_1 = op_O_4_0_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_0_2 = op_O_4_0_0_2; // @[Map2T.scala 17:7]
  assign O_5_0_0_0 = op_O_5_0_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_0_1 = op_O_5_0_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_0_2 = op_O_5_0_0_2; // @[Map2T.scala 17:7]
  assign O_6_0_0_0 = op_O_6_0_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_0_1 = op_O_6_0_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_0_2 = op_O_6_0_0_2; // @[Map2T.scala 17:7]
  assign O_7_0_0_0 = op_O_7_0_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_0_1 = op_O_7_0_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_0_2 = op_O_7_0_0_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0_0 = I0_0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_0_1 = I0_0_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0_0 = I0_1_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0_1 = I0_1_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0_0 = I0_2_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0_1 = I0_2_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0_0 = I0_3_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0_1 = I0_3_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0_0 = I0_4_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0_1 = I0_4_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0_0 = I0_5_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0_1 = I0_5_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0_0 = I0_6_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0_1 = I0_6_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0_0 = I0_7_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0_1 = I0_7_0_0_1; // @[Map2T.scala 15:11]
  assign op_I1_0_0_0 = I1_0_0_0; // @[Map2T.scala 16:11]
  assign op_I1_1_0_0 = I1_1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_2_0_0 = I1_2_0_0; // @[Map2T.scala 16:11]
  assign op_I1_3_0_0 = I1_3_0_0; // @[Map2T.scala 16:11]
  assign op_I1_4_0_0 = I1_4_0_0; // @[Map2T.scala 16:11]
  assign op_I1_5_0_0 = I1_5_0_0; // @[Map2T.scala 16:11]
  assign op_I1_6_0_0 = I1_6_0_0; // @[Map2T.scala 16:11]
  assign op_I1_7_0_0 = I1_7_0_0; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleToSSeq(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0 = I_0; // @[Tuple.scala 41:5]
  assign O_1 = I_1; // @[Tuple.scala 41:5]
  assign O_2 = I_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0(op_inst_I_0),
    .I_1(op_inst_I_1),
    .I_2(op_inst_I_2),
    .O_0(op_inst_O_0),
    .O_1(op_inst_O_1),
    .O_2(op_inst_O_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0 = op_inst_O_0; // @[Remove1S.scala 14:5]
  assign O_1 = op_inst_O_1; // @[Remove1S.scala 14:5]
  assign O_2 = op_inst_O_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0 = I_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1 = I_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2 = I_0_2; // @[Remove1S.scala 13:13]
endmodule
module MapS(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2; // @[MapS.scala 9:22]
  Remove1S fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
endmodule
module MapS_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0_0,
  input  [7:0] I_0_0_0_1,
  input  [7:0] I_0_0_0_2,
  input  [7:0] I_1_0_0_0,
  input  [7:0] I_1_0_0_1,
  input  [7:0] I_1_0_0_2,
  input  [7:0] I_2_0_0_0,
  input  [7:0] I_2_0_0_1,
  input  [7:0] I_2_0_0_2,
  input  [7:0] I_3_0_0_0,
  input  [7:0] I_3_0_0_1,
  input  [7:0] I_3_0_0_2,
  input  [7:0] I_4_0_0_0,
  input  [7:0] I_4_0_0_1,
  input  [7:0] I_4_0_0_2,
  input  [7:0] I_5_0_0_0,
  input  [7:0] I_5_0_0_1,
  input  [7:0] I_5_0_0_2,
  input  [7:0] I_6_0_0_0,
  input  [7:0] I_6_0_0_1,
  input  [7:0] I_6_0_0_2,
  input  [7:0] I_7_0_0_0,
  input  [7:0] I_7_0_0_1,
  input  [7:0] I_7_0_0_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  MapS fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0_0(fst_op_I_0_0_0),
    .I_0_0_1(fst_op_I_0_0_1),
    .I_0_0_2(fst_op_I_0_0_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2)
  );
  MapS other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0_0(other_ops_0_I_0_0_0),
    .I_0_0_1(other_ops_0_I_0_0_1),
    .I_0_0_2(other_ops_0_I_0_0_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2)
  );
  MapS other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0_0(other_ops_1_I_0_0_0),
    .I_0_0_1(other_ops_1_I_0_0_1),
    .I_0_0_2(other_ops_1_I_0_0_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2)
  );
  MapS other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0_0(other_ops_2_I_0_0_0),
    .I_0_0_1(other_ops_2_I_0_0_1),
    .I_0_0_2(other_ops_2_I_0_0_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2)
  );
  MapS other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0_0(other_ops_3_I_0_0_0),
    .I_0_0_1(other_ops_3_I_0_0_1),
    .I_0_0_2(other_ops_3_I_0_0_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2)
  );
  MapS other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0_0(other_ops_4_I_0_0_0),
    .I_0_0_1(other_ops_4_I_0_0_1),
    .I_0_0_2(other_ops_4_I_0_0_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2)
  );
  MapS other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0_0(other_ops_5_I_0_0_0),
    .I_0_0_1(other_ops_5_I_0_0_1),
    .I_0_0_2(other_ops_5_I_0_0_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2)
  );
  MapS other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0_0(other_ops_6_I_0_0_0),
    .I_0_0_1(other_ops_6_I_0_0_1),
    .I_0_0_2(other_ops_6_I_0_0_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[MapS.scala 17:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[MapS.scala 21:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[MapS.scala 21:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[MapS.scala 21:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[MapS.scala 21:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[MapS.scala 21:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[MapS.scala 21:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[MapS.scala 21:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0_0 = I_0_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_1 = I_0_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_2 = I_0_0_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0_0 = I_1_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_1 = I_1_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_2 = I_1_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0_0 = I_2_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_1 = I_2_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_2 = I_2_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0_0 = I_3_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_1 = I_3_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_2 = I_3_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0_0 = I_4_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_1 = I_4_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_2 = I_4_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0_0 = I_5_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_1 = I_5_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_2 = I_5_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0_0 = I_6_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_1 = I_6_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_2 = I_6_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0_0 = I_7_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_1 = I_7_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_2 = I_7_0_0_2; // @[MapS.scala 20:41]
endmodule
module MapT(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0_0,
  input  [7:0] I_0_0_0_1,
  input  [7:0] I_0_0_0_2,
  input  [7:0] I_1_0_0_0,
  input  [7:0] I_1_0_0_1,
  input  [7:0] I_1_0_0_2,
  input  [7:0] I_2_0_0_0,
  input  [7:0] I_2_0_0_1,
  input  [7:0] I_2_0_0_2,
  input  [7:0] I_3_0_0_0,
  input  [7:0] I_3_0_0_1,
  input  [7:0] I_3_0_0_2,
  input  [7:0] I_4_0_0_0,
  input  [7:0] I_4_0_0_1,
  input  [7:0] I_4_0_0_2,
  input  [7:0] I_5_0_0_0,
  input  [7:0] I_5_0_0_1,
  input  [7:0] I_5_0_0_2,
  input  [7:0] I_6_0_0_0,
  input  [7:0] I_6_0_0_1,
  input  [7:0] I_6_0_0_2,
  input  [7:0] I_7_0_0_0,
  input  [7:0] I_7_0_0_1,
  input  [7:0] I_7_0_0_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_2; // @[MapT.scala 8:20]
  MapS_1 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0_0(op_I_0_0_0_0),
    .I_0_0_0_1(op_I_0_0_0_1),
    .I_0_0_0_2(op_I_0_0_0_2),
    .I_1_0_0_0(op_I_1_0_0_0),
    .I_1_0_0_1(op_I_1_0_0_1),
    .I_1_0_0_2(op_I_1_0_0_2),
    .I_2_0_0_0(op_I_2_0_0_0),
    .I_2_0_0_1(op_I_2_0_0_1),
    .I_2_0_0_2(op_I_2_0_0_2),
    .I_3_0_0_0(op_I_3_0_0_0),
    .I_3_0_0_1(op_I_3_0_0_1),
    .I_3_0_0_2(op_I_3_0_0_2),
    .I_4_0_0_0(op_I_4_0_0_0),
    .I_4_0_0_1(op_I_4_0_0_1),
    .I_4_0_0_2(op_I_4_0_0_2),
    .I_5_0_0_0(op_I_5_0_0_0),
    .I_5_0_0_1(op_I_5_0_0_1),
    .I_5_0_0_2(op_I_5_0_0_2),
    .I_6_0_0_0(op_I_6_0_0_0),
    .I_6_0_0_1(op_I_6_0_0_1),
    .I_6_0_0_2(op_I_6_0_0_2),
    .I_7_0_0_0(op_I_7_0_0_0),
    .I_7_0_0_1(op_I_7_0_0_1),
    .I_7_0_0_2(op_I_7_0_0_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_4_0_2 = op_O_4_0_2; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_5_0_2 = op_O_5_0_2; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_6_0_2 = op_O_6_0_2; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_7_0_2 = op_O_7_0_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0_0 = I_0_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_0_1 = I_0_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_0_2 = I_0_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0_0 = I_1_0_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_0_1 = I_1_0_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0_2 = I_1_0_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0_0 = I_2_0_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_0_1 = I_2_0_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0_2 = I_2_0_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0_0 = I_3_0_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_0_1 = I_3_0_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0_2 = I_3_0_0_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0_0 = I_4_0_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_0_1 = I_4_0_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_0_2 = I_4_0_0_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0_0 = I_5_0_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_0_1 = I_5_0_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_0_2 = I_5_0_0_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0_0 = I_6_0_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_0_1 = I_6_0_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_0_2 = I_6_0_0_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0_0 = I_7_0_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_0_1 = I_7_0_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_0_2 = I_7_0_0_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleCreator_2(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0_0 = I0_0; // @[Tuple.scala 12:32]
  assign O_0_1 = I0_1; // @[Tuple.scala 12:32]
  assign O_0_2 = I0_2; // @[Tuple.scala 12:32]
  assign O_1_0 = I1_0; // @[Tuple.scala 13:32]
  assign O_1_1 = I1_1; // @[Tuple.scala 13:32]
  assign O_1_2 = I1_2; // @[Tuple.scala 13:32]
endmodule
module Map2S_12(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_0_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  SSeqTupleCreator_2 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
endmodule
module Map2S_13(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_0_0_1,
  input  [7:0] I0_0_0_2,
  input  [7:0] I0_1_0_0,
  input  [7:0] I0_1_0_1,
  input  [7:0] I0_1_0_2,
  input  [7:0] I0_2_0_0,
  input  [7:0] I0_2_0_1,
  input  [7:0] I0_2_0_2,
  input  [7:0] I0_3_0_0,
  input  [7:0] I0_3_0_1,
  input  [7:0] I0_3_0_2,
  input  [7:0] I0_4_0_0,
  input  [7:0] I0_4_0_1,
  input  [7:0] I0_4_0_2,
  input  [7:0] I0_5_0_0,
  input  [7:0] I0_5_0_1,
  input  [7:0] I0_5_0_2,
  input  [7:0] I0_6_0_0,
  input  [7:0] I0_6_0_1,
  input  [7:0] I0_6_0_2,
  input  [7:0] I0_7_0_0,
  input  [7:0] I0_7_0_1,
  input  [7:0] I0_7_0_2,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_0_0_1,
  input  [7:0] I1_0_0_2,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_1_0_1,
  input  [7:0] I1_1_0_2,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_2_0_1,
  input  [7:0] I1_2_0_2,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_3_0_1,
  input  [7:0] I1_3_0_2,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_4_0_1,
  input  [7:0] I1_4_0_2,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_5_0_1,
  input  [7:0] I1_5_0_2,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_6_0_1,
  input  [7:0] I1_6_0_2,
  input  [7:0] I1_7_0_0,
  input  [7:0] I1_7_0_1,
  input  [7:0] I1_7_0_2,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_0_0_1_0,
  output [7:0] O_0_0_1_1,
  output [7:0] O_0_0_1_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_1_0_1_0,
  output [7:0] O_1_0_1_1,
  output [7:0] O_1_0_1_2,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_0_2,
  output [7:0] O_2_0_1_0,
  output [7:0] O_2_0_1_1,
  output [7:0] O_2_0_1_2,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_0_2,
  output [7:0] O_3_0_1_0,
  output [7:0] O_3_0_1_1,
  output [7:0] O_3_0_1_2,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_0_2,
  output [7:0] O_4_0_1_0,
  output [7:0] O_4_0_1_1,
  output [7:0] O_4_0_1_2,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_0_2,
  output [7:0] O_5_0_1_0,
  output [7:0] O_5_0_1_1,
  output [7:0] O_5_0_1_2,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_0_2,
  output [7:0] O_6_0_1_0,
  output [7:0] O_6_0_1_1,
  output [7:0] O_6_0_1_2,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_0_2,
  output [7:0] O_7_0_1_0,
  output [7:0] O_7_0_1_1,
  output [7:0] O_7_0_1_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  Map2S_12 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I1_0_0(fst_op_I1_0_0),
    .I1_0_1(fst_op_I1_0_1),
    .I1_0_2(fst_op_I1_0_2),
    .O_0_0_0(fst_op_O_0_0_0),
    .O_0_0_1(fst_op_O_0_0_1),
    .O_0_0_2(fst_op_O_0_0_2),
    .O_0_1_0(fst_op_O_0_1_0),
    .O_0_1_1(fst_op_O_0_1_1),
    .O_0_1_2(fst_op_O_0_1_2)
  );
  Map2S_12 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0(other_ops_0_I0_0_0),
    .I0_0_1(other_ops_0_I0_0_1),
    .I0_0_2(other_ops_0_I0_0_2),
    .I1_0_0(other_ops_0_I1_0_0),
    .I1_0_1(other_ops_0_I1_0_1),
    .I1_0_2(other_ops_0_I1_0_2),
    .O_0_0_0(other_ops_0_O_0_0_0),
    .O_0_0_1(other_ops_0_O_0_0_1),
    .O_0_0_2(other_ops_0_O_0_0_2),
    .O_0_1_0(other_ops_0_O_0_1_0),
    .O_0_1_1(other_ops_0_O_0_1_1),
    .O_0_1_2(other_ops_0_O_0_1_2)
  );
  Map2S_12 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0(other_ops_1_I0_0_0),
    .I0_0_1(other_ops_1_I0_0_1),
    .I0_0_2(other_ops_1_I0_0_2),
    .I1_0_0(other_ops_1_I1_0_0),
    .I1_0_1(other_ops_1_I1_0_1),
    .I1_0_2(other_ops_1_I1_0_2),
    .O_0_0_0(other_ops_1_O_0_0_0),
    .O_0_0_1(other_ops_1_O_0_0_1),
    .O_0_0_2(other_ops_1_O_0_0_2),
    .O_0_1_0(other_ops_1_O_0_1_0),
    .O_0_1_1(other_ops_1_O_0_1_1),
    .O_0_1_2(other_ops_1_O_0_1_2)
  );
  Map2S_12 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0(other_ops_2_I0_0_0),
    .I0_0_1(other_ops_2_I0_0_1),
    .I0_0_2(other_ops_2_I0_0_2),
    .I1_0_0(other_ops_2_I1_0_0),
    .I1_0_1(other_ops_2_I1_0_1),
    .I1_0_2(other_ops_2_I1_0_2),
    .O_0_0_0(other_ops_2_O_0_0_0),
    .O_0_0_1(other_ops_2_O_0_0_1),
    .O_0_0_2(other_ops_2_O_0_0_2),
    .O_0_1_0(other_ops_2_O_0_1_0),
    .O_0_1_1(other_ops_2_O_0_1_1),
    .O_0_1_2(other_ops_2_O_0_1_2)
  );
  Map2S_12 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0(other_ops_3_I0_0_0),
    .I0_0_1(other_ops_3_I0_0_1),
    .I0_0_2(other_ops_3_I0_0_2),
    .I1_0_0(other_ops_3_I1_0_0),
    .I1_0_1(other_ops_3_I1_0_1),
    .I1_0_2(other_ops_3_I1_0_2),
    .O_0_0_0(other_ops_3_O_0_0_0),
    .O_0_0_1(other_ops_3_O_0_0_1),
    .O_0_0_2(other_ops_3_O_0_0_2),
    .O_0_1_0(other_ops_3_O_0_1_0),
    .O_0_1_1(other_ops_3_O_0_1_1),
    .O_0_1_2(other_ops_3_O_0_1_2)
  );
  Map2S_12 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0(other_ops_4_I0_0_0),
    .I0_0_1(other_ops_4_I0_0_1),
    .I0_0_2(other_ops_4_I0_0_2),
    .I1_0_0(other_ops_4_I1_0_0),
    .I1_0_1(other_ops_4_I1_0_1),
    .I1_0_2(other_ops_4_I1_0_2),
    .O_0_0_0(other_ops_4_O_0_0_0),
    .O_0_0_1(other_ops_4_O_0_0_1),
    .O_0_0_2(other_ops_4_O_0_0_2),
    .O_0_1_0(other_ops_4_O_0_1_0),
    .O_0_1_1(other_ops_4_O_0_1_1),
    .O_0_1_2(other_ops_4_O_0_1_2)
  );
  Map2S_12 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0(other_ops_5_I0_0_0),
    .I0_0_1(other_ops_5_I0_0_1),
    .I0_0_2(other_ops_5_I0_0_2),
    .I1_0_0(other_ops_5_I1_0_0),
    .I1_0_1(other_ops_5_I1_0_1),
    .I1_0_2(other_ops_5_I1_0_2),
    .O_0_0_0(other_ops_5_O_0_0_0),
    .O_0_0_1(other_ops_5_O_0_0_1),
    .O_0_0_2(other_ops_5_O_0_0_2),
    .O_0_1_0(other_ops_5_O_0_1_0),
    .O_0_1_1(other_ops_5_O_0_1_1),
    .O_0_1_2(other_ops_5_O_0_1_2)
  );
  Map2S_12 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0(other_ops_6_I0_0_0),
    .I0_0_1(other_ops_6_I0_0_1),
    .I0_0_2(other_ops_6_I0_0_2),
    .I1_0_0(other_ops_6_I1_0_0),
    .I1_0_1(other_ops_6_I1_0_1),
    .I1_0_2(other_ops_6_I1_0_2),
    .O_0_0_0(other_ops_6_O_0_0_0),
    .O_0_0_1(other_ops_6_O_0_0_1),
    .O_0_0_2(other_ops_6_O_0_0_2),
    .O_0_1_0(other_ops_6_O_0_1_0),
    .O_0_1_1(other_ops_6_O_0_1_1),
    .O_0_1_2(other_ops_6_O_0_1_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0_0 = fst_op_O_0_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_0_1 = fst_op_O_0_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_0_2 = fst_op_O_0_0_2; // @[Map2S.scala 19:8]
  assign O_0_0_1_0 = fst_op_O_0_1_0; // @[Map2S.scala 19:8]
  assign O_0_0_1_1 = fst_op_O_0_1_1; // @[Map2S.scala 19:8]
  assign O_0_0_1_2 = fst_op_O_0_1_2; // @[Map2S.scala 19:8]
  assign O_1_0_0_0 = other_ops_0_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_0_1 = other_ops_0_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_0_2 = other_ops_0_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_1_0_1_0 = other_ops_0_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_1_0_1_1 = other_ops_0_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_1_0_1_2 = other_ops_0_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_2_0_0_0 = other_ops_1_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_0_1 = other_ops_1_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_0_2 = other_ops_1_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_2_0_1_0 = other_ops_1_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_2_0_1_1 = other_ops_1_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_2_0_1_2 = other_ops_1_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_3_0_0_0 = other_ops_2_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_0_1 = other_ops_2_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_0_2 = other_ops_2_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_3_0_1_0 = other_ops_2_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_3_0_1_1 = other_ops_2_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_3_0_1_2 = other_ops_2_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_4_0_0_0 = other_ops_3_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_0_1 = other_ops_3_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_0_2 = other_ops_3_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_4_0_1_0 = other_ops_3_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_4_0_1_1 = other_ops_3_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_4_0_1_2 = other_ops_3_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_5_0_0_0 = other_ops_4_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_0_1 = other_ops_4_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_0_2 = other_ops_4_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_5_0_1_0 = other_ops_4_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_5_0_1_1 = other_ops_4_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_5_0_1_2 = other_ops_4_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_6_0_0_0 = other_ops_5_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_0_1 = other_ops_5_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_0_2 = other_ops_5_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_6_0_1_0 = other_ops_5_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_6_0_1_1 = other_ops_5_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_6_0_1_2 = other_ops_5_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_7_0_0_0 = other_ops_6_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_0_1 = other_ops_6_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_0_2 = other_ops_6_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_7_0_1_0 = other_ops_6_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_7_0_1_1 = other_ops_6_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_7_0_1_2 = other_ops_6_O_0_1_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_0 = I1_0_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_1 = I1_0_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_2 = I1_0_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0 = I0_1_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1 = I0_1_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_2 = I0_1_0_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0_0 = I1_1_0_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_0_1 = I1_1_0_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_0_2 = I1_1_0_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0 = I0_2_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1 = I0_2_0_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_2 = I0_2_0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0_0 = I1_2_0_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_0_1 = I1_2_0_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_0_2 = I1_2_0_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0 = I0_3_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1 = I0_3_0_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_2 = I0_3_0_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0_0 = I1_3_0_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_0_1 = I1_3_0_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_0_2 = I1_3_0_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0 = I0_4_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1 = I0_4_0_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_2 = I0_4_0_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0_0 = I1_4_0_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_0_1 = I1_4_0_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_0_2 = I1_4_0_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0 = I0_5_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1 = I0_5_0_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_2 = I0_5_0_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0_0 = I1_5_0_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_0_1 = I1_5_0_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_0_2 = I1_5_0_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0 = I0_6_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1 = I0_6_0_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_2 = I0_6_0_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0_0 = I1_6_0_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_0_1 = I1_6_0_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_0_2 = I1_6_0_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0 = I0_7_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1 = I0_7_0_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_2 = I0_7_0_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0_0 = I1_7_0_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_0_1 = I1_7_0_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_0_2 = I1_7_0_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_0_0_1,
  input  [7:0] I0_0_0_2,
  input  [7:0] I0_1_0_0,
  input  [7:0] I0_1_0_1,
  input  [7:0] I0_1_0_2,
  input  [7:0] I0_2_0_0,
  input  [7:0] I0_2_0_1,
  input  [7:0] I0_2_0_2,
  input  [7:0] I0_3_0_0,
  input  [7:0] I0_3_0_1,
  input  [7:0] I0_3_0_2,
  input  [7:0] I0_4_0_0,
  input  [7:0] I0_4_0_1,
  input  [7:0] I0_4_0_2,
  input  [7:0] I0_5_0_0,
  input  [7:0] I0_5_0_1,
  input  [7:0] I0_5_0_2,
  input  [7:0] I0_6_0_0,
  input  [7:0] I0_6_0_1,
  input  [7:0] I0_6_0_2,
  input  [7:0] I0_7_0_0,
  input  [7:0] I0_7_0_1,
  input  [7:0] I0_7_0_2,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_0_0_1,
  input  [7:0] I1_0_0_2,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_1_0_1,
  input  [7:0] I1_1_0_2,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_2_0_1,
  input  [7:0] I1_2_0_2,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_3_0_1,
  input  [7:0] I1_3_0_2,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_4_0_1,
  input  [7:0] I1_4_0_2,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_5_0_1,
  input  [7:0] I1_5_0_2,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_6_0_1,
  input  [7:0] I1_6_0_2,
  input  [7:0] I1_7_0_0,
  input  [7:0] I1_7_0_1,
  input  [7:0] I1_7_0_2,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_0_0_1_0,
  output [7:0] O_0_0_1_1,
  output [7:0] O_0_0_1_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_1_0_1_0,
  output [7:0] O_1_0_1_1,
  output [7:0] O_1_0_1_2,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_0_2,
  output [7:0] O_2_0_1_0,
  output [7:0] O_2_0_1_1,
  output [7:0] O_2_0_1_2,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_0_2,
  output [7:0] O_3_0_1_0,
  output [7:0] O_3_0_1_1,
  output [7:0] O_3_0_1_2,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_0_2,
  output [7:0] O_4_0_1_0,
  output [7:0] O_4_0_1_1,
  output [7:0] O_4_0_1_2,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_0_2,
  output [7:0] O_5_0_1_0,
  output [7:0] O_5_0_1_1,
  output [7:0] O_5_0_1_2,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_0_2,
  output [7:0] O_6_0_1_0,
  output [7:0] O_6_0_1_1,
  output [7:0] O_6_0_1_2,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_0_2,
  output [7:0] O_7_0_1_0,
  output [7:0] O_7_0_1_1,
  output [7:0] O_7_0_1_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_1_2; // @[Map2T.scala 8:20]
  Map2S_13 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0(op_I0_0_0_0),
    .I0_0_0_1(op_I0_0_0_1),
    .I0_0_0_2(op_I0_0_0_2),
    .I0_1_0_0(op_I0_1_0_0),
    .I0_1_0_1(op_I0_1_0_1),
    .I0_1_0_2(op_I0_1_0_2),
    .I0_2_0_0(op_I0_2_0_0),
    .I0_2_0_1(op_I0_2_0_1),
    .I0_2_0_2(op_I0_2_0_2),
    .I0_3_0_0(op_I0_3_0_0),
    .I0_3_0_1(op_I0_3_0_1),
    .I0_3_0_2(op_I0_3_0_2),
    .I0_4_0_0(op_I0_4_0_0),
    .I0_4_0_1(op_I0_4_0_1),
    .I0_4_0_2(op_I0_4_0_2),
    .I0_5_0_0(op_I0_5_0_0),
    .I0_5_0_1(op_I0_5_0_1),
    .I0_5_0_2(op_I0_5_0_2),
    .I0_6_0_0(op_I0_6_0_0),
    .I0_6_0_1(op_I0_6_0_1),
    .I0_6_0_2(op_I0_6_0_2),
    .I0_7_0_0(op_I0_7_0_0),
    .I0_7_0_1(op_I0_7_0_1),
    .I0_7_0_2(op_I0_7_0_2),
    .I1_0_0_0(op_I1_0_0_0),
    .I1_0_0_1(op_I1_0_0_1),
    .I1_0_0_2(op_I1_0_0_2),
    .I1_1_0_0(op_I1_1_0_0),
    .I1_1_0_1(op_I1_1_0_1),
    .I1_1_0_2(op_I1_1_0_2),
    .I1_2_0_0(op_I1_2_0_0),
    .I1_2_0_1(op_I1_2_0_1),
    .I1_2_0_2(op_I1_2_0_2),
    .I1_3_0_0(op_I1_3_0_0),
    .I1_3_0_1(op_I1_3_0_1),
    .I1_3_0_2(op_I1_3_0_2),
    .I1_4_0_0(op_I1_4_0_0),
    .I1_4_0_1(op_I1_4_0_1),
    .I1_4_0_2(op_I1_4_0_2),
    .I1_5_0_0(op_I1_5_0_0),
    .I1_5_0_1(op_I1_5_0_1),
    .I1_5_0_2(op_I1_5_0_2),
    .I1_6_0_0(op_I1_6_0_0),
    .I1_6_0_1(op_I1_6_0_1),
    .I1_6_0_2(op_I1_6_0_2),
    .I1_7_0_0(op_I1_7_0_0),
    .I1_7_0_1(op_I1_7_0_1),
    .I1_7_0_2(op_I1_7_0_2),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_0_0_0_2(op_O_0_0_0_2),
    .O_0_0_1_0(op_O_0_0_1_0),
    .O_0_0_1_1(op_O_0_0_1_1),
    .O_0_0_1_2(op_O_0_0_1_2),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_1_0_0_2(op_O_1_0_0_2),
    .O_1_0_1_0(op_O_1_0_1_0),
    .O_1_0_1_1(op_O_1_0_1_1),
    .O_1_0_1_2(op_O_1_0_1_2),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_2_0_0_2(op_O_2_0_0_2),
    .O_2_0_1_0(op_O_2_0_1_0),
    .O_2_0_1_1(op_O_2_0_1_1),
    .O_2_0_1_2(op_O_2_0_1_2),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_3_0_0_2(op_O_3_0_0_2),
    .O_3_0_1_0(op_O_3_0_1_0),
    .O_3_0_1_1(op_O_3_0_1_1),
    .O_3_0_1_2(op_O_3_0_1_2),
    .O_4_0_0_0(op_O_4_0_0_0),
    .O_4_0_0_1(op_O_4_0_0_1),
    .O_4_0_0_2(op_O_4_0_0_2),
    .O_4_0_1_0(op_O_4_0_1_0),
    .O_4_0_1_1(op_O_4_0_1_1),
    .O_4_0_1_2(op_O_4_0_1_2),
    .O_5_0_0_0(op_O_5_0_0_0),
    .O_5_0_0_1(op_O_5_0_0_1),
    .O_5_0_0_2(op_O_5_0_0_2),
    .O_5_0_1_0(op_O_5_0_1_0),
    .O_5_0_1_1(op_O_5_0_1_1),
    .O_5_0_1_2(op_O_5_0_1_2),
    .O_6_0_0_0(op_O_6_0_0_0),
    .O_6_0_0_1(op_O_6_0_0_1),
    .O_6_0_0_2(op_O_6_0_0_2),
    .O_6_0_1_0(op_O_6_0_1_0),
    .O_6_0_1_1(op_O_6_0_1_1),
    .O_6_0_1_2(op_O_6_0_1_2),
    .O_7_0_0_0(op_O_7_0_0_0),
    .O_7_0_0_1(op_O_7_0_0_1),
    .O_7_0_0_2(op_O_7_0_0_2),
    .O_7_0_1_0(op_O_7_0_1_0),
    .O_7_0_1_1(op_O_7_0_1_1),
    .O_7_0_1_2(op_O_7_0_1_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_0_2 = op_O_0_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_0_1_0 = op_O_0_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_0_1_1 = op_O_0_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_0_1_2 = op_O_0_0_1_2; // @[Map2T.scala 17:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_0_2 = op_O_1_0_0_2; // @[Map2T.scala 17:7]
  assign O_1_0_1_0 = op_O_1_0_1_0; // @[Map2T.scala 17:7]
  assign O_1_0_1_1 = op_O_1_0_1_1; // @[Map2T.scala 17:7]
  assign O_1_0_1_2 = op_O_1_0_1_2; // @[Map2T.scala 17:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_0_2 = op_O_2_0_0_2; // @[Map2T.scala 17:7]
  assign O_2_0_1_0 = op_O_2_0_1_0; // @[Map2T.scala 17:7]
  assign O_2_0_1_1 = op_O_2_0_1_1; // @[Map2T.scala 17:7]
  assign O_2_0_1_2 = op_O_2_0_1_2; // @[Map2T.scala 17:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_0_2 = op_O_3_0_0_2; // @[Map2T.scala 17:7]
  assign O_3_0_1_0 = op_O_3_0_1_0; // @[Map2T.scala 17:7]
  assign O_3_0_1_1 = op_O_3_0_1_1; // @[Map2T.scala 17:7]
  assign O_3_0_1_2 = op_O_3_0_1_2; // @[Map2T.scala 17:7]
  assign O_4_0_0_0 = op_O_4_0_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_0_1 = op_O_4_0_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_0_2 = op_O_4_0_0_2; // @[Map2T.scala 17:7]
  assign O_4_0_1_0 = op_O_4_0_1_0; // @[Map2T.scala 17:7]
  assign O_4_0_1_1 = op_O_4_0_1_1; // @[Map2T.scala 17:7]
  assign O_4_0_1_2 = op_O_4_0_1_2; // @[Map2T.scala 17:7]
  assign O_5_0_0_0 = op_O_5_0_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_0_1 = op_O_5_0_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_0_2 = op_O_5_0_0_2; // @[Map2T.scala 17:7]
  assign O_5_0_1_0 = op_O_5_0_1_0; // @[Map2T.scala 17:7]
  assign O_5_0_1_1 = op_O_5_0_1_1; // @[Map2T.scala 17:7]
  assign O_5_0_1_2 = op_O_5_0_1_2; // @[Map2T.scala 17:7]
  assign O_6_0_0_0 = op_O_6_0_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_0_1 = op_O_6_0_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_0_2 = op_O_6_0_0_2; // @[Map2T.scala 17:7]
  assign O_6_0_1_0 = op_O_6_0_1_0; // @[Map2T.scala 17:7]
  assign O_6_0_1_1 = op_O_6_0_1_1; // @[Map2T.scala 17:7]
  assign O_6_0_1_2 = op_O_6_0_1_2; // @[Map2T.scala 17:7]
  assign O_7_0_0_0 = op_O_7_0_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_0_1 = op_O_7_0_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_0_2 = op_O_7_0_0_2; // @[Map2T.scala 17:7]
  assign O_7_0_1_0 = op_O_7_0_1_0; // @[Map2T.scala 17:7]
  assign O_7_0_1_1 = op_O_7_0_1_1; // @[Map2T.scala 17:7]
  assign O_7_0_1_2 = op_O_7_0_1_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0 = I0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1 = I0_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_0_2 = I0_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0 = I0_1_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1 = I0_1_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_2 = I0_1_0_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0 = I0_2_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1 = I0_2_0_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_2 = I0_2_0_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0 = I0_3_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1 = I0_3_0_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_2 = I0_3_0_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0 = I0_4_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_1 = I0_4_0_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0_2 = I0_4_0_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0 = I0_5_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_1 = I0_5_0_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0_2 = I0_5_0_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0 = I0_6_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_1 = I0_6_0_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0_2 = I0_6_0_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0 = I0_7_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_1 = I0_7_0_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0_2 = I0_7_0_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0_0 = I1_0_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_0_1 = I1_0_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_0_2 = I1_0_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0_0 = I1_1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_1_0_1 = I1_1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_1_0_2 = I1_1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0_0 = I1_2_0_0; // @[Map2T.scala 16:11]
  assign op_I1_2_0_1 = I1_2_0_1; // @[Map2T.scala 16:11]
  assign op_I1_2_0_2 = I1_2_0_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0_0 = I1_3_0_0; // @[Map2T.scala 16:11]
  assign op_I1_3_0_1 = I1_3_0_1; // @[Map2T.scala 16:11]
  assign op_I1_3_0_2 = I1_3_0_2; // @[Map2T.scala 16:11]
  assign op_I1_4_0_0 = I1_4_0_0; // @[Map2T.scala 16:11]
  assign op_I1_4_0_1 = I1_4_0_1; // @[Map2T.scala 16:11]
  assign op_I1_4_0_2 = I1_4_0_2; // @[Map2T.scala 16:11]
  assign op_I1_5_0_0 = I1_5_0_0; // @[Map2T.scala 16:11]
  assign op_I1_5_0_1 = I1_5_0_1; // @[Map2T.scala 16:11]
  assign op_I1_5_0_2 = I1_5_0_2; // @[Map2T.scala 16:11]
  assign op_I1_6_0_0 = I1_6_0_0; // @[Map2T.scala 16:11]
  assign op_I1_6_0_1 = I1_6_0_1; // @[Map2T.scala 16:11]
  assign op_I1_6_0_2 = I1_6_0_2; // @[Map2T.scala 16:11]
  assign op_I1_7_0_0 = I1_7_0_0; // @[Map2T.scala 16:11]
  assign op_I1_7_0_1 = I1_7_0_1; // @[Map2T.scala 16:11]
  assign op_I1_7_0_2 = I1_7_0_2; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_1_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0_0 = I0_0_0; // @[Tuple.scala 24:34]
  assign O_0_1 = I0_0_1; // @[Tuple.scala 24:34]
  assign O_0_2 = I0_0_2; // @[Tuple.scala 24:34]
  assign O_1_0 = I0_1_0; // @[Tuple.scala 24:34]
  assign O_1_1 = I0_1_1; // @[Tuple.scala 24:34]
  assign O_1_2 = I0_1_2; // @[Tuple.scala 24:34]
  assign O_2_0 = I1_0; // @[Tuple.scala 26:32]
  assign O_2_1 = I1_1; // @[Tuple.scala 26:32]
  assign O_2_2 = I1_2; // @[Tuple.scala 26:32]
endmodule
module Map2S_20(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_0_0_1,
  input  [7:0] I0_0_0_2,
  input  [7:0] I0_0_1_0,
  input  [7:0] I0_0_1_1,
  input  [7:0] I0_0_1_2,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_0_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_2; // @[Map2S.scala 9:22]
  SSeqTupleAppender_3 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I0_1_0(fst_op_I0_1_0),
    .I0_1_1(fst_op_I0_1_1),
    .I0_1_2(fst_op_I0_1_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[Map2S.scala 19:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[Map2S.scala 19:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_0 = I0_0_1_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_1 = I0_0_1_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_2 = I0_0_1_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
endmodule
module Map2S_21(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0_0,
  input  [7:0] I0_0_0_0_1,
  input  [7:0] I0_0_0_0_2,
  input  [7:0] I0_0_0_1_0,
  input  [7:0] I0_0_0_1_1,
  input  [7:0] I0_0_0_1_2,
  input  [7:0] I0_1_0_0_0,
  input  [7:0] I0_1_0_0_1,
  input  [7:0] I0_1_0_0_2,
  input  [7:0] I0_1_0_1_0,
  input  [7:0] I0_1_0_1_1,
  input  [7:0] I0_1_0_1_2,
  input  [7:0] I0_2_0_0_0,
  input  [7:0] I0_2_0_0_1,
  input  [7:0] I0_2_0_0_2,
  input  [7:0] I0_2_0_1_0,
  input  [7:0] I0_2_0_1_1,
  input  [7:0] I0_2_0_1_2,
  input  [7:0] I0_3_0_0_0,
  input  [7:0] I0_3_0_0_1,
  input  [7:0] I0_3_0_0_2,
  input  [7:0] I0_3_0_1_0,
  input  [7:0] I0_3_0_1_1,
  input  [7:0] I0_3_0_1_2,
  input  [7:0] I0_4_0_0_0,
  input  [7:0] I0_4_0_0_1,
  input  [7:0] I0_4_0_0_2,
  input  [7:0] I0_4_0_1_0,
  input  [7:0] I0_4_0_1_1,
  input  [7:0] I0_4_0_1_2,
  input  [7:0] I0_5_0_0_0,
  input  [7:0] I0_5_0_0_1,
  input  [7:0] I0_5_0_0_2,
  input  [7:0] I0_5_0_1_0,
  input  [7:0] I0_5_0_1_1,
  input  [7:0] I0_5_0_1_2,
  input  [7:0] I0_6_0_0_0,
  input  [7:0] I0_6_0_0_1,
  input  [7:0] I0_6_0_0_2,
  input  [7:0] I0_6_0_1_0,
  input  [7:0] I0_6_0_1_1,
  input  [7:0] I0_6_0_1_2,
  input  [7:0] I0_7_0_0_0,
  input  [7:0] I0_7_0_0_1,
  input  [7:0] I0_7_0_0_2,
  input  [7:0] I0_7_0_1_0,
  input  [7:0] I0_7_0_1_1,
  input  [7:0] I0_7_0_1_2,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_0_0_1,
  input  [7:0] I1_0_0_2,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_1_0_1,
  input  [7:0] I1_1_0_2,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_2_0_1,
  input  [7:0] I1_2_0_2,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_3_0_1,
  input  [7:0] I1_3_0_2,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_4_0_1,
  input  [7:0] I1_4_0_2,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_5_0_1,
  input  [7:0] I1_5_0_2,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_6_0_1,
  input  [7:0] I1_6_0_2,
  input  [7:0] I1_7_0_0,
  input  [7:0] I1_7_0_1,
  input  [7:0] I1_7_0_2,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_0_0_1_0,
  output [7:0] O_0_0_1_1,
  output [7:0] O_0_0_1_2,
  output [7:0] O_0_0_2_0,
  output [7:0] O_0_0_2_1,
  output [7:0] O_0_0_2_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_1_0_1_0,
  output [7:0] O_1_0_1_1,
  output [7:0] O_1_0_1_2,
  output [7:0] O_1_0_2_0,
  output [7:0] O_1_0_2_1,
  output [7:0] O_1_0_2_2,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_0_2,
  output [7:0] O_2_0_1_0,
  output [7:0] O_2_0_1_1,
  output [7:0] O_2_0_1_2,
  output [7:0] O_2_0_2_0,
  output [7:0] O_2_0_2_1,
  output [7:0] O_2_0_2_2,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_0_2,
  output [7:0] O_3_0_1_0,
  output [7:0] O_3_0_1_1,
  output [7:0] O_3_0_1_2,
  output [7:0] O_3_0_2_0,
  output [7:0] O_3_0_2_1,
  output [7:0] O_3_0_2_2,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_0_2,
  output [7:0] O_4_0_1_0,
  output [7:0] O_4_0_1_1,
  output [7:0] O_4_0_1_2,
  output [7:0] O_4_0_2_0,
  output [7:0] O_4_0_2_1,
  output [7:0] O_4_0_2_2,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_0_2,
  output [7:0] O_5_0_1_0,
  output [7:0] O_5_0_1_1,
  output [7:0] O_5_0_1_2,
  output [7:0] O_5_0_2_0,
  output [7:0] O_5_0_2_1,
  output [7:0] O_5_0_2_2,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_0_2,
  output [7:0] O_6_0_1_0,
  output [7:0] O_6_0_1_1,
  output [7:0] O_6_0_1_2,
  output [7:0] O_6_0_2_0,
  output [7:0] O_6_0_2_1,
  output [7:0] O_6_0_2_2,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_0_2,
  output [7:0] O_7_0_1_0,
  output [7:0] O_7_0_1_1,
  output [7:0] O_7_0_1_2,
  output [7:0] O_7_0_2_0,
  output [7:0] O_7_0_2_1,
  output [7:0] O_7_0_2_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_2_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  Map2S_20 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0_0(fst_op_I0_0_0_0),
    .I0_0_0_1(fst_op_I0_0_0_1),
    .I0_0_0_2(fst_op_I0_0_0_2),
    .I0_0_1_0(fst_op_I0_0_1_0),
    .I0_0_1_1(fst_op_I0_0_1_1),
    .I0_0_1_2(fst_op_I0_0_1_2),
    .I1_0_0(fst_op_I1_0_0),
    .I1_0_1(fst_op_I1_0_1),
    .I1_0_2(fst_op_I1_0_2),
    .O_0_0_0(fst_op_O_0_0_0),
    .O_0_0_1(fst_op_O_0_0_1),
    .O_0_0_2(fst_op_O_0_0_2),
    .O_0_1_0(fst_op_O_0_1_0),
    .O_0_1_1(fst_op_O_0_1_1),
    .O_0_1_2(fst_op_O_0_1_2),
    .O_0_2_0(fst_op_O_0_2_0),
    .O_0_2_1(fst_op_O_0_2_1),
    .O_0_2_2(fst_op_O_0_2_2)
  );
  Map2S_20 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0_0(other_ops_0_I0_0_0_0),
    .I0_0_0_1(other_ops_0_I0_0_0_1),
    .I0_0_0_2(other_ops_0_I0_0_0_2),
    .I0_0_1_0(other_ops_0_I0_0_1_0),
    .I0_0_1_1(other_ops_0_I0_0_1_1),
    .I0_0_1_2(other_ops_0_I0_0_1_2),
    .I1_0_0(other_ops_0_I1_0_0),
    .I1_0_1(other_ops_0_I1_0_1),
    .I1_0_2(other_ops_0_I1_0_2),
    .O_0_0_0(other_ops_0_O_0_0_0),
    .O_0_0_1(other_ops_0_O_0_0_1),
    .O_0_0_2(other_ops_0_O_0_0_2),
    .O_0_1_0(other_ops_0_O_0_1_0),
    .O_0_1_1(other_ops_0_O_0_1_1),
    .O_0_1_2(other_ops_0_O_0_1_2),
    .O_0_2_0(other_ops_0_O_0_2_0),
    .O_0_2_1(other_ops_0_O_0_2_1),
    .O_0_2_2(other_ops_0_O_0_2_2)
  );
  Map2S_20 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0_0(other_ops_1_I0_0_0_0),
    .I0_0_0_1(other_ops_1_I0_0_0_1),
    .I0_0_0_2(other_ops_1_I0_0_0_2),
    .I0_0_1_0(other_ops_1_I0_0_1_0),
    .I0_0_1_1(other_ops_1_I0_0_1_1),
    .I0_0_1_2(other_ops_1_I0_0_1_2),
    .I1_0_0(other_ops_1_I1_0_0),
    .I1_0_1(other_ops_1_I1_0_1),
    .I1_0_2(other_ops_1_I1_0_2),
    .O_0_0_0(other_ops_1_O_0_0_0),
    .O_0_0_1(other_ops_1_O_0_0_1),
    .O_0_0_2(other_ops_1_O_0_0_2),
    .O_0_1_0(other_ops_1_O_0_1_0),
    .O_0_1_1(other_ops_1_O_0_1_1),
    .O_0_1_2(other_ops_1_O_0_1_2),
    .O_0_2_0(other_ops_1_O_0_2_0),
    .O_0_2_1(other_ops_1_O_0_2_1),
    .O_0_2_2(other_ops_1_O_0_2_2)
  );
  Map2S_20 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0_0(other_ops_2_I0_0_0_0),
    .I0_0_0_1(other_ops_2_I0_0_0_1),
    .I0_0_0_2(other_ops_2_I0_0_0_2),
    .I0_0_1_0(other_ops_2_I0_0_1_0),
    .I0_0_1_1(other_ops_2_I0_0_1_1),
    .I0_0_1_2(other_ops_2_I0_0_1_2),
    .I1_0_0(other_ops_2_I1_0_0),
    .I1_0_1(other_ops_2_I1_0_1),
    .I1_0_2(other_ops_2_I1_0_2),
    .O_0_0_0(other_ops_2_O_0_0_0),
    .O_0_0_1(other_ops_2_O_0_0_1),
    .O_0_0_2(other_ops_2_O_0_0_2),
    .O_0_1_0(other_ops_2_O_0_1_0),
    .O_0_1_1(other_ops_2_O_0_1_1),
    .O_0_1_2(other_ops_2_O_0_1_2),
    .O_0_2_0(other_ops_2_O_0_2_0),
    .O_0_2_1(other_ops_2_O_0_2_1),
    .O_0_2_2(other_ops_2_O_0_2_2)
  );
  Map2S_20 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0_0(other_ops_3_I0_0_0_0),
    .I0_0_0_1(other_ops_3_I0_0_0_1),
    .I0_0_0_2(other_ops_3_I0_0_0_2),
    .I0_0_1_0(other_ops_3_I0_0_1_0),
    .I0_0_1_1(other_ops_3_I0_0_1_1),
    .I0_0_1_2(other_ops_3_I0_0_1_2),
    .I1_0_0(other_ops_3_I1_0_0),
    .I1_0_1(other_ops_3_I1_0_1),
    .I1_0_2(other_ops_3_I1_0_2),
    .O_0_0_0(other_ops_3_O_0_0_0),
    .O_0_0_1(other_ops_3_O_0_0_1),
    .O_0_0_2(other_ops_3_O_0_0_2),
    .O_0_1_0(other_ops_3_O_0_1_0),
    .O_0_1_1(other_ops_3_O_0_1_1),
    .O_0_1_2(other_ops_3_O_0_1_2),
    .O_0_2_0(other_ops_3_O_0_2_0),
    .O_0_2_1(other_ops_3_O_0_2_1),
    .O_0_2_2(other_ops_3_O_0_2_2)
  );
  Map2S_20 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0_0(other_ops_4_I0_0_0_0),
    .I0_0_0_1(other_ops_4_I0_0_0_1),
    .I0_0_0_2(other_ops_4_I0_0_0_2),
    .I0_0_1_0(other_ops_4_I0_0_1_0),
    .I0_0_1_1(other_ops_4_I0_0_1_1),
    .I0_0_1_2(other_ops_4_I0_0_1_2),
    .I1_0_0(other_ops_4_I1_0_0),
    .I1_0_1(other_ops_4_I1_0_1),
    .I1_0_2(other_ops_4_I1_0_2),
    .O_0_0_0(other_ops_4_O_0_0_0),
    .O_0_0_1(other_ops_4_O_0_0_1),
    .O_0_0_2(other_ops_4_O_0_0_2),
    .O_0_1_0(other_ops_4_O_0_1_0),
    .O_0_1_1(other_ops_4_O_0_1_1),
    .O_0_1_2(other_ops_4_O_0_1_2),
    .O_0_2_0(other_ops_4_O_0_2_0),
    .O_0_2_1(other_ops_4_O_0_2_1),
    .O_0_2_2(other_ops_4_O_0_2_2)
  );
  Map2S_20 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0_0(other_ops_5_I0_0_0_0),
    .I0_0_0_1(other_ops_5_I0_0_0_1),
    .I0_0_0_2(other_ops_5_I0_0_0_2),
    .I0_0_1_0(other_ops_5_I0_0_1_0),
    .I0_0_1_1(other_ops_5_I0_0_1_1),
    .I0_0_1_2(other_ops_5_I0_0_1_2),
    .I1_0_0(other_ops_5_I1_0_0),
    .I1_0_1(other_ops_5_I1_0_1),
    .I1_0_2(other_ops_5_I1_0_2),
    .O_0_0_0(other_ops_5_O_0_0_0),
    .O_0_0_1(other_ops_5_O_0_0_1),
    .O_0_0_2(other_ops_5_O_0_0_2),
    .O_0_1_0(other_ops_5_O_0_1_0),
    .O_0_1_1(other_ops_5_O_0_1_1),
    .O_0_1_2(other_ops_5_O_0_1_2),
    .O_0_2_0(other_ops_5_O_0_2_0),
    .O_0_2_1(other_ops_5_O_0_2_1),
    .O_0_2_2(other_ops_5_O_0_2_2)
  );
  Map2S_20 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0_0(other_ops_6_I0_0_0_0),
    .I0_0_0_1(other_ops_6_I0_0_0_1),
    .I0_0_0_2(other_ops_6_I0_0_0_2),
    .I0_0_1_0(other_ops_6_I0_0_1_0),
    .I0_0_1_1(other_ops_6_I0_0_1_1),
    .I0_0_1_2(other_ops_6_I0_0_1_2),
    .I1_0_0(other_ops_6_I1_0_0),
    .I1_0_1(other_ops_6_I1_0_1),
    .I1_0_2(other_ops_6_I1_0_2),
    .O_0_0_0(other_ops_6_O_0_0_0),
    .O_0_0_1(other_ops_6_O_0_0_1),
    .O_0_0_2(other_ops_6_O_0_0_2),
    .O_0_1_0(other_ops_6_O_0_1_0),
    .O_0_1_1(other_ops_6_O_0_1_1),
    .O_0_1_2(other_ops_6_O_0_1_2),
    .O_0_2_0(other_ops_6_O_0_2_0),
    .O_0_2_1(other_ops_6_O_0_2_1),
    .O_0_2_2(other_ops_6_O_0_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0_0 = fst_op_O_0_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_0_1 = fst_op_O_0_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_0_2 = fst_op_O_0_0_2; // @[Map2S.scala 19:8]
  assign O_0_0_1_0 = fst_op_O_0_1_0; // @[Map2S.scala 19:8]
  assign O_0_0_1_1 = fst_op_O_0_1_1; // @[Map2S.scala 19:8]
  assign O_0_0_1_2 = fst_op_O_0_1_2; // @[Map2S.scala 19:8]
  assign O_0_0_2_0 = fst_op_O_0_2_0; // @[Map2S.scala 19:8]
  assign O_0_0_2_1 = fst_op_O_0_2_1; // @[Map2S.scala 19:8]
  assign O_0_0_2_2 = fst_op_O_0_2_2; // @[Map2S.scala 19:8]
  assign O_1_0_0_0 = other_ops_0_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_0_1 = other_ops_0_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_0_2 = other_ops_0_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_1_0_1_0 = other_ops_0_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_1_0_1_1 = other_ops_0_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_1_0_1_2 = other_ops_0_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_1_0_2_0 = other_ops_0_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_1_0_2_1 = other_ops_0_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_1_0_2_2 = other_ops_0_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_2_0_0_0 = other_ops_1_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_0_1 = other_ops_1_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_0_2 = other_ops_1_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_2_0_1_0 = other_ops_1_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_2_0_1_1 = other_ops_1_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_2_0_1_2 = other_ops_1_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_2_0_2_0 = other_ops_1_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_2_0_2_1 = other_ops_1_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_2_0_2_2 = other_ops_1_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_3_0_0_0 = other_ops_2_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_0_1 = other_ops_2_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_0_2 = other_ops_2_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_3_0_1_0 = other_ops_2_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_3_0_1_1 = other_ops_2_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_3_0_1_2 = other_ops_2_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_3_0_2_0 = other_ops_2_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_3_0_2_1 = other_ops_2_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_3_0_2_2 = other_ops_2_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_4_0_0_0 = other_ops_3_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_0_1 = other_ops_3_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_0_2 = other_ops_3_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_4_0_1_0 = other_ops_3_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_4_0_1_1 = other_ops_3_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_4_0_1_2 = other_ops_3_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_4_0_2_0 = other_ops_3_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_4_0_2_1 = other_ops_3_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_4_0_2_2 = other_ops_3_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_5_0_0_0 = other_ops_4_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_0_1 = other_ops_4_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_0_2 = other_ops_4_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_5_0_1_0 = other_ops_4_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_5_0_1_1 = other_ops_4_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_5_0_1_2 = other_ops_4_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_5_0_2_0 = other_ops_4_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_5_0_2_1 = other_ops_4_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_5_0_2_2 = other_ops_4_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_6_0_0_0 = other_ops_5_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_0_1 = other_ops_5_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_0_2 = other_ops_5_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_6_0_1_0 = other_ops_5_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_6_0_1_1 = other_ops_5_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_6_0_1_2 = other_ops_5_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_6_0_2_0 = other_ops_5_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_6_0_2_1 = other_ops_5_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_6_0_2_2 = other_ops_5_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_7_0_0_0 = other_ops_6_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_0_1 = other_ops_6_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_0_2 = other_ops_6_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_7_0_1_0 = other_ops_6_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_7_0_1_1 = other_ops_6_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_7_0_1_2 = other_ops_6_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_7_0_2_0 = other_ops_6_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_7_0_2_1 = other_ops_6_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_7_0_2_2 = other_ops_6_O_0_2_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0_0 = I0_0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_0_1 = I0_0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_0_2 = I0_0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1_0 = I0_0_0_1_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1_1 = I0_0_0_1_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1_2 = I0_0_0_1_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_0 = I1_0_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_1 = I1_0_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_2 = I1_0_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0_0 = I0_1_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_0_1 = I0_1_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_0_2 = I0_1_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1_0 = I0_1_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1_1 = I0_1_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1_2 = I0_1_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0_0 = I1_1_0_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_0_1 = I1_1_0_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_0_2 = I1_1_0_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0_0 = I0_2_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_0_1 = I0_2_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_0_2 = I0_2_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1_0 = I0_2_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1_1 = I0_2_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1_2 = I0_2_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0_0 = I1_2_0_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_0_1 = I1_2_0_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_0_2 = I1_2_0_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0_0 = I0_3_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_0_1 = I0_3_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_0_2 = I0_3_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1_0 = I0_3_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1_1 = I0_3_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1_2 = I0_3_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0_0 = I1_3_0_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_0_1 = I1_3_0_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_0_2 = I1_3_0_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0_0 = I0_4_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_0_1 = I0_4_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_0_2 = I0_4_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1_0 = I0_4_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1_1 = I0_4_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1_2 = I0_4_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0_0 = I1_4_0_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_0_1 = I1_4_0_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_0_2 = I1_4_0_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0_0 = I0_5_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_0_1 = I0_5_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_0_2 = I0_5_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1_0 = I0_5_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1_1 = I0_5_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1_2 = I0_5_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0_0 = I1_5_0_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_0_1 = I1_5_0_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_0_2 = I1_5_0_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0_0 = I0_6_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_0_1 = I0_6_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_0_2 = I0_6_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1_0 = I0_6_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1_1 = I0_6_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1_2 = I0_6_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0_0 = I1_6_0_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_0_1 = I1_6_0_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_0_2 = I1_6_0_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0_0 = I0_7_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_0_1 = I0_7_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_0_2 = I0_7_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1_0 = I0_7_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1_1 = I0_7_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1_2 = I0_7_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0_0 = I1_7_0_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_0_1 = I1_7_0_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_0_2 = I1_7_0_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_7(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0_0,
  input  [7:0] I0_0_0_0_1,
  input  [7:0] I0_0_0_0_2,
  input  [7:0] I0_0_0_1_0,
  input  [7:0] I0_0_0_1_1,
  input  [7:0] I0_0_0_1_2,
  input  [7:0] I0_1_0_0_0,
  input  [7:0] I0_1_0_0_1,
  input  [7:0] I0_1_0_0_2,
  input  [7:0] I0_1_0_1_0,
  input  [7:0] I0_1_0_1_1,
  input  [7:0] I0_1_0_1_2,
  input  [7:0] I0_2_0_0_0,
  input  [7:0] I0_2_0_0_1,
  input  [7:0] I0_2_0_0_2,
  input  [7:0] I0_2_0_1_0,
  input  [7:0] I0_2_0_1_1,
  input  [7:0] I0_2_0_1_2,
  input  [7:0] I0_3_0_0_0,
  input  [7:0] I0_3_0_0_1,
  input  [7:0] I0_3_0_0_2,
  input  [7:0] I0_3_0_1_0,
  input  [7:0] I0_3_0_1_1,
  input  [7:0] I0_3_0_1_2,
  input  [7:0] I0_4_0_0_0,
  input  [7:0] I0_4_0_0_1,
  input  [7:0] I0_4_0_0_2,
  input  [7:0] I0_4_0_1_0,
  input  [7:0] I0_4_0_1_1,
  input  [7:0] I0_4_0_1_2,
  input  [7:0] I0_5_0_0_0,
  input  [7:0] I0_5_0_0_1,
  input  [7:0] I0_5_0_0_2,
  input  [7:0] I0_5_0_1_0,
  input  [7:0] I0_5_0_1_1,
  input  [7:0] I0_5_0_1_2,
  input  [7:0] I0_6_0_0_0,
  input  [7:0] I0_6_0_0_1,
  input  [7:0] I0_6_0_0_2,
  input  [7:0] I0_6_0_1_0,
  input  [7:0] I0_6_0_1_1,
  input  [7:0] I0_6_0_1_2,
  input  [7:0] I0_7_0_0_0,
  input  [7:0] I0_7_0_0_1,
  input  [7:0] I0_7_0_0_2,
  input  [7:0] I0_7_0_1_0,
  input  [7:0] I0_7_0_1_1,
  input  [7:0] I0_7_0_1_2,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_0_0_1,
  input  [7:0] I1_0_0_2,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_1_0_1,
  input  [7:0] I1_1_0_2,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_2_0_1,
  input  [7:0] I1_2_0_2,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_3_0_1,
  input  [7:0] I1_3_0_2,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_4_0_1,
  input  [7:0] I1_4_0_2,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_5_0_1,
  input  [7:0] I1_5_0_2,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_6_0_1,
  input  [7:0] I1_6_0_2,
  input  [7:0] I1_7_0_0,
  input  [7:0] I1_7_0_1,
  input  [7:0] I1_7_0_2,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_0_0_1_0,
  output [7:0] O_0_0_1_1,
  output [7:0] O_0_0_1_2,
  output [7:0] O_0_0_2_0,
  output [7:0] O_0_0_2_1,
  output [7:0] O_0_0_2_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_1_0_1_0,
  output [7:0] O_1_0_1_1,
  output [7:0] O_1_0_1_2,
  output [7:0] O_1_0_2_0,
  output [7:0] O_1_0_2_1,
  output [7:0] O_1_0_2_2,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_0_2,
  output [7:0] O_2_0_1_0,
  output [7:0] O_2_0_1_1,
  output [7:0] O_2_0_1_2,
  output [7:0] O_2_0_2_0,
  output [7:0] O_2_0_2_1,
  output [7:0] O_2_0_2_2,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_0_2,
  output [7:0] O_3_0_1_0,
  output [7:0] O_3_0_1_1,
  output [7:0] O_3_0_1_2,
  output [7:0] O_3_0_2_0,
  output [7:0] O_3_0_2_1,
  output [7:0] O_3_0_2_2,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_0_2,
  output [7:0] O_4_0_1_0,
  output [7:0] O_4_0_1_1,
  output [7:0] O_4_0_1_2,
  output [7:0] O_4_0_2_0,
  output [7:0] O_4_0_2_1,
  output [7:0] O_4_0_2_2,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_0_2,
  output [7:0] O_5_0_1_0,
  output [7:0] O_5_0_1_1,
  output [7:0] O_5_0_1_2,
  output [7:0] O_5_0_2_0,
  output [7:0] O_5_0_2_1,
  output [7:0] O_5_0_2_2,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_0_2,
  output [7:0] O_6_0_1_0,
  output [7:0] O_6_0_1_1,
  output [7:0] O_6_0_1_2,
  output [7:0] O_6_0_2_0,
  output [7:0] O_6_0_2_1,
  output [7:0] O_6_0_2_2,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_0_2,
  output [7:0] O_7_0_1_0,
  output [7:0] O_7_0_1_1,
  output [7:0] O_7_0_1_2,
  output [7:0] O_7_0_2_0,
  output [7:0] O_7_0_2_1,
  output [7:0] O_7_0_2_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_2_2; // @[Map2T.scala 8:20]
  Map2S_21 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0_0(op_I0_0_0_0_0),
    .I0_0_0_0_1(op_I0_0_0_0_1),
    .I0_0_0_0_2(op_I0_0_0_0_2),
    .I0_0_0_1_0(op_I0_0_0_1_0),
    .I0_0_0_1_1(op_I0_0_0_1_1),
    .I0_0_0_1_2(op_I0_0_0_1_2),
    .I0_1_0_0_0(op_I0_1_0_0_0),
    .I0_1_0_0_1(op_I0_1_0_0_1),
    .I0_1_0_0_2(op_I0_1_0_0_2),
    .I0_1_0_1_0(op_I0_1_0_1_0),
    .I0_1_0_1_1(op_I0_1_0_1_1),
    .I0_1_0_1_2(op_I0_1_0_1_2),
    .I0_2_0_0_0(op_I0_2_0_0_0),
    .I0_2_0_0_1(op_I0_2_0_0_1),
    .I0_2_0_0_2(op_I0_2_0_0_2),
    .I0_2_0_1_0(op_I0_2_0_1_0),
    .I0_2_0_1_1(op_I0_2_0_1_1),
    .I0_2_0_1_2(op_I0_2_0_1_2),
    .I0_3_0_0_0(op_I0_3_0_0_0),
    .I0_3_0_0_1(op_I0_3_0_0_1),
    .I0_3_0_0_2(op_I0_3_0_0_2),
    .I0_3_0_1_0(op_I0_3_0_1_0),
    .I0_3_0_1_1(op_I0_3_0_1_1),
    .I0_3_0_1_2(op_I0_3_0_1_2),
    .I0_4_0_0_0(op_I0_4_0_0_0),
    .I0_4_0_0_1(op_I0_4_0_0_1),
    .I0_4_0_0_2(op_I0_4_0_0_2),
    .I0_4_0_1_0(op_I0_4_0_1_0),
    .I0_4_0_1_1(op_I0_4_0_1_1),
    .I0_4_0_1_2(op_I0_4_0_1_2),
    .I0_5_0_0_0(op_I0_5_0_0_0),
    .I0_5_0_0_1(op_I0_5_0_0_1),
    .I0_5_0_0_2(op_I0_5_0_0_2),
    .I0_5_0_1_0(op_I0_5_0_1_0),
    .I0_5_0_1_1(op_I0_5_0_1_1),
    .I0_5_0_1_2(op_I0_5_0_1_2),
    .I0_6_0_0_0(op_I0_6_0_0_0),
    .I0_6_0_0_1(op_I0_6_0_0_1),
    .I0_6_0_0_2(op_I0_6_0_0_2),
    .I0_6_0_1_0(op_I0_6_0_1_0),
    .I0_6_0_1_1(op_I0_6_0_1_1),
    .I0_6_0_1_2(op_I0_6_0_1_2),
    .I0_7_0_0_0(op_I0_7_0_0_0),
    .I0_7_0_0_1(op_I0_7_0_0_1),
    .I0_7_0_0_2(op_I0_7_0_0_2),
    .I0_7_0_1_0(op_I0_7_0_1_0),
    .I0_7_0_1_1(op_I0_7_0_1_1),
    .I0_7_0_1_2(op_I0_7_0_1_2),
    .I1_0_0_0(op_I1_0_0_0),
    .I1_0_0_1(op_I1_0_0_1),
    .I1_0_0_2(op_I1_0_0_2),
    .I1_1_0_0(op_I1_1_0_0),
    .I1_1_0_1(op_I1_1_0_1),
    .I1_1_0_2(op_I1_1_0_2),
    .I1_2_0_0(op_I1_2_0_0),
    .I1_2_0_1(op_I1_2_0_1),
    .I1_2_0_2(op_I1_2_0_2),
    .I1_3_0_0(op_I1_3_0_0),
    .I1_3_0_1(op_I1_3_0_1),
    .I1_3_0_2(op_I1_3_0_2),
    .I1_4_0_0(op_I1_4_0_0),
    .I1_4_0_1(op_I1_4_0_1),
    .I1_4_0_2(op_I1_4_0_2),
    .I1_5_0_0(op_I1_5_0_0),
    .I1_5_0_1(op_I1_5_0_1),
    .I1_5_0_2(op_I1_5_0_2),
    .I1_6_0_0(op_I1_6_0_0),
    .I1_6_0_1(op_I1_6_0_1),
    .I1_6_0_2(op_I1_6_0_2),
    .I1_7_0_0(op_I1_7_0_0),
    .I1_7_0_1(op_I1_7_0_1),
    .I1_7_0_2(op_I1_7_0_2),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_0_0_0_2(op_O_0_0_0_2),
    .O_0_0_1_0(op_O_0_0_1_0),
    .O_0_0_1_1(op_O_0_0_1_1),
    .O_0_0_1_2(op_O_0_0_1_2),
    .O_0_0_2_0(op_O_0_0_2_0),
    .O_0_0_2_1(op_O_0_0_2_1),
    .O_0_0_2_2(op_O_0_0_2_2),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_1_0_0_2(op_O_1_0_0_2),
    .O_1_0_1_0(op_O_1_0_1_0),
    .O_1_0_1_1(op_O_1_0_1_1),
    .O_1_0_1_2(op_O_1_0_1_2),
    .O_1_0_2_0(op_O_1_0_2_0),
    .O_1_0_2_1(op_O_1_0_2_1),
    .O_1_0_2_2(op_O_1_0_2_2),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_2_0_0_2(op_O_2_0_0_2),
    .O_2_0_1_0(op_O_2_0_1_0),
    .O_2_0_1_1(op_O_2_0_1_1),
    .O_2_0_1_2(op_O_2_0_1_2),
    .O_2_0_2_0(op_O_2_0_2_0),
    .O_2_0_2_1(op_O_2_0_2_1),
    .O_2_0_2_2(op_O_2_0_2_2),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_3_0_0_2(op_O_3_0_0_2),
    .O_3_0_1_0(op_O_3_0_1_0),
    .O_3_0_1_1(op_O_3_0_1_1),
    .O_3_0_1_2(op_O_3_0_1_2),
    .O_3_0_2_0(op_O_3_0_2_0),
    .O_3_0_2_1(op_O_3_0_2_1),
    .O_3_0_2_2(op_O_3_0_2_2),
    .O_4_0_0_0(op_O_4_0_0_0),
    .O_4_0_0_1(op_O_4_0_0_1),
    .O_4_0_0_2(op_O_4_0_0_2),
    .O_4_0_1_0(op_O_4_0_1_0),
    .O_4_0_1_1(op_O_4_0_1_1),
    .O_4_0_1_2(op_O_4_0_1_2),
    .O_4_0_2_0(op_O_4_0_2_0),
    .O_4_0_2_1(op_O_4_0_2_1),
    .O_4_0_2_2(op_O_4_0_2_2),
    .O_5_0_0_0(op_O_5_0_0_0),
    .O_5_0_0_1(op_O_5_0_0_1),
    .O_5_0_0_2(op_O_5_0_0_2),
    .O_5_0_1_0(op_O_5_0_1_0),
    .O_5_0_1_1(op_O_5_0_1_1),
    .O_5_0_1_2(op_O_5_0_1_2),
    .O_5_0_2_0(op_O_5_0_2_0),
    .O_5_0_2_1(op_O_5_0_2_1),
    .O_5_0_2_2(op_O_5_0_2_2),
    .O_6_0_0_0(op_O_6_0_0_0),
    .O_6_0_0_1(op_O_6_0_0_1),
    .O_6_0_0_2(op_O_6_0_0_2),
    .O_6_0_1_0(op_O_6_0_1_0),
    .O_6_0_1_1(op_O_6_0_1_1),
    .O_6_0_1_2(op_O_6_0_1_2),
    .O_6_0_2_0(op_O_6_0_2_0),
    .O_6_0_2_1(op_O_6_0_2_1),
    .O_6_0_2_2(op_O_6_0_2_2),
    .O_7_0_0_0(op_O_7_0_0_0),
    .O_7_0_0_1(op_O_7_0_0_1),
    .O_7_0_0_2(op_O_7_0_0_2),
    .O_7_0_1_0(op_O_7_0_1_0),
    .O_7_0_1_1(op_O_7_0_1_1),
    .O_7_0_1_2(op_O_7_0_1_2),
    .O_7_0_2_0(op_O_7_0_2_0),
    .O_7_0_2_1(op_O_7_0_2_1),
    .O_7_0_2_2(op_O_7_0_2_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_0_2 = op_O_0_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_0_1_0 = op_O_0_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_0_1_1 = op_O_0_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_0_1_2 = op_O_0_0_1_2; // @[Map2T.scala 17:7]
  assign O_0_0_2_0 = op_O_0_0_2_0; // @[Map2T.scala 17:7]
  assign O_0_0_2_1 = op_O_0_0_2_1; // @[Map2T.scala 17:7]
  assign O_0_0_2_2 = op_O_0_0_2_2; // @[Map2T.scala 17:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_0_2 = op_O_1_0_0_2; // @[Map2T.scala 17:7]
  assign O_1_0_1_0 = op_O_1_0_1_0; // @[Map2T.scala 17:7]
  assign O_1_0_1_1 = op_O_1_0_1_1; // @[Map2T.scala 17:7]
  assign O_1_0_1_2 = op_O_1_0_1_2; // @[Map2T.scala 17:7]
  assign O_1_0_2_0 = op_O_1_0_2_0; // @[Map2T.scala 17:7]
  assign O_1_0_2_1 = op_O_1_0_2_1; // @[Map2T.scala 17:7]
  assign O_1_0_2_2 = op_O_1_0_2_2; // @[Map2T.scala 17:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_0_2 = op_O_2_0_0_2; // @[Map2T.scala 17:7]
  assign O_2_0_1_0 = op_O_2_0_1_0; // @[Map2T.scala 17:7]
  assign O_2_0_1_1 = op_O_2_0_1_1; // @[Map2T.scala 17:7]
  assign O_2_0_1_2 = op_O_2_0_1_2; // @[Map2T.scala 17:7]
  assign O_2_0_2_0 = op_O_2_0_2_0; // @[Map2T.scala 17:7]
  assign O_2_0_2_1 = op_O_2_0_2_1; // @[Map2T.scala 17:7]
  assign O_2_0_2_2 = op_O_2_0_2_2; // @[Map2T.scala 17:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_0_2 = op_O_3_0_0_2; // @[Map2T.scala 17:7]
  assign O_3_0_1_0 = op_O_3_0_1_0; // @[Map2T.scala 17:7]
  assign O_3_0_1_1 = op_O_3_0_1_1; // @[Map2T.scala 17:7]
  assign O_3_0_1_2 = op_O_3_0_1_2; // @[Map2T.scala 17:7]
  assign O_3_0_2_0 = op_O_3_0_2_0; // @[Map2T.scala 17:7]
  assign O_3_0_2_1 = op_O_3_0_2_1; // @[Map2T.scala 17:7]
  assign O_3_0_2_2 = op_O_3_0_2_2; // @[Map2T.scala 17:7]
  assign O_4_0_0_0 = op_O_4_0_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_0_1 = op_O_4_0_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_0_2 = op_O_4_0_0_2; // @[Map2T.scala 17:7]
  assign O_4_0_1_0 = op_O_4_0_1_0; // @[Map2T.scala 17:7]
  assign O_4_0_1_1 = op_O_4_0_1_1; // @[Map2T.scala 17:7]
  assign O_4_0_1_2 = op_O_4_0_1_2; // @[Map2T.scala 17:7]
  assign O_4_0_2_0 = op_O_4_0_2_0; // @[Map2T.scala 17:7]
  assign O_4_0_2_1 = op_O_4_0_2_1; // @[Map2T.scala 17:7]
  assign O_4_0_2_2 = op_O_4_0_2_2; // @[Map2T.scala 17:7]
  assign O_5_0_0_0 = op_O_5_0_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_0_1 = op_O_5_0_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_0_2 = op_O_5_0_0_2; // @[Map2T.scala 17:7]
  assign O_5_0_1_0 = op_O_5_0_1_0; // @[Map2T.scala 17:7]
  assign O_5_0_1_1 = op_O_5_0_1_1; // @[Map2T.scala 17:7]
  assign O_5_0_1_2 = op_O_5_0_1_2; // @[Map2T.scala 17:7]
  assign O_5_0_2_0 = op_O_5_0_2_0; // @[Map2T.scala 17:7]
  assign O_5_0_2_1 = op_O_5_0_2_1; // @[Map2T.scala 17:7]
  assign O_5_0_2_2 = op_O_5_0_2_2; // @[Map2T.scala 17:7]
  assign O_6_0_0_0 = op_O_6_0_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_0_1 = op_O_6_0_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_0_2 = op_O_6_0_0_2; // @[Map2T.scala 17:7]
  assign O_6_0_1_0 = op_O_6_0_1_0; // @[Map2T.scala 17:7]
  assign O_6_0_1_1 = op_O_6_0_1_1; // @[Map2T.scala 17:7]
  assign O_6_0_1_2 = op_O_6_0_1_2; // @[Map2T.scala 17:7]
  assign O_6_0_2_0 = op_O_6_0_2_0; // @[Map2T.scala 17:7]
  assign O_6_0_2_1 = op_O_6_0_2_1; // @[Map2T.scala 17:7]
  assign O_6_0_2_2 = op_O_6_0_2_2; // @[Map2T.scala 17:7]
  assign O_7_0_0_0 = op_O_7_0_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_0_1 = op_O_7_0_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_0_2 = op_O_7_0_0_2; // @[Map2T.scala 17:7]
  assign O_7_0_1_0 = op_O_7_0_1_0; // @[Map2T.scala 17:7]
  assign O_7_0_1_1 = op_O_7_0_1_1; // @[Map2T.scala 17:7]
  assign O_7_0_1_2 = op_O_7_0_1_2; // @[Map2T.scala 17:7]
  assign O_7_0_2_0 = op_O_7_0_2_0; // @[Map2T.scala 17:7]
  assign O_7_0_2_1 = op_O_7_0_2_1; // @[Map2T.scala 17:7]
  assign O_7_0_2_2 = op_O_7_0_2_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0_0 = I0_0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_0_1 = I0_0_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_0_0_2 = I0_0_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1_0 = I0_0_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1_1 = I0_0_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1_2 = I0_0_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0_0 = I0_1_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0_1 = I0_1_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0_2 = I0_1_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1_0 = I0_1_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1_1 = I0_1_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1_2 = I0_1_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0_0 = I0_2_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0_1 = I0_2_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0_2 = I0_2_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1_0 = I0_2_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1_1 = I0_2_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1_2 = I0_2_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0_0 = I0_3_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0_1 = I0_3_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0_2 = I0_3_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1_0 = I0_3_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1_1 = I0_3_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1_2 = I0_3_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0_0 = I0_4_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0_1 = I0_4_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0_2 = I0_4_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0_1_0 = I0_4_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_1_1 = I0_4_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0_1_2 = I0_4_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0_0 = I0_5_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0_1 = I0_5_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0_2 = I0_5_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0_1_0 = I0_5_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_1_1 = I0_5_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0_1_2 = I0_5_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0_0 = I0_6_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0_1 = I0_6_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0_2 = I0_6_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0_1_0 = I0_6_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_1_1 = I0_6_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0_1_2 = I0_6_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0_0 = I0_7_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0_1 = I0_7_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0_2 = I0_7_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0_1_0 = I0_7_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_1_1 = I0_7_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0_1_2 = I0_7_0_1_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0_0 = I1_0_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_0_1 = I1_0_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_0_2 = I1_0_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0_0 = I1_1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_1_0_1 = I1_1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_1_0_2 = I1_1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0_0 = I1_2_0_0; // @[Map2T.scala 16:11]
  assign op_I1_2_0_1 = I1_2_0_1; // @[Map2T.scala 16:11]
  assign op_I1_2_0_2 = I1_2_0_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0_0 = I1_3_0_0; // @[Map2T.scala 16:11]
  assign op_I1_3_0_1 = I1_3_0_1; // @[Map2T.scala 16:11]
  assign op_I1_3_0_2 = I1_3_0_2; // @[Map2T.scala 16:11]
  assign op_I1_4_0_0 = I1_4_0_0; // @[Map2T.scala 16:11]
  assign op_I1_4_0_1 = I1_4_0_1; // @[Map2T.scala 16:11]
  assign op_I1_4_0_2 = I1_4_0_2; // @[Map2T.scala 16:11]
  assign op_I1_5_0_0 = I1_5_0_0; // @[Map2T.scala 16:11]
  assign op_I1_5_0_1 = I1_5_0_1; // @[Map2T.scala 16:11]
  assign op_I1_5_0_2 = I1_5_0_2; // @[Map2T.scala 16:11]
  assign op_I1_6_0_0 = I1_6_0_0; // @[Map2T.scala 16:11]
  assign op_I1_6_0_1 = I1_6_0_1; // @[Map2T.scala 16:11]
  assign op_I1_6_0_2 = I1_6_0_2; // @[Map2T.scala 16:11]
  assign op_I1_7_0_0 = I1_7_0_0; // @[Map2T.scala 16:11]
  assign op_I1_7_0_1 = I1_7_0_1; // @[Map2T.scala 16:11]
  assign op_I1_7_0_2 = I1_7_0_2; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleToSSeq_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0_0 = I_0_0; // @[Tuple.scala 41:5]
  assign O_0_1 = I_0_1; // @[Tuple.scala 41:5]
  assign O_0_2 = I_0_2; // @[Tuple.scala 41:5]
  assign O_1_0 = I_1_0; // @[Tuple.scala 41:5]
  assign O_1_1 = I_1_1; // @[Tuple.scala 41:5]
  assign O_1_2 = I_1_2; // @[Tuple.scala 41:5]
  assign O_2_0 = I_2_0; // @[Tuple.scala 41:5]
  assign O_2_1 = I_2_1; // @[Tuple.scala 41:5]
  assign O_2_2 = I_2_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_3 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0_0(op_inst_I_0_0),
    .I_0_1(op_inst_I_0_1),
    .I_0_2(op_inst_I_0_2),
    .I_1_0(op_inst_I_1_0),
    .I_1_1(op_inst_I_1_1),
    .I_1_2(op_inst_I_1_2),
    .I_2_0(op_inst_I_2_0),
    .I_2_1(op_inst_I_2_1),
    .I_2_2(op_inst_I_2_2),
    .O_0_0(op_inst_O_0_0),
    .O_0_1(op_inst_O_0_1),
    .O_0_2(op_inst_O_0_2),
    .O_1_0(op_inst_O_1_0),
    .O_1_1(op_inst_O_1_1),
    .O_1_2(op_inst_O_1_2),
    .O_2_0(op_inst_O_2_0),
    .O_2_1(op_inst_O_2_1),
    .O_2_2(op_inst_O_2_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0_0 = op_inst_O_0_0; // @[Remove1S.scala 14:5]
  assign O_0_1 = op_inst_O_0_1; // @[Remove1S.scala 14:5]
  assign O_0_2 = op_inst_O_0_2; // @[Remove1S.scala 14:5]
  assign O_1_0 = op_inst_O_1_0; // @[Remove1S.scala 14:5]
  assign O_1_1 = op_inst_O_1_1; // @[Remove1S.scala 14:5]
  assign O_1_2 = op_inst_O_1_2; // @[Remove1S.scala 14:5]
  assign O_2_0 = op_inst_O_2_0; // @[Remove1S.scala 14:5]
  assign O_2_1 = op_inst_O_2_1; // @[Remove1S.scala 14:5]
  assign O_2_2 = op_inst_O_2_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0_0 = I_0_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_1 = I_0_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_2 = I_0_0_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_0 = I_0_1_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_1 = I_0_1_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_2 = I_0_1_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_0 = I_0_2_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_1 = I_0_2_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_2 = I_0_2_2; // @[Remove1S.scala 13:13]
endmodule
module MapS_6(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0_0,
  input  [7:0] I_0_0_0_1,
  input  [7:0] I_0_0_0_2,
  input  [7:0] I_0_0_1_0,
  input  [7:0] I_0_0_1_1,
  input  [7:0] I_0_0_1_2,
  input  [7:0] I_0_0_2_0,
  input  [7:0] I_0_0_2_1,
  input  [7:0] I_0_0_2_2,
  input  [7:0] I_1_0_0_0,
  input  [7:0] I_1_0_0_1,
  input  [7:0] I_1_0_0_2,
  input  [7:0] I_1_0_1_0,
  input  [7:0] I_1_0_1_1,
  input  [7:0] I_1_0_1_2,
  input  [7:0] I_1_0_2_0,
  input  [7:0] I_1_0_2_1,
  input  [7:0] I_1_0_2_2,
  input  [7:0] I_2_0_0_0,
  input  [7:0] I_2_0_0_1,
  input  [7:0] I_2_0_0_2,
  input  [7:0] I_2_0_1_0,
  input  [7:0] I_2_0_1_1,
  input  [7:0] I_2_0_1_2,
  input  [7:0] I_2_0_2_0,
  input  [7:0] I_2_0_2_1,
  input  [7:0] I_2_0_2_2,
  input  [7:0] I_3_0_0_0,
  input  [7:0] I_3_0_0_1,
  input  [7:0] I_3_0_0_2,
  input  [7:0] I_3_0_1_0,
  input  [7:0] I_3_0_1_1,
  input  [7:0] I_3_0_1_2,
  input  [7:0] I_3_0_2_0,
  input  [7:0] I_3_0_2_1,
  input  [7:0] I_3_0_2_2,
  input  [7:0] I_4_0_0_0,
  input  [7:0] I_4_0_0_1,
  input  [7:0] I_4_0_0_2,
  input  [7:0] I_4_0_1_0,
  input  [7:0] I_4_0_1_1,
  input  [7:0] I_4_0_1_2,
  input  [7:0] I_4_0_2_0,
  input  [7:0] I_4_0_2_1,
  input  [7:0] I_4_0_2_2,
  input  [7:0] I_5_0_0_0,
  input  [7:0] I_5_0_0_1,
  input  [7:0] I_5_0_0_2,
  input  [7:0] I_5_0_1_0,
  input  [7:0] I_5_0_1_1,
  input  [7:0] I_5_0_1_2,
  input  [7:0] I_5_0_2_0,
  input  [7:0] I_5_0_2_1,
  input  [7:0] I_5_0_2_2,
  input  [7:0] I_6_0_0_0,
  input  [7:0] I_6_0_0_1,
  input  [7:0] I_6_0_0_2,
  input  [7:0] I_6_0_1_0,
  input  [7:0] I_6_0_1_1,
  input  [7:0] I_6_0_1_2,
  input  [7:0] I_6_0_2_0,
  input  [7:0] I_6_0_2_1,
  input  [7:0] I_6_0_2_2,
  input  [7:0] I_7_0_0_0,
  input  [7:0] I_7_0_0_1,
  input  [7:0] I_7_0_0_2,
  input  [7:0] I_7_0_1_0,
  input  [7:0] I_7_0_1_1,
  input  [7:0] I_7_0_1_2,
  input  [7:0] I_7_0_2_0,
  input  [7:0] I_7_0_2_1,
  input  [7:0] I_7_0_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_1_2_0,
  output [7:0] O_1_2_1,
  output [7:0] O_1_2_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_2_1_2,
  output [7:0] O_2_2_0,
  output [7:0] O_2_2_1,
  output [7:0] O_2_2_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_3_1_2,
  output [7:0] O_3_2_0,
  output [7:0] O_3_2_1,
  output [7:0] O_3_2_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_4_1_2,
  output [7:0] O_4_2_0,
  output [7:0] O_4_2_1,
  output [7:0] O_4_2_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_5_1_2,
  output [7:0] O_5_2_0,
  output [7:0] O_5_2_1,
  output [7:0] O_5_2_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_6_1_2,
  output [7:0] O_6_2_0,
  output [7:0] O_6_2_1,
  output [7:0] O_6_2_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_7_1_2,
  output [7:0] O_7_2_0,
  output [7:0] O_7_2_1,
  output [7:0] O_7_2_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_2_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  Remove1S_3 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0_0(fst_op_I_0_0_0),
    .I_0_0_1(fst_op_I_0_0_1),
    .I_0_0_2(fst_op_I_0_0_2),
    .I_0_1_0(fst_op_I_0_1_0),
    .I_0_1_1(fst_op_I_0_1_1),
    .I_0_1_2(fst_op_I_0_1_2),
    .I_0_2_0(fst_op_I_0_2_0),
    .I_0_2_1(fst_op_I_0_2_1),
    .I_0_2_2(fst_op_I_0_2_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  Remove1S_3 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0_0(other_ops_0_I_0_0_0),
    .I_0_0_1(other_ops_0_I_0_0_1),
    .I_0_0_2(other_ops_0_I_0_0_2),
    .I_0_1_0(other_ops_0_I_0_1_0),
    .I_0_1_1(other_ops_0_I_0_1_1),
    .I_0_1_2(other_ops_0_I_0_1_2),
    .I_0_2_0(other_ops_0_I_0_2_0),
    .I_0_2_1(other_ops_0_I_0_2_1),
    .I_0_2_2(other_ops_0_I_0_2_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  Remove1S_3 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0_0(other_ops_1_I_0_0_0),
    .I_0_0_1(other_ops_1_I_0_0_1),
    .I_0_0_2(other_ops_1_I_0_0_2),
    .I_0_1_0(other_ops_1_I_0_1_0),
    .I_0_1_1(other_ops_1_I_0_1_1),
    .I_0_1_2(other_ops_1_I_0_1_2),
    .I_0_2_0(other_ops_1_I_0_2_0),
    .I_0_2_1(other_ops_1_I_0_2_1),
    .I_0_2_2(other_ops_1_I_0_2_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  Remove1S_3 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0_0(other_ops_2_I_0_0_0),
    .I_0_0_1(other_ops_2_I_0_0_1),
    .I_0_0_2(other_ops_2_I_0_0_2),
    .I_0_1_0(other_ops_2_I_0_1_0),
    .I_0_1_1(other_ops_2_I_0_1_1),
    .I_0_1_2(other_ops_2_I_0_1_2),
    .I_0_2_0(other_ops_2_I_0_2_0),
    .I_0_2_1(other_ops_2_I_0_2_1),
    .I_0_2_2(other_ops_2_I_0_2_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  Remove1S_3 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0_0(other_ops_3_I_0_0_0),
    .I_0_0_1(other_ops_3_I_0_0_1),
    .I_0_0_2(other_ops_3_I_0_0_2),
    .I_0_1_0(other_ops_3_I_0_1_0),
    .I_0_1_1(other_ops_3_I_0_1_1),
    .I_0_1_2(other_ops_3_I_0_1_2),
    .I_0_2_0(other_ops_3_I_0_2_0),
    .I_0_2_1(other_ops_3_I_0_2_1),
    .I_0_2_2(other_ops_3_I_0_2_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2),
    .O_2_0(other_ops_3_O_2_0),
    .O_2_1(other_ops_3_O_2_1),
    .O_2_2(other_ops_3_O_2_2)
  );
  Remove1S_3 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0_0(other_ops_4_I_0_0_0),
    .I_0_0_1(other_ops_4_I_0_0_1),
    .I_0_0_2(other_ops_4_I_0_0_2),
    .I_0_1_0(other_ops_4_I_0_1_0),
    .I_0_1_1(other_ops_4_I_0_1_1),
    .I_0_1_2(other_ops_4_I_0_1_2),
    .I_0_2_0(other_ops_4_I_0_2_0),
    .I_0_2_1(other_ops_4_I_0_2_1),
    .I_0_2_2(other_ops_4_I_0_2_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2),
    .O_2_0(other_ops_4_O_2_0),
    .O_2_1(other_ops_4_O_2_1),
    .O_2_2(other_ops_4_O_2_2)
  );
  Remove1S_3 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0_0(other_ops_5_I_0_0_0),
    .I_0_0_1(other_ops_5_I_0_0_1),
    .I_0_0_2(other_ops_5_I_0_0_2),
    .I_0_1_0(other_ops_5_I_0_1_0),
    .I_0_1_1(other_ops_5_I_0_1_1),
    .I_0_1_2(other_ops_5_I_0_1_2),
    .I_0_2_0(other_ops_5_I_0_2_0),
    .I_0_2_1(other_ops_5_I_0_2_1),
    .I_0_2_2(other_ops_5_I_0_2_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2),
    .O_2_0(other_ops_5_O_2_0),
    .O_2_1(other_ops_5_O_2_1),
    .O_2_2(other_ops_5_O_2_2)
  );
  Remove1S_3 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0_0(other_ops_6_I_0_0_0),
    .I_0_0_1(other_ops_6_I_0_0_1),
    .I_0_0_2(other_ops_6_I_0_0_2),
    .I_0_1_0(other_ops_6_I_0_1_0),
    .I_0_1_1(other_ops_6_I_0_1_1),
    .I_0_1_2(other_ops_6_I_0_1_2),
    .I_0_2_0(other_ops_6_I_0_2_0),
    .I_0_2_1(other_ops_6_I_0_2_1),
    .I_0_2_2(other_ops_6_I_0_2_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2),
    .O_2_0(other_ops_6_O_2_0),
    .O_2_1(other_ops_6_O_2_1),
    .O_2_2(other_ops_6_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[MapS.scala 17:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[MapS.scala 17:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[MapS.scala 17:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[MapS.scala 17:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[MapS.scala 17:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[MapS.scala 17:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[MapS.scala 17:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[MapS.scala 21:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[MapS.scala 21:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[MapS.scala 21:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[MapS.scala 21:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[MapS.scala 21:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[MapS.scala 21:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[MapS.scala 21:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[MapS.scala 21:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[MapS.scala 21:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[MapS.scala 21:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[MapS.scala 21:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[MapS.scala 21:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[MapS.scala 21:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[MapS.scala 21:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[MapS.scala 21:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[MapS.scala 21:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[MapS.scala 21:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[MapS.scala 21:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[MapS.scala 21:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[MapS.scala 21:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[MapS.scala 21:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[MapS.scala 21:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[MapS.scala 21:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[MapS.scala 21:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[MapS.scala 21:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[MapS.scala 21:12]
  assign O_4_2_0 = other_ops_3_O_2_0; // @[MapS.scala 21:12]
  assign O_4_2_1 = other_ops_3_O_2_1; // @[MapS.scala 21:12]
  assign O_4_2_2 = other_ops_3_O_2_2; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[MapS.scala 21:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[MapS.scala 21:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[MapS.scala 21:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[MapS.scala 21:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[MapS.scala 21:12]
  assign O_5_2_0 = other_ops_4_O_2_0; // @[MapS.scala 21:12]
  assign O_5_2_1 = other_ops_4_O_2_1; // @[MapS.scala 21:12]
  assign O_5_2_2 = other_ops_4_O_2_2; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[MapS.scala 21:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[MapS.scala 21:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[MapS.scala 21:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[MapS.scala 21:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[MapS.scala 21:12]
  assign O_6_2_0 = other_ops_5_O_2_0; // @[MapS.scala 21:12]
  assign O_6_2_1 = other_ops_5_O_2_1; // @[MapS.scala 21:12]
  assign O_6_2_2 = other_ops_5_O_2_2; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[MapS.scala 21:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[MapS.scala 21:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[MapS.scala 21:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[MapS.scala 21:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[MapS.scala 21:12]
  assign O_7_2_0 = other_ops_6_O_2_0; // @[MapS.scala 21:12]
  assign O_7_2_1 = other_ops_6_O_2_1; // @[MapS.scala 21:12]
  assign O_7_2_2 = other_ops_6_O_2_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0_0 = I_0_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_1 = I_0_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_2 = I_0_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_0 = I_0_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_1 = I_0_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_2 = I_0_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_0 = I_0_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_1 = I_0_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_2 = I_0_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0_0 = I_1_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_1 = I_1_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_2 = I_1_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_0 = I_1_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_1 = I_1_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_2 = I_1_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_0 = I_1_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_1 = I_1_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_2 = I_1_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0_0 = I_2_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_1 = I_2_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_2 = I_2_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_0 = I_2_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_1 = I_2_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_2 = I_2_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_0 = I_2_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_1 = I_2_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_2 = I_2_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0_0 = I_3_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_1 = I_3_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_2 = I_3_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_0 = I_3_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_1 = I_3_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_2 = I_3_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_0 = I_3_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_1 = I_3_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_2 = I_3_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0_0 = I_4_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_1 = I_4_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_2 = I_4_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_0 = I_4_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_1 = I_4_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_2 = I_4_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_0 = I_4_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_1 = I_4_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_2 = I_4_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0_0 = I_5_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_1 = I_5_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_2 = I_5_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_0 = I_5_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_1 = I_5_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_2 = I_5_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_0 = I_5_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_1 = I_5_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_2 = I_5_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0_0 = I_6_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_1 = I_6_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_2 = I_6_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_0 = I_6_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_1 = I_6_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_2 = I_6_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_0 = I_6_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_1 = I_6_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_2 = I_6_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0_0 = I_7_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_1 = I_7_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_2 = I_7_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_0 = I_7_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_1 = I_7_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_2 = I_7_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_0 = I_7_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_1 = I_7_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_2 = I_7_0_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0_0,
  input  [7:0] I_0_0_0_1,
  input  [7:0] I_0_0_0_2,
  input  [7:0] I_0_0_1_0,
  input  [7:0] I_0_0_1_1,
  input  [7:0] I_0_0_1_2,
  input  [7:0] I_0_0_2_0,
  input  [7:0] I_0_0_2_1,
  input  [7:0] I_0_0_2_2,
  input  [7:0] I_1_0_0_0,
  input  [7:0] I_1_0_0_1,
  input  [7:0] I_1_0_0_2,
  input  [7:0] I_1_0_1_0,
  input  [7:0] I_1_0_1_1,
  input  [7:0] I_1_0_1_2,
  input  [7:0] I_1_0_2_0,
  input  [7:0] I_1_0_2_1,
  input  [7:0] I_1_0_2_2,
  input  [7:0] I_2_0_0_0,
  input  [7:0] I_2_0_0_1,
  input  [7:0] I_2_0_0_2,
  input  [7:0] I_2_0_1_0,
  input  [7:0] I_2_0_1_1,
  input  [7:0] I_2_0_1_2,
  input  [7:0] I_2_0_2_0,
  input  [7:0] I_2_0_2_1,
  input  [7:0] I_2_0_2_2,
  input  [7:0] I_3_0_0_0,
  input  [7:0] I_3_0_0_1,
  input  [7:0] I_3_0_0_2,
  input  [7:0] I_3_0_1_0,
  input  [7:0] I_3_0_1_1,
  input  [7:0] I_3_0_1_2,
  input  [7:0] I_3_0_2_0,
  input  [7:0] I_3_0_2_1,
  input  [7:0] I_3_0_2_2,
  input  [7:0] I_4_0_0_0,
  input  [7:0] I_4_0_0_1,
  input  [7:0] I_4_0_0_2,
  input  [7:0] I_4_0_1_0,
  input  [7:0] I_4_0_1_1,
  input  [7:0] I_4_0_1_2,
  input  [7:0] I_4_0_2_0,
  input  [7:0] I_4_0_2_1,
  input  [7:0] I_4_0_2_2,
  input  [7:0] I_5_0_0_0,
  input  [7:0] I_5_0_0_1,
  input  [7:0] I_5_0_0_2,
  input  [7:0] I_5_0_1_0,
  input  [7:0] I_5_0_1_1,
  input  [7:0] I_5_0_1_2,
  input  [7:0] I_5_0_2_0,
  input  [7:0] I_5_0_2_1,
  input  [7:0] I_5_0_2_2,
  input  [7:0] I_6_0_0_0,
  input  [7:0] I_6_0_0_1,
  input  [7:0] I_6_0_0_2,
  input  [7:0] I_6_0_1_0,
  input  [7:0] I_6_0_1_1,
  input  [7:0] I_6_0_1_2,
  input  [7:0] I_6_0_2_0,
  input  [7:0] I_6_0_2_1,
  input  [7:0] I_6_0_2_2,
  input  [7:0] I_7_0_0_0,
  input  [7:0] I_7_0_0_1,
  input  [7:0] I_7_0_0_2,
  input  [7:0] I_7_0_1_0,
  input  [7:0] I_7_0_1_1,
  input  [7:0] I_7_0_1_2,
  input  [7:0] I_7_0_2_0,
  input  [7:0] I_7_0_2_1,
  input  [7:0] I_7_0_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_1_2_0,
  output [7:0] O_1_2_1,
  output [7:0] O_1_2_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_2_1_2,
  output [7:0] O_2_2_0,
  output [7:0] O_2_2_1,
  output [7:0] O_2_2_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_3_1_2,
  output [7:0] O_3_2_0,
  output [7:0] O_3_2_1,
  output [7:0] O_3_2_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_4_1_2,
  output [7:0] O_4_2_0,
  output [7:0] O_4_2_1,
  output [7:0] O_4_2_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_5_1_2,
  output [7:0] O_5_2_0,
  output [7:0] O_5_2_1,
  output [7:0] O_5_2_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_6_1_2,
  output [7:0] O_6_2_0,
  output [7:0] O_6_2_1,
  output [7:0] O_6_2_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_7_1_2,
  output [7:0] O_7_2_0,
  output [7:0] O_7_2_1,
  output [7:0] O_7_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_2_2; // @[MapT.scala 8:20]
  MapS_6 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0_0(op_I_0_0_0_0),
    .I_0_0_0_1(op_I_0_0_0_1),
    .I_0_0_0_2(op_I_0_0_0_2),
    .I_0_0_1_0(op_I_0_0_1_0),
    .I_0_0_1_1(op_I_0_0_1_1),
    .I_0_0_1_2(op_I_0_0_1_2),
    .I_0_0_2_0(op_I_0_0_2_0),
    .I_0_0_2_1(op_I_0_0_2_1),
    .I_0_0_2_2(op_I_0_0_2_2),
    .I_1_0_0_0(op_I_1_0_0_0),
    .I_1_0_0_1(op_I_1_0_0_1),
    .I_1_0_0_2(op_I_1_0_0_2),
    .I_1_0_1_0(op_I_1_0_1_0),
    .I_1_0_1_1(op_I_1_0_1_1),
    .I_1_0_1_2(op_I_1_0_1_2),
    .I_1_0_2_0(op_I_1_0_2_0),
    .I_1_0_2_1(op_I_1_0_2_1),
    .I_1_0_2_2(op_I_1_0_2_2),
    .I_2_0_0_0(op_I_2_0_0_0),
    .I_2_0_0_1(op_I_2_0_0_1),
    .I_2_0_0_2(op_I_2_0_0_2),
    .I_2_0_1_0(op_I_2_0_1_0),
    .I_2_0_1_1(op_I_2_0_1_1),
    .I_2_0_1_2(op_I_2_0_1_2),
    .I_2_0_2_0(op_I_2_0_2_0),
    .I_2_0_2_1(op_I_2_0_2_1),
    .I_2_0_2_2(op_I_2_0_2_2),
    .I_3_0_0_0(op_I_3_0_0_0),
    .I_3_0_0_1(op_I_3_0_0_1),
    .I_3_0_0_2(op_I_3_0_0_2),
    .I_3_0_1_0(op_I_3_0_1_0),
    .I_3_0_1_1(op_I_3_0_1_1),
    .I_3_0_1_2(op_I_3_0_1_2),
    .I_3_0_2_0(op_I_3_0_2_0),
    .I_3_0_2_1(op_I_3_0_2_1),
    .I_3_0_2_2(op_I_3_0_2_2),
    .I_4_0_0_0(op_I_4_0_0_0),
    .I_4_0_0_1(op_I_4_0_0_1),
    .I_4_0_0_2(op_I_4_0_0_2),
    .I_4_0_1_0(op_I_4_0_1_0),
    .I_4_0_1_1(op_I_4_0_1_1),
    .I_4_0_1_2(op_I_4_0_1_2),
    .I_4_0_2_0(op_I_4_0_2_0),
    .I_4_0_2_1(op_I_4_0_2_1),
    .I_4_0_2_2(op_I_4_0_2_2),
    .I_5_0_0_0(op_I_5_0_0_0),
    .I_5_0_0_1(op_I_5_0_0_1),
    .I_5_0_0_2(op_I_5_0_0_2),
    .I_5_0_1_0(op_I_5_0_1_0),
    .I_5_0_1_1(op_I_5_0_1_1),
    .I_5_0_1_2(op_I_5_0_1_2),
    .I_5_0_2_0(op_I_5_0_2_0),
    .I_5_0_2_1(op_I_5_0_2_1),
    .I_5_0_2_2(op_I_5_0_2_2),
    .I_6_0_0_0(op_I_6_0_0_0),
    .I_6_0_0_1(op_I_6_0_0_1),
    .I_6_0_0_2(op_I_6_0_0_2),
    .I_6_0_1_0(op_I_6_0_1_0),
    .I_6_0_1_1(op_I_6_0_1_1),
    .I_6_0_1_2(op_I_6_0_1_2),
    .I_6_0_2_0(op_I_6_0_2_0),
    .I_6_0_2_1(op_I_6_0_2_1),
    .I_6_0_2_2(op_I_6_0_2_2),
    .I_7_0_0_0(op_I_7_0_0_0),
    .I_7_0_0_1(op_I_7_0_0_1),
    .I_7_0_0_2(op_I_7_0_0_2),
    .I_7_0_1_0(op_I_7_0_1_0),
    .I_7_0_1_1(op_I_7_0_1_1),
    .I_7_0_1_2(op_I_7_0_1_2),
    .I_7_0_2_0(op_I_7_0_2_0),
    .I_7_0_2_1(op_I_7_0_2_1),
    .I_7_0_2_2(op_I_7_0_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_2_2_0(op_O_2_2_0),
    .O_2_2_1(op_O_2_2_1),
    .O_2_2_2(op_O_2_2_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_3_2_0(op_O_3_2_0),
    .O_3_2_1(op_O_3_2_1),
    .O_3_2_2(op_O_3_2_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_4_2_0(op_O_4_2_0),
    .O_4_2_1(op_O_4_2_1),
    .O_4_2_2(op_O_4_2_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_5_2_0(op_O_5_2_0),
    .O_5_2_1(op_O_5_2_1),
    .O_5_2_2(op_O_5_2_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_6_2_0(op_O_6_2_0),
    .O_6_2_1(op_O_6_2_1),
    .O_6_2_2(op_O_6_2_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2),
    .O_7_2_0(op_O_7_2_0),
    .O_7_2_1(op_O_7_2_1),
    .O_7_2_2(op_O_7_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_0_1_0 = op_O_0_1_0; // @[MapT.scala 15:7]
  assign O_0_1_1 = op_O_0_1_1; // @[MapT.scala 15:7]
  assign O_0_1_2 = op_O_0_1_2; // @[MapT.scala 15:7]
  assign O_0_2_0 = op_O_0_2_0; // @[MapT.scala 15:7]
  assign O_0_2_1 = op_O_0_2_1; // @[MapT.scala 15:7]
  assign O_0_2_2 = op_O_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_1_1_0 = op_O_1_1_0; // @[MapT.scala 15:7]
  assign O_1_1_1 = op_O_1_1_1; // @[MapT.scala 15:7]
  assign O_1_1_2 = op_O_1_1_2; // @[MapT.scala 15:7]
  assign O_1_2_0 = op_O_1_2_0; // @[MapT.scala 15:7]
  assign O_1_2_1 = op_O_1_2_1; // @[MapT.scala 15:7]
  assign O_1_2_2 = op_O_1_2_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_2_1_0 = op_O_2_1_0; // @[MapT.scala 15:7]
  assign O_2_1_1 = op_O_2_1_1; // @[MapT.scala 15:7]
  assign O_2_1_2 = op_O_2_1_2; // @[MapT.scala 15:7]
  assign O_2_2_0 = op_O_2_2_0; // @[MapT.scala 15:7]
  assign O_2_2_1 = op_O_2_2_1; // @[MapT.scala 15:7]
  assign O_2_2_2 = op_O_2_2_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign O_3_1_0 = op_O_3_1_0; // @[MapT.scala 15:7]
  assign O_3_1_1 = op_O_3_1_1; // @[MapT.scala 15:7]
  assign O_3_1_2 = op_O_3_1_2; // @[MapT.scala 15:7]
  assign O_3_2_0 = op_O_3_2_0; // @[MapT.scala 15:7]
  assign O_3_2_1 = op_O_3_2_1; // @[MapT.scala 15:7]
  assign O_3_2_2 = op_O_3_2_2; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_4_0_2 = op_O_4_0_2; // @[MapT.scala 15:7]
  assign O_4_1_0 = op_O_4_1_0; // @[MapT.scala 15:7]
  assign O_4_1_1 = op_O_4_1_1; // @[MapT.scala 15:7]
  assign O_4_1_2 = op_O_4_1_2; // @[MapT.scala 15:7]
  assign O_4_2_0 = op_O_4_2_0; // @[MapT.scala 15:7]
  assign O_4_2_1 = op_O_4_2_1; // @[MapT.scala 15:7]
  assign O_4_2_2 = op_O_4_2_2; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_5_0_2 = op_O_5_0_2; // @[MapT.scala 15:7]
  assign O_5_1_0 = op_O_5_1_0; // @[MapT.scala 15:7]
  assign O_5_1_1 = op_O_5_1_1; // @[MapT.scala 15:7]
  assign O_5_1_2 = op_O_5_1_2; // @[MapT.scala 15:7]
  assign O_5_2_0 = op_O_5_2_0; // @[MapT.scala 15:7]
  assign O_5_2_1 = op_O_5_2_1; // @[MapT.scala 15:7]
  assign O_5_2_2 = op_O_5_2_2; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_6_0_2 = op_O_6_0_2; // @[MapT.scala 15:7]
  assign O_6_1_0 = op_O_6_1_0; // @[MapT.scala 15:7]
  assign O_6_1_1 = op_O_6_1_1; // @[MapT.scala 15:7]
  assign O_6_1_2 = op_O_6_1_2; // @[MapT.scala 15:7]
  assign O_6_2_0 = op_O_6_2_0; // @[MapT.scala 15:7]
  assign O_6_2_1 = op_O_6_2_1; // @[MapT.scala 15:7]
  assign O_6_2_2 = op_O_6_2_2; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_7_0_2 = op_O_7_0_2; // @[MapT.scala 15:7]
  assign O_7_1_0 = op_O_7_1_0; // @[MapT.scala 15:7]
  assign O_7_1_1 = op_O_7_1_1; // @[MapT.scala 15:7]
  assign O_7_1_2 = op_O_7_1_2; // @[MapT.scala 15:7]
  assign O_7_2_0 = op_O_7_2_0; // @[MapT.scala 15:7]
  assign O_7_2_1 = op_O_7_2_1; // @[MapT.scala 15:7]
  assign O_7_2_2 = op_O_7_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0_0 = I_0_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_0_1 = I_0_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_0_2 = I_0_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_0_1_0 = I_0_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1_1 = I_0_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_0_1_2 = I_0_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_0_2_0 = I_0_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_0_2_1 = I_0_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2_2 = I_0_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0_0 = I_1_0_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_0_1 = I_1_0_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0_2 = I_1_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_1_0 = I_1_0_1_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1_1 = I_1_0_1_1; // @[MapT.scala 14:10]
  assign op_I_1_0_1_2 = I_1_0_1_2; // @[MapT.scala 14:10]
  assign op_I_1_0_2_0 = I_1_0_2_0; // @[MapT.scala 14:10]
  assign op_I_1_0_2_1 = I_1_0_2_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2_2 = I_1_0_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0_0 = I_2_0_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_0_1 = I_2_0_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0_2 = I_2_0_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_1_0 = I_2_0_1_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1_1 = I_2_0_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0_1_2 = I_2_0_1_2; // @[MapT.scala 14:10]
  assign op_I_2_0_2_0 = I_2_0_2_0; // @[MapT.scala 14:10]
  assign op_I_2_0_2_1 = I_2_0_2_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2_2 = I_2_0_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0_0 = I_3_0_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_0_1 = I_3_0_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0_2 = I_3_0_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_1_0 = I_3_0_1_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1_1 = I_3_0_1_1; // @[MapT.scala 14:10]
  assign op_I_3_0_1_2 = I_3_0_1_2; // @[MapT.scala 14:10]
  assign op_I_3_0_2_0 = I_3_0_2_0; // @[MapT.scala 14:10]
  assign op_I_3_0_2_1 = I_3_0_2_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2_2 = I_3_0_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0_0 = I_4_0_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_0_1 = I_4_0_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_0_2 = I_4_0_0_2; // @[MapT.scala 14:10]
  assign op_I_4_0_1_0 = I_4_0_1_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1_1 = I_4_0_1_1; // @[MapT.scala 14:10]
  assign op_I_4_0_1_2 = I_4_0_1_2; // @[MapT.scala 14:10]
  assign op_I_4_0_2_0 = I_4_0_2_0; // @[MapT.scala 14:10]
  assign op_I_4_0_2_1 = I_4_0_2_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2_2 = I_4_0_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0_0 = I_5_0_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_0_1 = I_5_0_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_0_2 = I_5_0_0_2; // @[MapT.scala 14:10]
  assign op_I_5_0_1_0 = I_5_0_1_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1_1 = I_5_0_1_1; // @[MapT.scala 14:10]
  assign op_I_5_0_1_2 = I_5_0_1_2; // @[MapT.scala 14:10]
  assign op_I_5_0_2_0 = I_5_0_2_0; // @[MapT.scala 14:10]
  assign op_I_5_0_2_1 = I_5_0_2_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2_2 = I_5_0_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0_0 = I_6_0_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_0_1 = I_6_0_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_0_2 = I_6_0_0_2; // @[MapT.scala 14:10]
  assign op_I_6_0_1_0 = I_6_0_1_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1_1 = I_6_0_1_1; // @[MapT.scala 14:10]
  assign op_I_6_0_1_2 = I_6_0_1_2; // @[MapT.scala 14:10]
  assign op_I_6_0_2_0 = I_6_0_2_0; // @[MapT.scala 14:10]
  assign op_I_6_0_2_1 = I_6_0_2_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2_2 = I_6_0_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0_0 = I_7_0_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_0_1 = I_7_0_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_0_2 = I_7_0_0_2; // @[MapT.scala 14:10]
  assign op_I_7_0_1_0 = I_7_0_1_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1_1 = I_7_0_1_1; // @[MapT.scala 14:10]
  assign op_I_7_0_1_2 = I_7_0_1_2; // @[MapT.scala 14:10]
  assign op_I_7_0_2_0 = I_7_0_2_0; // @[MapT.scala 14:10]
  assign op_I_7_0_2_1 = I_7_0_2_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2_2 = I_7_0_2_2; // @[MapT.scala 14:10]
endmodule
module InitialDelayCounter(
  input   clock,
  input   reset,
  output  valid_down
);
  reg  value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire  _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 1'h1; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 1'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 1'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module AtomTuple(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_t0b,
  output [7:0] O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Map2S_22(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_t0b,
  output [7:0] O_0_t1b,
  output [7:0] O_1_t0b,
  output [7:0] O_1_t1b,
  output [7:0] O_2_t0b,
  output [7:0] O_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  AtomTuple other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  AtomTuple other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_t0b(other_ops_1_O_t0b),
    .O_t1b(other_ops_1_O_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign O_2_t0b = other_ops_1_O_t0b; // @[Map2S.scala 24:12]
  assign O_2_t1b = other_ops_1_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
endmodule
module Map2S_23(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_1_2,
  input  [7:0] I0_2_0,
  input  [7:0] I0_2_1,
  input  [7:0] I0_2_2,
  output [7:0] O_0_0_t0b,
  output [7:0] O_0_0_t1b,
  output [7:0] O_0_1_t0b,
  output [7:0] O_0_1_t1b,
  output [7:0] O_0_2_t0b,
  output [7:0] O_0_2_t1b,
  output [7:0] O_1_0_t0b,
  output [7:0] O_1_0_t1b,
  output [7:0] O_1_1_t0b,
  output [7:0] O_1_1_t1b,
  output [7:0] O_1_2_t0b,
  output [7:0] O_1_2_t1b,
  output [7:0] O_2_0_t0b,
  output [7:0] O_2_0_t1b,
  output [7:0] O_2_1_t0b,
  output [7:0] O_2_1_t1b,
  output [7:0] O_2_2_t0b,
  output [7:0] O_2_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_t1b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  Map2S_22 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b),
    .O_1_t0b(fst_op_O_1_t0b),
    .O_1_t1b(fst_op_O_1_t1b),
    .O_2_t0b(fst_op_O_2_t0b),
    .O_2_t1b(fst_op_O_2_t1b)
  );
  Map2S_22 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_t0b(other_ops_0_O_0_t0b),
    .O_0_t1b(other_ops_0_O_0_t1b),
    .O_1_t0b(other_ops_0_O_1_t0b),
    .O_1_t1b(other_ops_0_O_1_t1b),
    .O_2_t0b(other_ops_0_O_2_t0b),
    .O_2_t1b(other_ops_0_O_2_t1b)
  );
  Map2S_22 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_t0b(other_ops_1_O_0_t0b),
    .O_0_t1b(other_ops_1_O_0_t1b),
    .O_1_t0b(other_ops_1_O_1_t0b),
    .O_1_t1b(other_ops_1_O_1_t1b),
    .O_2_t0b(other_ops_1_O_2_t0b),
    .O_2_t1b(other_ops_1_O_2_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign O_0_1_t0b = fst_op_O_1_t0b; // @[Map2S.scala 19:8]
  assign O_0_1_t1b = fst_op_O_1_t1b; // @[Map2S.scala 19:8]
  assign O_0_2_t0b = fst_op_O_2_t0b; // @[Map2S.scala 19:8]
  assign O_0_2_t1b = fst_op_O_2_t1b; // @[Map2S.scala 19:8]
  assign O_1_0_t0b = other_ops_0_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_1_0_t1b = other_ops_0_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_1_1_t0b = other_ops_0_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_1_1_t1b = other_ops_0_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_1_2_t0b = other_ops_0_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_1_2_t1b = other_ops_0_O_2_t1b; // @[Map2S.scala 24:12]
  assign O_2_0_t0b = other_ops_1_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_2_0_t1b = other_ops_1_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_2_1_t0b = other_ops_1_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_2_1_t1b = other_ops_1_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_2_2_t0b = other_ops_1_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_2_2_t1b = other_ops_1_O_2_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = 8'h0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = 8'h1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = 8'h0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = 8'h2; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = 8'h0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = 8'h0; // @[Map2S.scala 23:43]
endmodule
module LShift(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  wire [262:0] _GEN_0; // @[Arithmetic.scala 163:23]
  wire [262:0] _T; // @[Arithmetic.scala 163:23]
  assign _GEN_0 = {{255'd0}, I_t0b}; // @[Arithmetic.scala 163:23]
  assign _T = _GEN_0 << I_t1b; // @[Arithmetic.scala 163:23]
  assign valid_down = valid_up; // @[Arithmetic.scala 164:14]
  assign O = _T[7:0]; // @[Arithmetic.scala 163:5]
endmodule
module MapS_7(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  input  [7:0] I_1_t0b,
  input  [7:0] I_1_t1b,
  input  [7:0] I_2_t0b,
  input  [7:0] I_2_t1b,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  LShift fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  LShift other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t0b(other_ops_0_I_t0b),
    .I_t1b(other_ops_0_I_t1b),
    .O(other_ops_0_O)
  );
  LShift other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_t0b(other_ops_1_I_t0b),
    .I_t1b(other_ops_1_I_t1b),
    .O(other_ops_1_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t0b = I_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_t1b = I_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_t0b = I_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_t1b = I_2_t1b; // @[MapS.scala 20:41]
endmodule
module MapS_8(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_t0b,
  input  [7:0] I_0_0_t1b,
  input  [7:0] I_0_1_t0b,
  input  [7:0] I_0_1_t1b,
  input  [7:0] I_0_2_t0b,
  input  [7:0] I_0_2_t1b,
  input  [7:0] I_1_0_t0b,
  input  [7:0] I_1_0_t1b,
  input  [7:0] I_1_1_t0b,
  input  [7:0] I_1_1_t1b,
  input  [7:0] I_1_2_t0b,
  input  [7:0] I_1_2_t1b,
  input  [7:0] I_2_0_t0b,
  input  [7:0] I_2_0_t1b,
  input  [7:0] I_2_1_t0b,
  input  [7:0] I_2_1_t1b,
  input  [7:0] I_2_2_t0b,
  input  [7:0] I_2_2_t1b,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  MapS_7 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .I_1_t0b(fst_op_I_1_t0b),
    .I_1_t1b(fst_op_I_1_t1b),
    .I_2_t0b(fst_op_I_2_t0b),
    .I_2_t1b(fst_op_I_2_t1b),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  MapS_7 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_t0b(other_ops_0_I_0_t0b),
    .I_0_t1b(other_ops_0_I_0_t1b),
    .I_1_t0b(other_ops_0_I_1_t0b),
    .I_1_t1b(other_ops_0_I_1_t1b),
    .I_2_t0b(other_ops_0_I_2_t0b),
    .I_2_t1b(other_ops_0_I_2_t1b),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  MapS_7 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_t0b(other_ops_1_I_0_t0b),
    .I_0_t1b(other_ops_1_I_0_t1b),
    .I_1_t0b(other_ops_1_I_1_t0b),
    .I_1_t1b(other_ops_1_I_1_t1b),
    .I_2_t0b(other_ops_1_I_2_t0b),
    .I_2_t1b(other_ops_1_I_2_t1b),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t0b = I_0_1_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t1b = I_0_1_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t0b = I_0_2_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t1b = I_0_2_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_t0b = I_1_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_t1b = I_1_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t0b = I_1_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t1b = I_1_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t0b = I_1_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t1b = I_1_2_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_t0b = I_2_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_t1b = I_2_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t0b = I_2_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t1b = I_2_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t0b = I_2_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t1b = I_2_2_t1b; // @[MapS.scala 20:41]
endmodule
module AddNoValid(
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  assign O = I_t0b + I_t1b; // @[Arithmetic.scala 69:5]
endmodule
module ReduceS(
  input        clock,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O_0
);
  wire [7:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_1_O; // @[ReduceS.scala 20:43]
  reg [7:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_1;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  AddNoValid AddNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_1_I_t0b),
    .I_t1b(AddNoValid_1_I_t1b),
    .O(AddNoValid_1_O)
  );
  assign valid_down = _T_1; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = I_1; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = AddNoValid_1_O; // @[ReduceS.scala 36:18]
  assign AddNoValid_1_I_t0b = I_0; // @[ReduceS.scala 43:18]
  assign AddNoValid_1_I_t1b = I_2; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    _T_1 <= valid_up;
  end
endmodule
module MapS_9(
  input        clock,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  output [7:0] O_0_0,
  output [7:0] O_1_0,
  output [7:0] O_2_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  ReduceS fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .O_0(fst_op_O_0)
  );
  ReduceS other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0(other_ops_0_I_0),
    .I_1(other_ops_0_I_1),
    .I_2(other_ops_0_I_2),
    .O_0(other_ops_0_O_0)
  );
  ReduceS other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0(other_ops_1_I_0),
    .I_1(other_ops_1_I_1),
    .I_2(other_ops_1_I_2),
    .O_0(other_ops_1_O_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0 = I_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1 = I_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2 = I_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0 = I_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1 = I_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2 = I_2_2; // @[MapS.scala 20:41]
endmodule
module MapSNoValid(
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  output [7:0] O_0
);
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 28:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 28:22]
  wire [7:0] fst_op_O; // @[MapS.scala 28:22]
  AddNoValid fst_op ( // @[MapS.scala 28:22]
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign O_0 = fst_op_O; // @[MapS.scala 35:8]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 34:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 34:12]
endmodule
module ReduceS_1(
  input        clock,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_1_0,
  input  [7:0] I_2_0,
  output [7:0] O_0_0
);
  wire [7:0] MapSNoValid_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_O_0; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_1_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_1_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_1_O_0; // @[ReduceS.scala 20:43]
  reg [7:0] _T_0; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_1;
  MapSNoValid MapSNoValid ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_I_0_t0b),
    .I_0_t1b(MapSNoValid_I_0_t1b),
    .O_0(MapSNoValid_O_0)
  );
  MapSNoValid MapSNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_1_I_0_t0b),
    .I_0_t1b(MapSNoValid_1_I_0_t1b),
    .O_0(MapSNoValid_1_O_0)
  );
  assign valid_down = _T_1; // @[ReduceS.scala 47:14]
  assign O_0_0 = _T_0; // @[ReduceS.scala 27:14]
  assign MapSNoValid_I_0_t0b = I_2_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_I_0_t1b = MapSNoValid_1_O_0; // @[ReduceS.scala 36:18]
  assign MapSNoValid_1_I_0_t0b = I_0_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_1_I_0_t1b = I_1_0; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= MapSNoValid_O_0;
    _T_1 <= valid_up;
  end
endmodule
module InitialDelayCounter_1(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [1:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [1:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 2'h3; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 2'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 2'h3; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 2'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Map2S_24(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  output [7:0] O_0_t0b,
  output [7:0] O_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = 8'h4; // @[Map2S.scala 18:13]
endmodule
module Map2S_25(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  output [7:0] O_0_0_t0b,
  output [7:0] O_0_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  Map2S_24 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
endmodule
module RShift(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 143:14]
  assign O = I_t0b >> I_t1b; // @[Arithmetic.scala 142:5]
endmodule
module MapS_10(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  output [7:0] O_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  RShift fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
endmodule
module MapS_11(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_t0b,
  input  [7:0] I_0_0_t1b,
  output [7:0] O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  MapS_10 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
endmodule
module Module_0(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  output [7:0] O_0_0
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n146_valid_up; // @[Top.scala 16:22]
  wire  n146_valid_down; // @[Top.scala 16:22]
  wire [7:0] n146_I0_0_0; // @[Top.scala 16:22]
  wire [7:0] n146_I0_0_1; // @[Top.scala 16:22]
  wire [7:0] n146_I0_0_2; // @[Top.scala 16:22]
  wire [7:0] n146_I0_1_0; // @[Top.scala 16:22]
  wire [7:0] n146_I0_1_1; // @[Top.scala 16:22]
  wire [7:0] n146_I0_1_2; // @[Top.scala 16:22]
  wire [7:0] n146_I0_2_0; // @[Top.scala 16:22]
  wire [7:0] n146_I0_2_1; // @[Top.scala 16:22]
  wire [7:0] n146_I0_2_2; // @[Top.scala 16:22]
  wire [7:0] n146_O_0_0_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_0_0_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_0_1_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_0_1_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_0_2_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_0_2_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_1_0_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_1_0_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_1_1_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_1_1_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_1_2_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_1_2_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_2_0_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_2_0_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_2_1_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_2_1_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_2_2_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_2_2_t1b; // @[Top.scala 16:22]
  wire  n157_valid_up; // @[Top.scala 20:22]
  wire  n157_valid_down; // @[Top.scala 20:22]
  wire [7:0] n157_I_0_0_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_0_0_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_0_1_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_0_1_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_0_2_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_0_2_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_1_0_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_1_0_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_1_1_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_1_1_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_1_2_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_1_2_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_2_0_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_2_0_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_2_1_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_2_1_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_2_2_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_2_2_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_O_0_0; // @[Top.scala 20:22]
  wire [7:0] n157_O_0_1; // @[Top.scala 20:22]
  wire [7:0] n157_O_0_2; // @[Top.scala 20:22]
  wire [7:0] n157_O_1_0; // @[Top.scala 20:22]
  wire [7:0] n157_O_1_1; // @[Top.scala 20:22]
  wire [7:0] n157_O_1_2; // @[Top.scala 20:22]
  wire [7:0] n157_O_2_0; // @[Top.scala 20:22]
  wire [7:0] n157_O_2_1; // @[Top.scala 20:22]
  wire [7:0] n157_O_2_2; // @[Top.scala 20:22]
  wire  n162_clock; // @[Top.scala 23:22]
  wire  n162_valid_up; // @[Top.scala 23:22]
  wire  n162_valid_down; // @[Top.scala 23:22]
  wire [7:0] n162_I_0_0; // @[Top.scala 23:22]
  wire [7:0] n162_I_0_1; // @[Top.scala 23:22]
  wire [7:0] n162_I_0_2; // @[Top.scala 23:22]
  wire [7:0] n162_I_1_0; // @[Top.scala 23:22]
  wire [7:0] n162_I_1_1; // @[Top.scala 23:22]
  wire [7:0] n162_I_1_2; // @[Top.scala 23:22]
  wire [7:0] n162_I_2_0; // @[Top.scala 23:22]
  wire [7:0] n162_I_2_1; // @[Top.scala 23:22]
  wire [7:0] n162_I_2_2; // @[Top.scala 23:22]
  wire [7:0] n162_O_0_0; // @[Top.scala 23:22]
  wire [7:0] n162_O_1_0; // @[Top.scala 23:22]
  wire [7:0] n162_O_2_0; // @[Top.scala 23:22]
  wire  n167_clock; // @[Top.scala 26:22]
  wire  n167_valid_up; // @[Top.scala 26:22]
  wire  n167_valid_down; // @[Top.scala 26:22]
  wire [7:0] n167_I_0_0; // @[Top.scala 26:22]
  wire [7:0] n167_I_1_0; // @[Top.scala 26:22]
  wire [7:0] n167_I_2_0; // @[Top.scala 26:22]
  wire [7:0] n167_O_0_0; // @[Top.scala 26:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n170_valid_up; // @[Top.scala 30:22]
  wire  n170_valid_down; // @[Top.scala 30:22]
  wire [7:0] n170_I0_0_0; // @[Top.scala 30:22]
  wire [7:0] n170_O_0_0_t0b; // @[Top.scala 30:22]
  wire [7:0] n170_O_0_0_t1b; // @[Top.scala 30:22]
  wire  n181_valid_up; // @[Top.scala 34:22]
  wire  n181_valid_down; // @[Top.scala 34:22]
  wire [7:0] n181_I_0_0_t0b; // @[Top.scala 34:22]
  wire [7:0] n181_I_0_0_t1b; // @[Top.scala 34:22]
  wire [7:0] n181_O_0_0; // @[Top.scala 34:22]
  InitialDelayCounter InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  Map2S_23 n146 ( // @[Top.scala 16:22]
    .valid_up(n146_valid_up),
    .valid_down(n146_valid_down),
    .I0_0_0(n146_I0_0_0),
    .I0_0_1(n146_I0_0_1),
    .I0_0_2(n146_I0_0_2),
    .I0_1_0(n146_I0_1_0),
    .I0_1_1(n146_I0_1_1),
    .I0_1_2(n146_I0_1_2),
    .I0_2_0(n146_I0_2_0),
    .I0_2_1(n146_I0_2_1),
    .I0_2_2(n146_I0_2_2),
    .O_0_0_t0b(n146_O_0_0_t0b),
    .O_0_0_t1b(n146_O_0_0_t1b),
    .O_0_1_t0b(n146_O_0_1_t0b),
    .O_0_1_t1b(n146_O_0_1_t1b),
    .O_0_2_t0b(n146_O_0_2_t0b),
    .O_0_2_t1b(n146_O_0_2_t1b),
    .O_1_0_t0b(n146_O_1_0_t0b),
    .O_1_0_t1b(n146_O_1_0_t1b),
    .O_1_1_t0b(n146_O_1_1_t0b),
    .O_1_1_t1b(n146_O_1_1_t1b),
    .O_1_2_t0b(n146_O_1_2_t0b),
    .O_1_2_t1b(n146_O_1_2_t1b),
    .O_2_0_t0b(n146_O_2_0_t0b),
    .O_2_0_t1b(n146_O_2_0_t1b),
    .O_2_1_t0b(n146_O_2_1_t0b),
    .O_2_1_t1b(n146_O_2_1_t1b),
    .O_2_2_t0b(n146_O_2_2_t0b),
    .O_2_2_t1b(n146_O_2_2_t1b)
  );
  MapS_8 n157 ( // @[Top.scala 20:22]
    .valid_up(n157_valid_up),
    .valid_down(n157_valid_down),
    .I_0_0_t0b(n157_I_0_0_t0b),
    .I_0_0_t1b(n157_I_0_0_t1b),
    .I_0_1_t0b(n157_I_0_1_t0b),
    .I_0_1_t1b(n157_I_0_1_t1b),
    .I_0_2_t0b(n157_I_0_2_t0b),
    .I_0_2_t1b(n157_I_0_2_t1b),
    .I_1_0_t0b(n157_I_1_0_t0b),
    .I_1_0_t1b(n157_I_1_0_t1b),
    .I_1_1_t0b(n157_I_1_1_t0b),
    .I_1_1_t1b(n157_I_1_1_t1b),
    .I_1_2_t0b(n157_I_1_2_t0b),
    .I_1_2_t1b(n157_I_1_2_t1b),
    .I_2_0_t0b(n157_I_2_0_t0b),
    .I_2_0_t1b(n157_I_2_0_t1b),
    .I_2_1_t0b(n157_I_2_1_t0b),
    .I_2_1_t1b(n157_I_2_1_t1b),
    .I_2_2_t0b(n157_I_2_2_t0b),
    .I_2_2_t1b(n157_I_2_2_t1b),
    .O_0_0(n157_O_0_0),
    .O_0_1(n157_O_0_1),
    .O_0_2(n157_O_0_2),
    .O_1_0(n157_O_1_0),
    .O_1_1(n157_O_1_1),
    .O_1_2(n157_O_1_2),
    .O_2_0(n157_O_2_0),
    .O_2_1(n157_O_2_1),
    .O_2_2(n157_O_2_2)
  );
  MapS_9 n162 ( // @[Top.scala 23:22]
    .clock(n162_clock),
    .valid_up(n162_valid_up),
    .valid_down(n162_valid_down),
    .I_0_0(n162_I_0_0),
    .I_0_1(n162_I_0_1),
    .I_0_2(n162_I_0_2),
    .I_1_0(n162_I_1_0),
    .I_1_1(n162_I_1_1),
    .I_1_2(n162_I_1_2),
    .I_2_0(n162_I_2_0),
    .I_2_1(n162_I_2_1),
    .I_2_2(n162_I_2_2),
    .O_0_0(n162_O_0_0),
    .O_1_0(n162_O_1_0),
    .O_2_0(n162_O_2_0)
  );
  ReduceS_1 n167 ( // @[Top.scala 26:22]
    .clock(n167_clock),
    .valid_up(n167_valid_up),
    .valid_down(n167_valid_down),
    .I_0_0(n167_I_0_0),
    .I_1_0(n167_I_1_0),
    .I_2_0(n167_I_2_0),
    .O_0_0(n167_O_0_0)
  );
  InitialDelayCounter_1 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  Map2S_25 n170 ( // @[Top.scala 30:22]
    .valid_up(n170_valid_up),
    .valid_down(n170_valid_down),
    .I0_0_0(n170_I0_0_0),
    .O_0_0_t0b(n170_O_0_0_t0b),
    .O_0_0_t1b(n170_O_0_0_t1b)
  );
  MapS_11 n181 ( // @[Top.scala 34:22]
    .valid_up(n181_valid_up),
    .valid_down(n181_valid_down),
    .I_0_0_t0b(n181_I_0_0_t0b),
    .I_0_0_t1b(n181_I_0_0_t1b),
    .O_0_0(n181_O_0_0)
  );
  assign valid_down = n181_valid_down; // @[Top.scala 38:16]
  assign O_0_0 = n181_O_0_0; // @[Top.scala 37:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n146_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 19:19]
  assign n146_I0_0_0 = I_0_0; // @[Top.scala 17:13]
  assign n146_I0_0_1 = I_0_1; // @[Top.scala 17:13]
  assign n146_I0_0_2 = I_0_2; // @[Top.scala 17:13]
  assign n146_I0_1_0 = I_1_0; // @[Top.scala 17:13]
  assign n146_I0_1_1 = I_1_1; // @[Top.scala 17:13]
  assign n146_I0_1_2 = I_1_2; // @[Top.scala 17:13]
  assign n146_I0_2_0 = I_2_0; // @[Top.scala 17:13]
  assign n146_I0_2_1 = I_2_1; // @[Top.scala 17:13]
  assign n146_I0_2_2 = I_2_2; // @[Top.scala 17:13]
  assign n157_valid_up = n146_valid_down; // @[Top.scala 22:19]
  assign n157_I_0_0_t0b = n146_O_0_0_t0b; // @[Top.scala 21:12]
  assign n157_I_0_0_t1b = n146_O_0_0_t1b; // @[Top.scala 21:12]
  assign n157_I_0_1_t0b = n146_O_0_1_t0b; // @[Top.scala 21:12]
  assign n157_I_0_1_t1b = n146_O_0_1_t1b; // @[Top.scala 21:12]
  assign n157_I_0_2_t0b = n146_O_0_2_t0b; // @[Top.scala 21:12]
  assign n157_I_0_2_t1b = n146_O_0_2_t1b; // @[Top.scala 21:12]
  assign n157_I_1_0_t0b = n146_O_1_0_t0b; // @[Top.scala 21:12]
  assign n157_I_1_0_t1b = n146_O_1_0_t1b; // @[Top.scala 21:12]
  assign n157_I_1_1_t0b = n146_O_1_1_t0b; // @[Top.scala 21:12]
  assign n157_I_1_1_t1b = n146_O_1_1_t1b; // @[Top.scala 21:12]
  assign n157_I_1_2_t0b = n146_O_1_2_t0b; // @[Top.scala 21:12]
  assign n157_I_1_2_t1b = n146_O_1_2_t1b; // @[Top.scala 21:12]
  assign n157_I_2_0_t0b = n146_O_2_0_t0b; // @[Top.scala 21:12]
  assign n157_I_2_0_t1b = n146_O_2_0_t1b; // @[Top.scala 21:12]
  assign n157_I_2_1_t0b = n146_O_2_1_t0b; // @[Top.scala 21:12]
  assign n157_I_2_1_t1b = n146_O_2_1_t1b; // @[Top.scala 21:12]
  assign n157_I_2_2_t0b = n146_O_2_2_t0b; // @[Top.scala 21:12]
  assign n157_I_2_2_t1b = n146_O_2_2_t1b; // @[Top.scala 21:12]
  assign n162_clock = clock;
  assign n162_valid_up = n157_valid_down; // @[Top.scala 25:19]
  assign n162_I_0_0 = n157_O_0_0; // @[Top.scala 24:12]
  assign n162_I_0_1 = n157_O_0_1; // @[Top.scala 24:12]
  assign n162_I_0_2 = n157_O_0_2; // @[Top.scala 24:12]
  assign n162_I_1_0 = n157_O_1_0; // @[Top.scala 24:12]
  assign n162_I_1_1 = n157_O_1_1; // @[Top.scala 24:12]
  assign n162_I_1_2 = n157_O_1_2; // @[Top.scala 24:12]
  assign n162_I_2_0 = n157_O_2_0; // @[Top.scala 24:12]
  assign n162_I_2_1 = n157_O_2_1; // @[Top.scala 24:12]
  assign n162_I_2_2 = n157_O_2_2; // @[Top.scala 24:12]
  assign n167_clock = clock;
  assign n167_valid_up = n162_valid_down; // @[Top.scala 28:19]
  assign n167_I_0_0 = n162_O_0_0; // @[Top.scala 27:12]
  assign n167_I_1_0 = n162_O_1_0; // @[Top.scala 27:12]
  assign n167_I_2_0 = n162_O_2_0; // @[Top.scala 27:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n170_valid_up = n167_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 33:19]
  assign n170_I0_0_0 = n167_O_0_0; // @[Top.scala 31:13]
  assign n181_valid_up = n170_valid_down; // @[Top.scala 36:19]
  assign n181_I_0_0_t0b = n170_O_0_0_t0b; // @[Top.scala 35:12]
  assign n181_I_0_0_t1b = n170_O_0_0_t1b; // @[Top.scala 35:12]
endmodule
module MapS_12(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_1_1_2,
  input  [7:0] I_1_2_0,
  input  [7:0] I_1_2_1,
  input  [7:0] I_1_2_2,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_0_2,
  input  [7:0] I_2_1_0,
  input  [7:0] I_2_1_1,
  input  [7:0] I_2_1_2,
  input  [7:0] I_2_2_0,
  input  [7:0] I_2_2_1,
  input  [7:0] I_2_2_2,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_0_2,
  input  [7:0] I_3_1_0,
  input  [7:0] I_3_1_1,
  input  [7:0] I_3_1_2,
  input  [7:0] I_3_2_0,
  input  [7:0] I_3_2_1,
  input  [7:0] I_3_2_2,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_0_2,
  input  [7:0] I_4_1_0,
  input  [7:0] I_4_1_1,
  input  [7:0] I_4_1_2,
  input  [7:0] I_4_2_0,
  input  [7:0] I_4_2_1,
  input  [7:0] I_4_2_2,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_0_2,
  input  [7:0] I_5_1_0,
  input  [7:0] I_5_1_1,
  input  [7:0] I_5_1_2,
  input  [7:0] I_5_2_0,
  input  [7:0] I_5_2_1,
  input  [7:0] I_5_2_2,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_0_2,
  input  [7:0] I_6_1_0,
  input  [7:0] I_6_1_1,
  input  [7:0] I_6_1_2,
  input  [7:0] I_6_2_0,
  input  [7:0] I_6_2_1,
  input  [7:0] I_6_2_2,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_0_2,
  input  [7:0] I_7_1_0,
  input  [7:0] I_7_1_1,
  input  [7:0] I_7_1_2,
  input  [7:0] I_7_2_0,
  input  [7:0] I_7_2_1,
  input  [7:0] I_7_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_2_clock; // @[MapS.scala 10:86]
  wire  other_ops_2_reset; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_3_clock; // @[MapS.scala 10:86]
  wire  other_ops_3_reset; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_4_clock; // @[MapS.scala 10:86]
  wire  other_ops_4_reset; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_5_clock; // @[MapS.scala 10:86]
  wire  other_ops_5_reset; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_6_clock; // @[MapS.scala 10:86]
  wire  other_ops_6_reset; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  Module_0 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .I_1_0(fst_op_I_1_0),
    .I_1_1(fst_op_I_1_1),
    .I_1_2(fst_op_I_1_2),
    .I_2_0(fst_op_I_2_0),
    .I_2_1(fst_op_I_2_1),
    .I_2_2(fst_op_I_2_2),
    .O_0_0(fst_op_O_0_0)
  );
  Module_0 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .I_1_0(other_ops_0_I_1_0),
    .I_1_1(other_ops_0_I_1_1),
    .I_1_2(other_ops_0_I_1_2),
    .I_2_0(other_ops_0_I_2_0),
    .I_2_1(other_ops_0_I_2_1),
    .I_2_2(other_ops_0_I_2_2),
    .O_0_0(other_ops_0_O_0_0)
  );
  Module_0 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .I_1_0(other_ops_1_I_1_0),
    .I_1_1(other_ops_1_I_1_1),
    .I_1_2(other_ops_1_I_1_2),
    .I_2_0(other_ops_1_I_2_0),
    .I_2_1(other_ops_1_I_2_1),
    .I_2_2(other_ops_1_I_2_2),
    .O_0_0(other_ops_1_O_0_0)
  );
  Module_0 other_ops_2 ( // @[MapS.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .I_1_0(other_ops_2_I_1_0),
    .I_1_1(other_ops_2_I_1_1),
    .I_1_2(other_ops_2_I_1_2),
    .I_2_0(other_ops_2_I_2_0),
    .I_2_1(other_ops_2_I_2_1),
    .I_2_2(other_ops_2_I_2_2),
    .O_0_0(other_ops_2_O_0_0)
  );
  Module_0 other_ops_3 ( // @[MapS.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_0_2(other_ops_3_I_0_2),
    .I_1_0(other_ops_3_I_1_0),
    .I_1_1(other_ops_3_I_1_1),
    .I_1_2(other_ops_3_I_1_2),
    .I_2_0(other_ops_3_I_2_0),
    .I_2_1(other_ops_3_I_2_1),
    .I_2_2(other_ops_3_I_2_2),
    .O_0_0(other_ops_3_O_0_0)
  );
  Module_0 other_ops_4 ( // @[MapS.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_0_2(other_ops_4_I_0_2),
    .I_1_0(other_ops_4_I_1_0),
    .I_1_1(other_ops_4_I_1_1),
    .I_1_2(other_ops_4_I_1_2),
    .I_2_0(other_ops_4_I_2_0),
    .I_2_1(other_ops_4_I_2_1),
    .I_2_2(other_ops_4_I_2_2),
    .O_0_0(other_ops_4_O_0_0)
  );
  Module_0 other_ops_5 ( // @[MapS.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_0_2(other_ops_5_I_0_2),
    .I_1_0(other_ops_5_I_1_0),
    .I_1_1(other_ops_5_I_1_1),
    .I_1_2(other_ops_5_I_1_2),
    .I_2_0(other_ops_5_I_2_0),
    .I_2_1(other_ops_5_I_2_1),
    .I_2_2(other_ops_5_I_2_2),
    .O_0_0(other_ops_5_O_0_0)
  );
  Module_0 other_ops_6 ( // @[MapS.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_0_2(other_ops_6_I_0_2),
    .I_1_0(other_ops_6_I_1_0),
    .I_1_1(other_ops_6_I_1_1),
    .I_1_2(other_ops_6_I_1_2),
    .I_2_0(other_ops_6_I_2_0),
    .I_2_1(other_ops_6_I_2_1),
    .I_2_2(other_ops_6_I_2_2),
    .O_0_0(other_ops_6_O_0_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_1_0 = I_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_1_1 = I_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_1_2 = I_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_2_0 = I_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_2_1 = I_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_2_2 = I_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_0 = I_1_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_1 = I_1_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_2 = I_1_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_0 = I_1_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_1 = I_1_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_2 = I_1_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_0 = I_2_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_1 = I_2_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_2 = I_2_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_0 = I_2_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_1 = I_2_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_2 = I_2_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_2_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_0 = I_3_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_1 = I_3_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_2 = I_3_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_0 = I_3_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_1 = I_3_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_2 = I_3_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_3_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2 = I_4_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_0 = I_4_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_1 = I_4_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_2 = I_4_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_0 = I_4_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_1 = I_4_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_2 = I_4_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_4_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2 = I_5_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_0 = I_5_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_1 = I_5_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_2 = I_5_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_0 = I_5_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_1 = I_5_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_2 = I_5_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_5_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2 = I_6_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_0 = I_6_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_1 = I_6_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_2 = I_6_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_0 = I_6_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_1 = I_6_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_2 = I_6_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_6_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2 = I_7_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_0 = I_7_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_1 = I_7_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_2 = I_7_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_0 = I_7_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_1 = I_7_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_2 = I_7_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_4(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_1_1_2,
  input  [7:0] I_1_2_0,
  input  [7:0] I_1_2_1,
  input  [7:0] I_1_2_2,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_0_2,
  input  [7:0] I_2_1_0,
  input  [7:0] I_2_1_1,
  input  [7:0] I_2_1_2,
  input  [7:0] I_2_2_0,
  input  [7:0] I_2_2_1,
  input  [7:0] I_2_2_2,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_0_2,
  input  [7:0] I_3_1_0,
  input  [7:0] I_3_1_1,
  input  [7:0] I_3_1_2,
  input  [7:0] I_3_2_0,
  input  [7:0] I_3_2_1,
  input  [7:0] I_3_2_2,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_0_2,
  input  [7:0] I_4_1_0,
  input  [7:0] I_4_1_1,
  input  [7:0] I_4_1_2,
  input  [7:0] I_4_2_0,
  input  [7:0] I_4_2_1,
  input  [7:0] I_4_2_2,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_0_2,
  input  [7:0] I_5_1_0,
  input  [7:0] I_5_1_1,
  input  [7:0] I_5_1_2,
  input  [7:0] I_5_2_0,
  input  [7:0] I_5_2_1,
  input  [7:0] I_5_2_2,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_0_2,
  input  [7:0] I_6_1_0,
  input  [7:0] I_6_1_1,
  input  [7:0] I_6_1_2,
  input  [7:0] I_6_2_0,
  input  [7:0] I_6_2_1,
  input  [7:0] I_6_2_2,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_0_2,
  input  [7:0] I_7_1_0,
  input  [7:0] I_7_1_1,
  input  [7:0] I_7_1_2,
  input  [7:0] I_7_2_0,
  input  [7:0] I_7_2_1,
  input  [7:0] I_7_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[MapT.scala 8:20]
  MapS_12 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_4_1_2(op_I_4_1_2),
    .I_4_2_0(op_I_4_2_0),
    .I_4_2_1(op_I_4_2_1),
    .I_4_2_2(op_I_4_2_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_5_1_2(op_I_5_1_2),
    .I_5_2_0(op_I_5_2_0),
    .I_5_2_1(op_I_5_2_1),
    .I_5_2_2(op_I_5_2_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_6_1_2(op_I_6_1_2),
    .I_6_2_0(op_I_6_2_0),
    .I_6_2_1(op_I_6_2_1),
    .I_6_2_2(op_I_6_2_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_7_1_2(op_I_7_1_2),
    .I_7_2_0(op_I_7_2_0),
    .I_7_2_1(op_I_7_2_1),
    .I_7_2_2(op_I_7_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_1_0_0(op_O_1_0_0),
    .O_2_0_0(op_O_2_0_0),
    .O_3_0_0(op_O_3_0_0),
    .O_4_0_0(op_O_4_0_0),
    .O_5_0_0(op_O_5_0_0),
    .O_6_0_0(op_O_6_0_0),
    .O_7_0_0(op_O_7_0_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_4_1_2 = I_4_1_2; // @[MapT.scala 14:10]
  assign op_I_4_2_0 = I_4_2_0; // @[MapT.scala 14:10]
  assign op_I_4_2_1 = I_4_2_1; // @[MapT.scala 14:10]
  assign op_I_4_2_2 = I_4_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_5_1_2 = I_5_1_2; // @[MapT.scala 14:10]
  assign op_I_5_2_0 = I_5_2_0; // @[MapT.scala 14:10]
  assign op_I_5_2_1 = I_5_2_1; // @[MapT.scala 14:10]
  assign op_I_5_2_2 = I_5_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_6_1_2 = I_6_1_2; // @[MapT.scala 14:10]
  assign op_I_6_2_0 = I_6_2_0; // @[MapT.scala 14:10]
  assign op_I_6_2_1 = I_6_2_1; // @[MapT.scala 14:10]
  assign op_I_6_2_2 = I_6_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_7_1_2 = I_7_1_2; // @[MapT.scala 14:10]
  assign op_I_7_2_0 = I_7_2_0; // @[MapT.scala 14:10]
  assign op_I_7_2_1 = I_7_2_1; // @[MapT.scala 14:10]
  assign op_I_7_2_2 = I_7_2_2; // @[MapT.scala 14:10]
endmodule
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_1_0_0,
  input  [7:0] I_2_0_0,
  input  [7:0] I_3_0_0,
  input  [7:0] I_4_0_0,
  input  [7:0] I_5_0_0,
  input  [7:0] I_6_0_0,
  input  [7:0] I_7_0_0,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0
);
  wire  n1_clock; // @[Top.scala 44:20]
  wire  n1_valid_up; // @[Top.scala 44:20]
  wire  n1_valid_down; // @[Top.scala 44:20]
  wire [7:0] n1_I_0_0_0; // @[Top.scala 44:20]
  wire [7:0] n1_I_1_0_0; // @[Top.scala 44:20]
  wire [7:0] n1_I_2_0_0; // @[Top.scala 44:20]
  wire [7:0] n1_I_3_0_0; // @[Top.scala 44:20]
  wire [7:0] n1_I_4_0_0; // @[Top.scala 44:20]
  wire [7:0] n1_I_5_0_0; // @[Top.scala 44:20]
  wire [7:0] n1_I_6_0_0; // @[Top.scala 44:20]
  wire [7:0] n1_I_7_0_0; // @[Top.scala 44:20]
  wire [7:0] n1_O_0_0_0; // @[Top.scala 44:20]
  wire [7:0] n1_O_1_0_0; // @[Top.scala 44:20]
  wire [7:0] n1_O_2_0_0; // @[Top.scala 44:20]
  wire [7:0] n1_O_3_0_0; // @[Top.scala 44:20]
  wire [7:0] n1_O_4_0_0; // @[Top.scala 44:20]
  wire [7:0] n1_O_5_0_0; // @[Top.scala 44:20]
  wire [7:0] n1_O_6_0_0; // @[Top.scala 44:20]
  wire [7:0] n1_O_7_0_0; // @[Top.scala 44:20]
  wire  n2_clock; // @[Top.scala 47:20]
  wire  n2_reset; // @[Top.scala 47:20]
  wire  n2_valid_up; // @[Top.scala 47:20]
  wire  n2_valid_down; // @[Top.scala 47:20]
  wire [7:0] n2_I_0_0_0; // @[Top.scala 47:20]
  wire [7:0] n2_I_1_0_0; // @[Top.scala 47:20]
  wire [7:0] n2_I_2_0_0; // @[Top.scala 47:20]
  wire [7:0] n2_I_3_0_0; // @[Top.scala 47:20]
  wire [7:0] n2_I_4_0_0; // @[Top.scala 47:20]
  wire [7:0] n2_I_5_0_0; // @[Top.scala 47:20]
  wire [7:0] n2_I_6_0_0; // @[Top.scala 47:20]
  wire [7:0] n2_I_7_0_0; // @[Top.scala 47:20]
  wire [7:0] n2_O_0_0_0; // @[Top.scala 47:20]
  wire [7:0] n2_O_1_0_0; // @[Top.scala 47:20]
  wire [7:0] n2_O_2_0_0; // @[Top.scala 47:20]
  wire [7:0] n2_O_3_0_0; // @[Top.scala 47:20]
  wire [7:0] n2_O_4_0_0; // @[Top.scala 47:20]
  wire [7:0] n2_O_5_0_0; // @[Top.scala 47:20]
  wire [7:0] n2_O_6_0_0; // @[Top.scala 47:20]
  wire [7:0] n2_O_7_0_0; // @[Top.scala 47:20]
  wire  n3_clock; // @[Top.scala 50:20]
  wire  n3_reset; // @[Top.scala 50:20]
  wire  n3_valid_up; // @[Top.scala 50:20]
  wire  n3_valid_down; // @[Top.scala 50:20]
  wire [7:0] n3_I_0_0_0; // @[Top.scala 50:20]
  wire [7:0] n3_I_1_0_0; // @[Top.scala 50:20]
  wire [7:0] n3_I_2_0_0; // @[Top.scala 50:20]
  wire [7:0] n3_I_3_0_0; // @[Top.scala 50:20]
  wire [7:0] n3_I_4_0_0; // @[Top.scala 50:20]
  wire [7:0] n3_I_5_0_0; // @[Top.scala 50:20]
  wire [7:0] n3_I_6_0_0; // @[Top.scala 50:20]
  wire [7:0] n3_I_7_0_0; // @[Top.scala 50:20]
  wire [7:0] n3_O_0_0_0; // @[Top.scala 50:20]
  wire [7:0] n3_O_1_0_0; // @[Top.scala 50:20]
  wire [7:0] n3_O_2_0_0; // @[Top.scala 50:20]
  wire [7:0] n3_O_3_0_0; // @[Top.scala 50:20]
  wire [7:0] n3_O_4_0_0; // @[Top.scala 50:20]
  wire [7:0] n3_O_5_0_0; // @[Top.scala 50:20]
  wire [7:0] n3_O_6_0_0; // @[Top.scala 50:20]
  wire [7:0] n3_O_7_0_0; // @[Top.scala 50:20]
  wire  n4_clock; // @[Top.scala 53:20]
  wire  n4_valid_up; // @[Top.scala 53:20]
  wire  n4_valid_down; // @[Top.scala 53:20]
  wire [7:0] n4_I_0_0_0; // @[Top.scala 53:20]
  wire [7:0] n4_I_1_0_0; // @[Top.scala 53:20]
  wire [7:0] n4_I_2_0_0; // @[Top.scala 53:20]
  wire [7:0] n4_I_3_0_0; // @[Top.scala 53:20]
  wire [7:0] n4_I_4_0_0; // @[Top.scala 53:20]
  wire [7:0] n4_I_5_0_0; // @[Top.scala 53:20]
  wire [7:0] n4_I_6_0_0; // @[Top.scala 53:20]
  wire [7:0] n4_I_7_0_0; // @[Top.scala 53:20]
  wire [7:0] n4_O_0_0_0; // @[Top.scala 53:20]
  wire [7:0] n4_O_1_0_0; // @[Top.scala 53:20]
  wire [7:0] n4_O_2_0_0; // @[Top.scala 53:20]
  wire [7:0] n4_O_3_0_0; // @[Top.scala 53:20]
  wire [7:0] n4_O_4_0_0; // @[Top.scala 53:20]
  wire [7:0] n4_O_5_0_0; // @[Top.scala 53:20]
  wire [7:0] n4_O_6_0_0; // @[Top.scala 53:20]
  wire [7:0] n4_O_7_0_0; // @[Top.scala 53:20]
  wire  n5_clock; // @[Top.scala 56:20]
  wire  n5_valid_up; // @[Top.scala 56:20]
  wire  n5_valid_down; // @[Top.scala 56:20]
  wire [7:0] n5_I_0_0_0; // @[Top.scala 56:20]
  wire [7:0] n5_I_1_0_0; // @[Top.scala 56:20]
  wire [7:0] n5_I_2_0_0; // @[Top.scala 56:20]
  wire [7:0] n5_I_3_0_0; // @[Top.scala 56:20]
  wire [7:0] n5_I_4_0_0; // @[Top.scala 56:20]
  wire [7:0] n5_I_5_0_0; // @[Top.scala 56:20]
  wire [7:0] n5_I_6_0_0; // @[Top.scala 56:20]
  wire [7:0] n5_I_7_0_0; // @[Top.scala 56:20]
  wire [7:0] n5_O_0_0_0; // @[Top.scala 56:20]
  wire [7:0] n5_O_1_0_0; // @[Top.scala 56:20]
  wire [7:0] n5_O_2_0_0; // @[Top.scala 56:20]
  wire [7:0] n5_O_3_0_0; // @[Top.scala 56:20]
  wire [7:0] n5_O_4_0_0; // @[Top.scala 56:20]
  wire [7:0] n5_O_5_0_0; // @[Top.scala 56:20]
  wire [7:0] n5_O_6_0_0; // @[Top.scala 56:20]
  wire [7:0] n5_O_7_0_0; // @[Top.scala 56:20]
  wire  n6_valid_up; // @[Top.scala 59:20]
  wire  n6_valid_down; // @[Top.scala 59:20]
  wire [7:0] n6_I0_0_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_I0_1_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_I0_2_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_I0_3_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_I0_4_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_I0_5_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_I0_6_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_I0_7_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_I1_0_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_I1_1_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_I1_2_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_I1_3_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_I1_4_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_I1_5_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_I1_6_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_I1_7_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_O_0_0_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_O_0_0_0_1; // @[Top.scala 59:20]
  wire [7:0] n6_O_1_0_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_O_1_0_0_1; // @[Top.scala 59:20]
  wire [7:0] n6_O_2_0_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_O_2_0_0_1; // @[Top.scala 59:20]
  wire [7:0] n6_O_3_0_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_O_3_0_0_1; // @[Top.scala 59:20]
  wire [7:0] n6_O_4_0_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_O_4_0_0_1; // @[Top.scala 59:20]
  wire [7:0] n6_O_5_0_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_O_5_0_0_1; // @[Top.scala 59:20]
  wire [7:0] n6_O_6_0_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_O_6_0_0_1; // @[Top.scala 59:20]
  wire [7:0] n6_O_7_0_0_0; // @[Top.scala 59:20]
  wire [7:0] n6_O_7_0_0_1; // @[Top.scala 59:20]
  wire  n19_valid_up; // @[Top.scala 63:21]
  wire  n19_valid_down; // @[Top.scala 63:21]
  wire [7:0] n19_I0_0_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_I0_0_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_I0_1_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_I0_1_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_I0_2_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_I0_2_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_I0_3_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_I0_3_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_I0_4_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_I0_4_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_I0_5_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_I0_5_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_I0_6_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_I0_6_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_I0_7_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_I0_7_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_I1_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_I1_1_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_I1_2_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_I1_3_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_I1_4_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_I1_5_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_I1_6_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_I1_7_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_O_0_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_O_0_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_O_0_0_0_2; // @[Top.scala 63:21]
  wire [7:0] n19_O_1_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_O_1_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_O_1_0_0_2; // @[Top.scala 63:21]
  wire [7:0] n19_O_2_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_O_2_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_O_2_0_0_2; // @[Top.scala 63:21]
  wire [7:0] n19_O_3_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_O_3_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_O_3_0_0_2; // @[Top.scala 63:21]
  wire [7:0] n19_O_4_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_O_4_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_O_4_0_0_2; // @[Top.scala 63:21]
  wire [7:0] n19_O_5_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_O_5_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_O_5_0_0_2; // @[Top.scala 63:21]
  wire [7:0] n19_O_6_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_O_6_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_O_6_0_0_2; // @[Top.scala 63:21]
  wire [7:0] n19_O_7_0_0_0; // @[Top.scala 63:21]
  wire [7:0] n19_O_7_0_0_1; // @[Top.scala 63:21]
  wire [7:0] n19_O_7_0_0_2; // @[Top.scala 63:21]
  wire  n40_valid_up; // @[Top.scala 67:21]
  wire  n40_valid_down; // @[Top.scala 67:21]
  wire [7:0] n40_I_0_0_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_I_0_0_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_I_0_0_0_2; // @[Top.scala 67:21]
  wire [7:0] n40_I_1_0_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_I_1_0_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_I_1_0_0_2; // @[Top.scala 67:21]
  wire [7:0] n40_I_2_0_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_I_2_0_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_I_2_0_0_2; // @[Top.scala 67:21]
  wire [7:0] n40_I_3_0_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_I_3_0_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_I_3_0_0_2; // @[Top.scala 67:21]
  wire [7:0] n40_I_4_0_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_I_4_0_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_I_4_0_0_2; // @[Top.scala 67:21]
  wire [7:0] n40_I_5_0_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_I_5_0_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_I_5_0_0_2; // @[Top.scala 67:21]
  wire [7:0] n40_I_6_0_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_I_6_0_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_I_6_0_0_2; // @[Top.scala 67:21]
  wire [7:0] n40_I_7_0_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_I_7_0_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_I_7_0_0_2; // @[Top.scala 67:21]
  wire [7:0] n40_O_0_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_O_0_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_O_0_0_2; // @[Top.scala 67:21]
  wire [7:0] n40_O_1_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_O_1_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_O_1_0_2; // @[Top.scala 67:21]
  wire [7:0] n40_O_2_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_O_2_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_O_2_0_2; // @[Top.scala 67:21]
  wire [7:0] n40_O_3_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_O_3_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_O_3_0_2; // @[Top.scala 67:21]
  wire [7:0] n40_O_4_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_O_4_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_O_4_0_2; // @[Top.scala 67:21]
  wire [7:0] n40_O_5_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_O_5_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_O_5_0_2; // @[Top.scala 67:21]
  wire [7:0] n40_O_6_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_O_6_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_O_6_0_2; // @[Top.scala 67:21]
  wire [7:0] n40_O_7_0_0; // @[Top.scala 67:21]
  wire [7:0] n40_O_7_0_1; // @[Top.scala 67:21]
  wire [7:0] n40_O_7_0_2; // @[Top.scala 67:21]
  wire  n41_clock; // @[Top.scala 70:21]
  wire  n41_valid_up; // @[Top.scala 70:21]
  wire  n41_valid_down; // @[Top.scala 70:21]
  wire [7:0] n41_I_0_0_0; // @[Top.scala 70:21]
  wire [7:0] n41_I_1_0_0; // @[Top.scala 70:21]
  wire [7:0] n41_I_2_0_0; // @[Top.scala 70:21]
  wire [7:0] n41_I_3_0_0; // @[Top.scala 70:21]
  wire [7:0] n41_I_4_0_0; // @[Top.scala 70:21]
  wire [7:0] n41_I_5_0_0; // @[Top.scala 70:21]
  wire [7:0] n41_I_6_0_0; // @[Top.scala 70:21]
  wire [7:0] n41_I_7_0_0; // @[Top.scala 70:21]
  wire [7:0] n41_O_0_0_0; // @[Top.scala 70:21]
  wire [7:0] n41_O_1_0_0; // @[Top.scala 70:21]
  wire [7:0] n41_O_2_0_0; // @[Top.scala 70:21]
  wire [7:0] n41_O_3_0_0; // @[Top.scala 70:21]
  wire [7:0] n41_O_4_0_0; // @[Top.scala 70:21]
  wire [7:0] n41_O_5_0_0; // @[Top.scala 70:21]
  wire [7:0] n41_O_6_0_0; // @[Top.scala 70:21]
  wire [7:0] n41_O_7_0_0; // @[Top.scala 70:21]
  wire  n42_clock; // @[Top.scala 73:21]
  wire  n42_valid_up; // @[Top.scala 73:21]
  wire  n42_valid_down; // @[Top.scala 73:21]
  wire [7:0] n42_I_0_0_0; // @[Top.scala 73:21]
  wire [7:0] n42_I_1_0_0; // @[Top.scala 73:21]
  wire [7:0] n42_I_2_0_0; // @[Top.scala 73:21]
  wire [7:0] n42_I_3_0_0; // @[Top.scala 73:21]
  wire [7:0] n42_I_4_0_0; // @[Top.scala 73:21]
  wire [7:0] n42_I_5_0_0; // @[Top.scala 73:21]
  wire [7:0] n42_I_6_0_0; // @[Top.scala 73:21]
  wire [7:0] n42_I_7_0_0; // @[Top.scala 73:21]
  wire [7:0] n42_O_0_0_0; // @[Top.scala 73:21]
  wire [7:0] n42_O_1_0_0; // @[Top.scala 73:21]
  wire [7:0] n42_O_2_0_0; // @[Top.scala 73:21]
  wire [7:0] n42_O_3_0_0; // @[Top.scala 73:21]
  wire [7:0] n42_O_4_0_0; // @[Top.scala 73:21]
  wire [7:0] n42_O_5_0_0; // @[Top.scala 73:21]
  wire [7:0] n42_O_6_0_0; // @[Top.scala 73:21]
  wire [7:0] n42_O_7_0_0; // @[Top.scala 73:21]
  wire  n43_valid_up; // @[Top.scala 76:21]
  wire  n43_valid_down; // @[Top.scala 76:21]
  wire [7:0] n43_I0_0_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_I0_1_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_I0_2_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_I0_3_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_I0_4_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_I0_5_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_I0_6_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_I0_7_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_I1_0_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_I1_1_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_I1_2_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_I1_3_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_I1_4_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_I1_5_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_I1_6_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_I1_7_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_O_0_0_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_O_0_0_0_1; // @[Top.scala 76:21]
  wire [7:0] n43_O_1_0_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_O_1_0_0_1; // @[Top.scala 76:21]
  wire [7:0] n43_O_2_0_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_O_2_0_0_1; // @[Top.scala 76:21]
  wire [7:0] n43_O_3_0_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_O_3_0_0_1; // @[Top.scala 76:21]
  wire [7:0] n43_O_4_0_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_O_4_0_0_1; // @[Top.scala 76:21]
  wire [7:0] n43_O_5_0_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_O_5_0_0_1; // @[Top.scala 76:21]
  wire [7:0] n43_O_6_0_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_O_6_0_0_1; // @[Top.scala 76:21]
  wire [7:0] n43_O_7_0_0_0; // @[Top.scala 76:21]
  wire [7:0] n43_O_7_0_0_1; // @[Top.scala 76:21]
  wire  n56_valid_up; // @[Top.scala 80:21]
  wire  n56_valid_down; // @[Top.scala 80:21]
  wire [7:0] n56_I0_0_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_I0_0_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_I0_1_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_I0_1_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_I0_2_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_I0_2_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_I0_3_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_I0_3_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_I0_4_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_I0_4_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_I0_5_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_I0_5_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_I0_6_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_I0_6_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_I0_7_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_I0_7_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_I1_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_I1_1_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_I1_2_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_I1_3_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_I1_4_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_I1_5_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_I1_6_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_I1_7_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_O_0_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_O_0_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_O_0_0_0_2; // @[Top.scala 80:21]
  wire [7:0] n56_O_1_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_O_1_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_O_1_0_0_2; // @[Top.scala 80:21]
  wire [7:0] n56_O_2_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_O_2_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_O_2_0_0_2; // @[Top.scala 80:21]
  wire [7:0] n56_O_3_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_O_3_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_O_3_0_0_2; // @[Top.scala 80:21]
  wire [7:0] n56_O_4_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_O_4_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_O_4_0_0_2; // @[Top.scala 80:21]
  wire [7:0] n56_O_5_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_O_5_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_O_5_0_0_2; // @[Top.scala 80:21]
  wire [7:0] n56_O_6_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_O_6_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_O_6_0_0_2; // @[Top.scala 80:21]
  wire [7:0] n56_O_7_0_0_0; // @[Top.scala 80:21]
  wire [7:0] n56_O_7_0_0_1; // @[Top.scala 80:21]
  wire [7:0] n56_O_7_0_0_2; // @[Top.scala 80:21]
  wire  n77_valid_up; // @[Top.scala 84:21]
  wire  n77_valid_down; // @[Top.scala 84:21]
  wire [7:0] n77_I_0_0_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_I_0_0_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_I_0_0_0_2; // @[Top.scala 84:21]
  wire [7:0] n77_I_1_0_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_I_1_0_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_I_1_0_0_2; // @[Top.scala 84:21]
  wire [7:0] n77_I_2_0_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_I_2_0_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_I_2_0_0_2; // @[Top.scala 84:21]
  wire [7:0] n77_I_3_0_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_I_3_0_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_I_3_0_0_2; // @[Top.scala 84:21]
  wire [7:0] n77_I_4_0_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_I_4_0_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_I_4_0_0_2; // @[Top.scala 84:21]
  wire [7:0] n77_I_5_0_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_I_5_0_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_I_5_0_0_2; // @[Top.scala 84:21]
  wire [7:0] n77_I_6_0_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_I_6_0_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_I_6_0_0_2; // @[Top.scala 84:21]
  wire [7:0] n77_I_7_0_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_I_7_0_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_I_7_0_0_2; // @[Top.scala 84:21]
  wire [7:0] n77_O_0_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_O_0_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_O_0_0_2; // @[Top.scala 84:21]
  wire [7:0] n77_O_1_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_O_1_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_O_1_0_2; // @[Top.scala 84:21]
  wire [7:0] n77_O_2_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_O_2_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_O_2_0_2; // @[Top.scala 84:21]
  wire [7:0] n77_O_3_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_O_3_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_O_3_0_2; // @[Top.scala 84:21]
  wire [7:0] n77_O_4_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_O_4_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_O_4_0_2; // @[Top.scala 84:21]
  wire [7:0] n77_O_5_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_O_5_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_O_5_0_2; // @[Top.scala 84:21]
  wire [7:0] n77_O_6_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_O_6_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_O_6_0_2; // @[Top.scala 84:21]
  wire [7:0] n77_O_7_0_0; // @[Top.scala 84:21]
  wire [7:0] n77_O_7_0_1; // @[Top.scala 84:21]
  wire [7:0] n77_O_7_0_2; // @[Top.scala 84:21]
  wire  n78_valid_up; // @[Top.scala 87:21]
  wire  n78_valid_down; // @[Top.scala 87:21]
  wire [7:0] n78_I0_0_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I0_0_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I0_0_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_I0_1_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I0_1_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I0_1_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_I0_2_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I0_2_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I0_2_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_I0_3_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I0_3_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I0_3_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_I0_4_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I0_4_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I0_4_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_I0_5_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I0_5_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I0_5_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_I0_6_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I0_6_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I0_6_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_I0_7_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I0_7_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I0_7_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_I1_0_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I1_0_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I1_0_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_I1_1_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I1_1_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I1_1_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_I1_2_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I1_2_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I1_2_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_I1_3_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I1_3_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I1_3_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_I1_4_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I1_4_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I1_4_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_I1_5_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I1_5_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I1_5_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_I1_6_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I1_6_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I1_6_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_I1_7_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_I1_7_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_I1_7_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_0_0_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_0_0_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_0_0_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_0_0_1_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_0_0_1_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_0_0_1_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_1_0_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_1_0_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_1_0_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_1_0_1_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_1_0_1_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_1_0_1_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_2_0_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_2_0_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_2_0_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_2_0_1_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_2_0_1_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_2_0_1_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_3_0_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_3_0_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_3_0_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_3_0_1_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_3_0_1_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_3_0_1_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_4_0_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_4_0_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_4_0_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_4_0_1_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_4_0_1_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_4_0_1_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_5_0_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_5_0_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_5_0_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_5_0_1_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_5_0_1_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_5_0_1_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_6_0_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_6_0_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_6_0_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_6_0_1_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_6_0_1_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_6_0_1_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_7_0_0_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_7_0_0_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_7_0_0_2; // @[Top.scala 87:21]
  wire [7:0] n78_O_7_0_1_0; // @[Top.scala 87:21]
  wire [7:0] n78_O_7_0_1_1; // @[Top.scala 87:21]
  wire [7:0] n78_O_7_0_1_2; // @[Top.scala 87:21]
  wire  n88_clock; // @[Top.scala 91:21]
  wire  n88_valid_up; // @[Top.scala 91:21]
  wire  n88_valid_down; // @[Top.scala 91:21]
  wire [7:0] n88_I_0_0_0; // @[Top.scala 91:21]
  wire [7:0] n88_I_1_0_0; // @[Top.scala 91:21]
  wire [7:0] n88_I_2_0_0; // @[Top.scala 91:21]
  wire [7:0] n88_I_3_0_0; // @[Top.scala 91:21]
  wire [7:0] n88_I_4_0_0; // @[Top.scala 91:21]
  wire [7:0] n88_I_5_0_0; // @[Top.scala 91:21]
  wire [7:0] n88_I_6_0_0; // @[Top.scala 91:21]
  wire [7:0] n88_I_7_0_0; // @[Top.scala 91:21]
  wire [7:0] n88_O_0_0_0; // @[Top.scala 91:21]
  wire [7:0] n88_O_1_0_0; // @[Top.scala 91:21]
  wire [7:0] n88_O_2_0_0; // @[Top.scala 91:21]
  wire [7:0] n88_O_3_0_0; // @[Top.scala 91:21]
  wire [7:0] n88_O_4_0_0; // @[Top.scala 91:21]
  wire [7:0] n88_O_5_0_0; // @[Top.scala 91:21]
  wire [7:0] n88_O_6_0_0; // @[Top.scala 91:21]
  wire [7:0] n88_O_7_0_0; // @[Top.scala 91:21]
  wire  n89_clock; // @[Top.scala 94:21]
  wire  n89_valid_up; // @[Top.scala 94:21]
  wire  n89_valid_down; // @[Top.scala 94:21]
  wire [7:0] n89_I_0_0_0; // @[Top.scala 94:21]
  wire [7:0] n89_I_1_0_0; // @[Top.scala 94:21]
  wire [7:0] n89_I_2_0_0; // @[Top.scala 94:21]
  wire [7:0] n89_I_3_0_0; // @[Top.scala 94:21]
  wire [7:0] n89_I_4_0_0; // @[Top.scala 94:21]
  wire [7:0] n89_I_5_0_0; // @[Top.scala 94:21]
  wire [7:0] n89_I_6_0_0; // @[Top.scala 94:21]
  wire [7:0] n89_I_7_0_0; // @[Top.scala 94:21]
  wire [7:0] n89_O_0_0_0; // @[Top.scala 94:21]
  wire [7:0] n89_O_1_0_0; // @[Top.scala 94:21]
  wire [7:0] n89_O_2_0_0; // @[Top.scala 94:21]
  wire [7:0] n89_O_3_0_0; // @[Top.scala 94:21]
  wire [7:0] n89_O_4_0_0; // @[Top.scala 94:21]
  wire [7:0] n89_O_5_0_0; // @[Top.scala 94:21]
  wire [7:0] n89_O_6_0_0; // @[Top.scala 94:21]
  wire [7:0] n89_O_7_0_0; // @[Top.scala 94:21]
  wire  n90_valid_up; // @[Top.scala 97:21]
  wire  n90_valid_down; // @[Top.scala 97:21]
  wire [7:0] n90_I0_0_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_I0_1_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_I0_2_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_I0_3_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_I0_4_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_I0_5_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_I0_6_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_I0_7_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_I1_0_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_I1_1_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_I1_2_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_I1_3_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_I1_4_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_I1_5_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_I1_6_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_I1_7_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_O_0_0_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_O_0_0_0_1; // @[Top.scala 97:21]
  wire [7:0] n90_O_1_0_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_O_1_0_0_1; // @[Top.scala 97:21]
  wire [7:0] n90_O_2_0_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_O_2_0_0_1; // @[Top.scala 97:21]
  wire [7:0] n90_O_3_0_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_O_3_0_0_1; // @[Top.scala 97:21]
  wire [7:0] n90_O_4_0_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_O_4_0_0_1; // @[Top.scala 97:21]
  wire [7:0] n90_O_5_0_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_O_5_0_0_1; // @[Top.scala 97:21]
  wire [7:0] n90_O_6_0_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_O_6_0_0_1; // @[Top.scala 97:21]
  wire [7:0] n90_O_7_0_0_0; // @[Top.scala 97:21]
  wire [7:0] n90_O_7_0_0_1; // @[Top.scala 97:21]
  wire  n103_valid_up; // @[Top.scala 101:22]
  wire  n103_valid_down; // @[Top.scala 101:22]
  wire [7:0] n103_I0_0_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_I0_0_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_I0_1_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_I0_1_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_I0_2_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_I0_2_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_I0_3_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_I0_3_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_I0_4_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_I0_4_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_I0_5_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_I0_5_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_I0_6_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_I0_6_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_I0_7_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_I0_7_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_I1_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_I1_1_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_I1_2_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_I1_3_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_I1_4_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_I1_5_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_I1_6_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_I1_7_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_O_0_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_O_0_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_O_0_0_0_2; // @[Top.scala 101:22]
  wire [7:0] n103_O_1_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_O_1_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_O_1_0_0_2; // @[Top.scala 101:22]
  wire [7:0] n103_O_2_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_O_2_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_O_2_0_0_2; // @[Top.scala 101:22]
  wire [7:0] n103_O_3_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_O_3_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_O_3_0_0_2; // @[Top.scala 101:22]
  wire [7:0] n103_O_4_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_O_4_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_O_4_0_0_2; // @[Top.scala 101:22]
  wire [7:0] n103_O_5_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_O_5_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_O_5_0_0_2; // @[Top.scala 101:22]
  wire [7:0] n103_O_6_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_O_6_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_O_6_0_0_2; // @[Top.scala 101:22]
  wire [7:0] n103_O_7_0_0_0; // @[Top.scala 101:22]
  wire [7:0] n103_O_7_0_0_1; // @[Top.scala 101:22]
  wire [7:0] n103_O_7_0_0_2; // @[Top.scala 101:22]
  wire  n124_valid_up; // @[Top.scala 105:22]
  wire  n124_valid_down; // @[Top.scala 105:22]
  wire [7:0] n124_I_0_0_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_I_0_0_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_I_0_0_0_2; // @[Top.scala 105:22]
  wire [7:0] n124_I_1_0_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_I_1_0_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_I_1_0_0_2; // @[Top.scala 105:22]
  wire [7:0] n124_I_2_0_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_I_2_0_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_I_2_0_0_2; // @[Top.scala 105:22]
  wire [7:0] n124_I_3_0_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_I_3_0_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_I_3_0_0_2; // @[Top.scala 105:22]
  wire [7:0] n124_I_4_0_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_I_4_0_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_I_4_0_0_2; // @[Top.scala 105:22]
  wire [7:0] n124_I_5_0_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_I_5_0_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_I_5_0_0_2; // @[Top.scala 105:22]
  wire [7:0] n124_I_6_0_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_I_6_0_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_I_6_0_0_2; // @[Top.scala 105:22]
  wire [7:0] n124_I_7_0_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_I_7_0_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_I_7_0_0_2; // @[Top.scala 105:22]
  wire [7:0] n124_O_0_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_O_0_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_O_0_0_2; // @[Top.scala 105:22]
  wire [7:0] n124_O_1_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_O_1_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_O_1_0_2; // @[Top.scala 105:22]
  wire [7:0] n124_O_2_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_O_2_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_O_2_0_2; // @[Top.scala 105:22]
  wire [7:0] n124_O_3_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_O_3_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_O_3_0_2; // @[Top.scala 105:22]
  wire [7:0] n124_O_4_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_O_4_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_O_4_0_2; // @[Top.scala 105:22]
  wire [7:0] n124_O_5_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_O_5_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_O_5_0_2; // @[Top.scala 105:22]
  wire [7:0] n124_O_6_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_O_6_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_O_6_0_2; // @[Top.scala 105:22]
  wire [7:0] n124_O_7_0_0; // @[Top.scala 105:22]
  wire [7:0] n124_O_7_0_1; // @[Top.scala 105:22]
  wire [7:0] n124_O_7_0_2; // @[Top.scala 105:22]
  wire  n125_valid_up; // @[Top.scala 108:22]
  wire  n125_valid_down; // @[Top.scala 108:22]
  wire [7:0] n125_I0_0_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_0_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_0_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_I0_0_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_0_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_0_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_I0_1_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_1_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_1_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_I0_1_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_1_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_1_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_I0_2_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_2_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_2_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_I0_2_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_2_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_2_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_I0_3_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_3_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_3_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_I0_3_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_3_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_3_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_I0_4_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_4_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_4_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_I0_4_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_4_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_4_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_I0_5_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_5_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_5_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_I0_5_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_5_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_5_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_I0_6_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_6_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_6_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_I0_6_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_6_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_6_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_I0_7_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_7_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_7_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_I0_7_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_I0_7_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_I0_7_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_I1_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I1_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I1_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_I1_1_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I1_1_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I1_1_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_I1_2_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I1_2_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I1_2_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_I1_3_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I1_3_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I1_3_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_I1_4_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I1_4_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I1_4_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_I1_5_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I1_5_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I1_5_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_I1_6_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I1_6_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I1_6_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_I1_7_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_I1_7_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_I1_7_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_0_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_0_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_0_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_0_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_0_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_0_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_0_0_2_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_0_0_2_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_0_0_2_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_1_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_1_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_1_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_1_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_1_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_1_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_1_0_2_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_1_0_2_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_1_0_2_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_2_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_2_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_2_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_2_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_2_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_2_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_2_0_2_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_2_0_2_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_2_0_2_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_3_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_3_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_3_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_3_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_3_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_3_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_3_0_2_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_3_0_2_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_3_0_2_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_4_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_4_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_4_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_4_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_4_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_4_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_4_0_2_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_4_0_2_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_4_0_2_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_5_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_5_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_5_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_5_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_5_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_5_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_5_0_2_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_5_0_2_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_5_0_2_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_6_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_6_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_6_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_6_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_6_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_6_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_6_0_2_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_6_0_2_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_6_0_2_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_7_0_0_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_7_0_0_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_7_0_0_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_7_0_1_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_7_0_1_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_7_0_1_2; // @[Top.scala 108:22]
  wire [7:0] n125_O_7_0_2_0; // @[Top.scala 108:22]
  wire [7:0] n125_O_7_0_2_1; // @[Top.scala 108:22]
  wire [7:0] n125_O_7_0_2_2; // @[Top.scala 108:22]
  wire  n141_valid_up; // @[Top.scala 112:22]
  wire  n141_valid_down; // @[Top.scala 112:22]
  wire [7:0] n141_I_0_0_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_0_0_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_0_0_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_0_0_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_0_0_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_0_0_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_0_0_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_0_0_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_0_0_2_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_1_0_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_1_0_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_1_0_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_1_0_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_1_0_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_1_0_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_1_0_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_1_0_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_1_0_2_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_2_0_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_2_0_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_2_0_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_2_0_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_2_0_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_2_0_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_2_0_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_2_0_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_2_0_2_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_3_0_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_3_0_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_3_0_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_3_0_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_3_0_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_3_0_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_3_0_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_3_0_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_3_0_2_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_4_0_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_4_0_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_4_0_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_4_0_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_4_0_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_4_0_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_4_0_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_4_0_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_4_0_2_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_5_0_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_5_0_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_5_0_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_5_0_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_5_0_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_5_0_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_5_0_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_5_0_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_5_0_2_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_6_0_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_6_0_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_6_0_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_6_0_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_6_0_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_6_0_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_6_0_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_6_0_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_6_0_2_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_7_0_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_7_0_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_7_0_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_7_0_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_7_0_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_7_0_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_I_7_0_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_I_7_0_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_I_7_0_2_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_0_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_0_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_0_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_0_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_0_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_0_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_0_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_0_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_0_2_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_1_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_1_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_1_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_1_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_1_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_1_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_1_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_1_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_1_2_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_2_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_2_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_2_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_2_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_2_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_2_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_2_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_2_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_2_2_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_3_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_3_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_3_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_3_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_3_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_3_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_3_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_3_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_3_2_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_4_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_4_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_4_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_4_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_4_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_4_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_4_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_4_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_4_2_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_5_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_5_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_5_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_5_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_5_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_5_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_5_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_5_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_5_2_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_6_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_6_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_6_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_6_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_6_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_6_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_6_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_6_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_6_2_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_7_0_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_7_0_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_7_0_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_7_1_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_7_1_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_7_1_2; // @[Top.scala 112:22]
  wire [7:0] n141_O_7_2_0; // @[Top.scala 112:22]
  wire [7:0] n141_O_7_2_1; // @[Top.scala 112:22]
  wire [7:0] n141_O_7_2_2; // @[Top.scala 112:22]
  wire  n183_clock; // @[Top.scala 115:22]
  wire  n183_reset; // @[Top.scala 115:22]
  wire  n183_valid_up; // @[Top.scala 115:22]
  wire  n183_valid_down; // @[Top.scala 115:22]
  wire [7:0] n183_I_0_0_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_0_0_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_0_0_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_0_1_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_0_1_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_0_1_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_0_2_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_0_2_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_0_2_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_1_0_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_1_0_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_1_0_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_1_1_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_1_1_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_1_1_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_1_2_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_1_2_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_1_2_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_2_0_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_2_0_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_2_0_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_2_1_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_2_1_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_2_1_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_2_2_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_2_2_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_2_2_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_3_0_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_3_0_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_3_0_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_3_1_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_3_1_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_3_1_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_3_2_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_3_2_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_3_2_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_4_0_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_4_0_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_4_0_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_4_1_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_4_1_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_4_1_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_4_2_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_4_2_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_4_2_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_5_0_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_5_0_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_5_0_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_5_1_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_5_1_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_5_1_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_5_2_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_5_2_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_5_2_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_6_0_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_6_0_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_6_0_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_6_1_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_6_1_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_6_1_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_6_2_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_6_2_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_6_2_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_7_0_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_7_0_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_7_0_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_7_1_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_7_1_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_7_1_2; // @[Top.scala 115:22]
  wire [7:0] n183_I_7_2_0; // @[Top.scala 115:22]
  wire [7:0] n183_I_7_2_1; // @[Top.scala 115:22]
  wire [7:0] n183_I_7_2_2; // @[Top.scala 115:22]
  wire [7:0] n183_O_0_0_0; // @[Top.scala 115:22]
  wire [7:0] n183_O_1_0_0; // @[Top.scala 115:22]
  wire [7:0] n183_O_2_0_0; // @[Top.scala 115:22]
  wire [7:0] n183_O_3_0_0; // @[Top.scala 115:22]
  wire [7:0] n183_O_4_0_0; // @[Top.scala 115:22]
  wire [7:0] n183_O_5_0_0; // @[Top.scala 115:22]
  wire [7:0] n183_O_6_0_0; // @[Top.scala 115:22]
  wire [7:0] n183_O_7_0_0; // @[Top.scala 115:22]
  wire  n184_clock; // @[Top.scala 118:22]
  wire  n184_valid_up; // @[Top.scala 118:22]
  wire  n184_valid_down; // @[Top.scala 118:22]
  wire [7:0] n184_I_0_0_0; // @[Top.scala 118:22]
  wire [7:0] n184_I_1_0_0; // @[Top.scala 118:22]
  wire [7:0] n184_I_2_0_0; // @[Top.scala 118:22]
  wire [7:0] n184_I_3_0_0; // @[Top.scala 118:22]
  wire [7:0] n184_I_4_0_0; // @[Top.scala 118:22]
  wire [7:0] n184_I_5_0_0; // @[Top.scala 118:22]
  wire [7:0] n184_I_6_0_0; // @[Top.scala 118:22]
  wire [7:0] n184_I_7_0_0; // @[Top.scala 118:22]
  wire [7:0] n184_O_0_0_0; // @[Top.scala 118:22]
  wire [7:0] n184_O_1_0_0; // @[Top.scala 118:22]
  wire [7:0] n184_O_2_0_0; // @[Top.scala 118:22]
  wire [7:0] n184_O_3_0_0; // @[Top.scala 118:22]
  wire [7:0] n184_O_4_0_0; // @[Top.scala 118:22]
  wire [7:0] n184_O_5_0_0; // @[Top.scala 118:22]
  wire [7:0] n184_O_6_0_0; // @[Top.scala 118:22]
  wire [7:0] n184_O_7_0_0; // @[Top.scala 118:22]
  wire  n185_clock; // @[Top.scala 121:22]
  wire  n185_valid_up; // @[Top.scala 121:22]
  wire  n185_valid_down; // @[Top.scala 121:22]
  wire [7:0] n185_I_0_0_0; // @[Top.scala 121:22]
  wire [7:0] n185_I_1_0_0; // @[Top.scala 121:22]
  wire [7:0] n185_I_2_0_0; // @[Top.scala 121:22]
  wire [7:0] n185_I_3_0_0; // @[Top.scala 121:22]
  wire [7:0] n185_I_4_0_0; // @[Top.scala 121:22]
  wire [7:0] n185_I_5_0_0; // @[Top.scala 121:22]
  wire [7:0] n185_I_6_0_0; // @[Top.scala 121:22]
  wire [7:0] n185_I_7_0_0; // @[Top.scala 121:22]
  wire [7:0] n185_O_0_0_0; // @[Top.scala 121:22]
  wire [7:0] n185_O_1_0_0; // @[Top.scala 121:22]
  wire [7:0] n185_O_2_0_0; // @[Top.scala 121:22]
  wire [7:0] n185_O_3_0_0; // @[Top.scala 121:22]
  wire [7:0] n185_O_4_0_0; // @[Top.scala 121:22]
  wire [7:0] n185_O_5_0_0; // @[Top.scala 121:22]
  wire [7:0] n185_O_6_0_0; // @[Top.scala 121:22]
  wire [7:0] n185_O_7_0_0; // @[Top.scala 121:22]
  wire  n186_clock; // @[Top.scala 124:22]
  wire  n186_valid_up; // @[Top.scala 124:22]
  wire  n186_valid_down; // @[Top.scala 124:22]
  wire [7:0] n186_I_0_0_0; // @[Top.scala 124:22]
  wire [7:0] n186_I_1_0_0; // @[Top.scala 124:22]
  wire [7:0] n186_I_2_0_0; // @[Top.scala 124:22]
  wire [7:0] n186_I_3_0_0; // @[Top.scala 124:22]
  wire [7:0] n186_I_4_0_0; // @[Top.scala 124:22]
  wire [7:0] n186_I_5_0_0; // @[Top.scala 124:22]
  wire [7:0] n186_I_6_0_0; // @[Top.scala 124:22]
  wire [7:0] n186_I_7_0_0; // @[Top.scala 124:22]
  wire [7:0] n186_O_0_0_0; // @[Top.scala 124:22]
  wire [7:0] n186_O_1_0_0; // @[Top.scala 124:22]
  wire [7:0] n186_O_2_0_0; // @[Top.scala 124:22]
  wire [7:0] n186_O_3_0_0; // @[Top.scala 124:22]
  wire [7:0] n186_O_4_0_0; // @[Top.scala 124:22]
  wire [7:0] n186_O_5_0_0; // @[Top.scala 124:22]
  wire [7:0] n186_O_6_0_0; // @[Top.scala 124:22]
  wire [7:0] n186_O_7_0_0; // @[Top.scala 124:22]
  FIFO n1 ( // @[Top.scala 44:20]
    .clock(n1_clock),
    .valid_up(n1_valid_up),
    .valid_down(n1_valid_down),
    .I_0_0_0(n1_I_0_0_0),
    .I_1_0_0(n1_I_1_0_0),
    .I_2_0_0(n1_I_2_0_0),
    .I_3_0_0(n1_I_3_0_0),
    .I_4_0_0(n1_I_4_0_0),
    .I_5_0_0(n1_I_5_0_0),
    .I_6_0_0(n1_I_6_0_0),
    .I_7_0_0(n1_I_7_0_0),
    .O_0_0_0(n1_O_0_0_0),
    .O_1_0_0(n1_O_1_0_0),
    .O_2_0_0(n1_O_2_0_0),
    .O_3_0_0(n1_O_3_0_0),
    .O_4_0_0(n1_O_4_0_0),
    .O_5_0_0(n1_O_5_0_0),
    .O_6_0_0(n1_O_6_0_0),
    .O_7_0_0(n1_O_7_0_0)
  );
  ShiftTS n2 ( // @[Top.scala 47:20]
    .clock(n2_clock),
    .reset(n2_reset),
    .valid_up(n2_valid_up),
    .valid_down(n2_valid_down),
    .I_0_0_0(n2_I_0_0_0),
    .I_1_0_0(n2_I_1_0_0),
    .I_2_0_0(n2_I_2_0_0),
    .I_3_0_0(n2_I_3_0_0),
    .I_4_0_0(n2_I_4_0_0),
    .I_5_0_0(n2_I_5_0_0),
    .I_6_0_0(n2_I_6_0_0),
    .I_7_0_0(n2_I_7_0_0),
    .O_0_0_0(n2_O_0_0_0),
    .O_1_0_0(n2_O_1_0_0),
    .O_2_0_0(n2_O_2_0_0),
    .O_3_0_0(n2_O_3_0_0),
    .O_4_0_0(n2_O_4_0_0),
    .O_5_0_0(n2_O_5_0_0),
    .O_6_0_0(n2_O_6_0_0),
    .O_7_0_0(n2_O_7_0_0)
  );
  ShiftTS n3 ( // @[Top.scala 50:20]
    .clock(n3_clock),
    .reset(n3_reset),
    .valid_up(n3_valid_up),
    .valid_down(n3_valid_down),
    .I_0_0_0(n3_I_0_0_0),
    .I_1_0_0(n3_I_1_0_0),
    .I_2_0_0(n3_I_2_0_0),
    .I_3_0_0(n3_I_3_0_0),
    .I_4_0_0(n3_I_4_0_0),
    .I_5_0_0(n3_I_5_0_0),
    .I_6_0_0(n3_I_6_0_0),
    .I_7_0_0(n3_I_7_0_0),
    .O_0_0_0(n3_O_0_0_0),
    .O_1_0_0(n3_O_1_0_0),
    .O_2_0_0(n3_O_2_0_0),
    .O_3_0_0(n3_O_3_0_0),
    .O_4_0_0(n3_O_4_0_0),
    .O_5_0_0(n3_O_5_0_0),
    .O_6_0_0(n3_O_6_0_0),
    .O_7_0_0(n3_O_7_0_0)
  );
  ShiftTS_2 n4 ( // @[Top.scala 53:20]
    .clock(n4_clock),
    .valid_up(n4_valid_up),
    .valid_down(n4_valid_down),
    .I_0_0_0(n4_I_0_0_0),
    .I_1_0_0(n4_I_1_0_0),
    .I_2_0_0(n4_I_2_0_0),
    .I_3_0_0(n4_I_3_0_0),
    .I_4_0_0(n4_I_4_0_0),
    .I_5_0_0(n4_I_5_0_0),
    .I_6_0_0(n4_I_6_0_0),
    .I_7_0_0(n4_I_7_0_0),
    .O_0_0_0(n4_O_0_0_0),
    .O_1_0_0(n4_O_1_0_0),
    .O_2_0_0(n4_O_2_0_0),
    .O_3_0_0(n4_O_3_0_0),
    .O_4_0_0(n4_O_4_0_0),
    .O_5_0_0(n4_O_5_0_0),
    .O_6_0_0(n4_O_6_0_0),
    .O_7_0_0(n4_O_7_0_0)
  );
  ShiftTS_2 n5 ( // @[Top.scala 56:20]
    .clock(n5_clock),
    .valid_up(n5_valid_up),
    .valid_down(n5_valid_down),
    .I_0_0_0(n5_I_0_0_0),
    .I_1_0_0(n5_I_1_0_0),
    .I_2_0_0(n5_I_2_0_0),
    .I_3_0_0(n5_I_3_0_0),
    .I_4_0_0(n5_I_4_0_0),
    .I_5_0_0(n5_I_5_0_0),
    .I_6_0_0(n5_I_6_0_0),
    .I_7_0_0(n5_I_7_0_0),
    .O_0_0_0(n5_O_0_0_0),
    .O_1_0_0(n5_O_1_0_0),
    .O_2_0_0(n5_O_2_0_0),
    .O_3_0_0(n5_O_3_0_0),
    .O_4_0_0(n5_O_4_0_0),
    .O_5_0_0(n5_O_5_0_0),
    .O_6_0_0(n5_O_6_0_0),
    .O_7_0_0(n5_O_7_0_0)
  );
  Map2T n6 ( // @[Top.scala 59:20]
    .valid_up(n6_valid_up),
    .valid_down(n6_valid_down),
    .I0_0_0_0(n6_I0_0_0_0),
    .I0_1_0_0(n6_I0_1_0_0),
    .I0_2_0_0(n6_I0_2_0_0),
    .I0_3_0_0(n6_I0_3_0_0),
    .I0_4_0_0(n6_I0_4_0_0),
    .I0_5_0_0(n6_I0_5_0_0),
    .I0_6_0_0(n6_I0_6_0_0),
    .I0_7_0_0(n6_I0_7_0_0),
    .I1_0_0_0(n6_I1_0_0_0),
    .I1_1_0_0(n6_I1_1_0_0),
    .I1_2_0_0(n6_I1_2_0_0),
    .I1_3_0_0(n6_I1_3_0_0),
    .I1_4_0_0(n6_I1_4_0_0),
    .I1_5_0_0(n6_I1_5_0_0),
    .I1_6_0_0(n6_I1_6_0_0),
    .I1_7_0_0(n6_I1_7_0_0),
    .O_0_0_0_0(n6_O_0_0_0_0),
    .O_0_0_0_1(n6_O_0_0_0_1),
    .O_1_0_0_0(n6_O_1_0_0_0),
    .O_1_0_0_1(n6_O_1_0_0_1),
    .O_2_0_0_0(n6_O_2_0_0_0),
    .O_2_0_0_1(n6_O_2_0_0_1),
    .O_3_0_0_0(n6_O_3_0_0_0),
    .O_3_0_0_1(n6_O_3_0_0_1),
    .O_4_0_0_0(n6_O_4_0_0_0),
    .O_4_0_0_1(n6_O_4_0_0_1),
    .O_5_0_0_0(n6_O_5_0_0_0),
    .O_5_0_0_1(n6_O_5_0_0_1),
    .O_6_0_0_0(n6_O_6_0_0_0),
    .O_6_0_0_1(n6_O_6_0_0_1),
    .O_7_0_0_0(n6_O_7_0_0_0),
    .O_7_0_0_1(n6_O_7_0_0_1)
  );
  Map2T_1 n19 ( // @[Top.scala 63:21]
    .valid_up(n19_valid_up),
    .valid_down(n19_valid_down),
    .I0_0_0_0_0(n19_I0_0_0_0_0),
    .I0_0_0_0_1(n19_I0_0_0_0_1),
    .I0_1_0_0_0(n19_I0_1_0_0_0),
    .I0_1_0_0_1(n19_I0_1_0_0_1),
    .I0_2_0_0_0(n19_I0_2_0_0_0),
    .I0_2_0_0_1(n19_I0_2_0_0_1),
    .I0_3_0_0_0(n19_I0_3_0_0_0),
    .I0_3_0_0_1(n19_I0_3_0_0_1),
    .I0_4_0_0_0(n19_I0_4_0_0_0),
    .I0_4_0_0_1(n19_I0_4_0_0_1),
    .I0_5_0_0_0(n19_I0_5_0_0_0),
    .I0_5_0_0_1(n19_I0_5_0_0_1),
    .I0_6_0_0_0(n19_I0_6_0_0_0),
    .I0_6_0_0_1(n19_I0_6_0_0_1),
    .I0_7_0_0_0(n19_I0_7_0_0_0),
    .I0_7_0_0_1(n19_I0_7_0_0_1),
    .I1_0_0_0(n19_I1_0_0_0),
    .I1_1_0_0(n19_I1_1_0_0),
    .I1_2_0_0(n19_I1_2_0_0),
    .I1_3_0_0(n19_I1_3_0_0),
    .I1_4_0_0(n19_I1_4_0_0),
    .I1_5_0_0(n19_I1_5_0_0),
    .I1_6_0_0(n19_I1_6_0_0),
    .I1_7_0_0(n19_I1_7_0_0),
    .O_0_0_0_0(n19_O_0_0_0_0),
    .O_0_0_0_1(n19_O_0_0_0_1),
    .O_0_0_0_2(n19_O_0_0_0_2),
    .O_1_0_0_0(n19_O_1_0_0_0),
    .O_1_0_0_1(n19_O_1_0_0_1),
    .O_1_0_0_2(n19_O_1_0_0_2),
    .O_2_0_0_0(n19_O_2_0_0_0),
    .O_2_0_0_1(n19_O_2_0_0_1),
    .O_2_0_0_2(n19_O_2_0_0_2),
    .O_3_0_0_0(n19_O_3_0_0_0),
    .O_3_0_0_1(n19_O_3_0_0_1),
    .O_3_0_0_2(n19_O_3_0_0_2),
    .O_4_0_0_0(n19_O_4_0_0_0),
    .O_4_0_0_1(n19_O_4_0_0_1),
    .O_4_0_0_2(n19_O_4_0_0_2),
    .O_5_0_0_0(n19_O_5_0_0_0),
    .O_5_0_0_1(n19_O_5_0_0_1),
    .O_5_0_0_2(n19_O_5_0_0_2),
    .O_6_0_0_0(n19_O_6_0_0_0),
    .O_6_0_0_1(n19_O_6_0_0_1),
    .O_6_0_0_2(n19_O_6_0_0_2),
    .O_7_0_0_0(n19_O_7_0_0_0),
    .O_7_0_0_1(n19_O_7_0_0_1),
    .O_7_0_0_2(n19_O_7_0_0_2)
  );
  MapT n40 ( // @[Top.scala 67:21]
    .valid_up(n40_valid_up),
    .valid_down(n40_valid_down),
    .I_0_0_0_0(n40_I_0_0_0_0),
    .I_0_0_0_1(n40_I_0_0_0_1),
    .I_0_0_0_2(n40_I_0_0_0_2),
    .I_1_0_0_0(n40_I_1_0_0_0),
    .I_1_0_0_1(n40_I_1_0_0_1),
    .I_1_0_0_2(n40_I_1_0_0_2),
    .I_2_0_0_0(n40_I_2_0_0_0),
    .I_2_0_0_1(n40_I_2_0_0_1),
    .I_2_0_0_2(n40_I_2_0_0_2),
    .I_3_0_0_0(n40_I_3_0_0_0),
    .I_3_0_0_1(n40_I_3_0_0_1),
    .I_3_0_0_2(n40_I_3_0_0_2),
    .I_4_0_0_0(n40_I_4_0_0_0),
    .I_4_0_0_1(n40_I_4_0_0_1),
    .I_4_0_0_2(n40_I_4_0_0_2),
    .I_5_0_0_0(n40_I_5_0_0_0),
    .I_5_0_0_1(n40_I_5_0_0_1),
    .I_5_0_0_2(n40_I_5_0_0_2),
    .I_6_0_0_0(n40_I_6_0_0_0),
    .I_6_0_0_1(n40_I_6_0_0_1),
    .I_6_0_0_2(n40_I_6_0_0_2),
    .I_7_0_0_0(n40_I_7_0_0_0),
    .I_7_0_0_1(n40_I_7_0_0_1),
    .I_7_0_0_2(n40_I_7_0_0_2),
    .O_0_0_0(n40_O_0_0_0),
    .O_0_0_1(n40_O_0_0_1),
    .O_0_0_2(n40_O_0_0_2),
    .O_1_0_0(n40_O_1_0_0),
    .O_1_0_1(n40_O_1_0_1),
    .O_1_0_2(n40_O_1_0_2),
    .O_2_0_0(n40_O_2_0_0),
    .O_2_0_1(n40_O_2_0_1),
    .O_2_0_2(n40_O_2_0_2),
    .O_3_0_0(n40_O_3_0_0),
    .O_3_0_1(n40_O_3_0_1),
    .O_3_0_2(n40_O_3_0_2),
    .O_4_0_0(n40_O_4_0_0),
    .O_4_0_1(n40_O_4_0_1),
    .O_4_0_2(n40_O_4_0_2),
    .O_5_0_0(n40_O_5_0_0),
    .O_5_0_1(n40_O_5_0_1),
    .O_5_0_2(n40_O_5_0_2),
    .O_6_0_0(n40_O_6_0_0),
    .O_6_0_1(n40_O_6_0_1),
    .O_6_0_2(n40_O_6_0_2),
    .O_7_0_0(n40_O_7_0_0),
    .O_7_0_1(n40_O_7_0_1),
    .O_7_0_2(n40_O_7_0_2)
  );
  ShiftTS_2 n41 ( // @[Top.scala 70:21]
    .clock(n41_clock),
    .valid_up(n41_valid_up),
    .valid_down(n41_valid_down),
    .I_0_0_0(n41_I_0_0_0),
    .I_1_0_0(n41_I_1_0_0),
    .I_2_0_0(n41_I_2_0_0),
    .I_3_0_0(n41_I_3_0_0),
    .I_4_0_0(n41_I_4_0_0),
    .I_5_0_0(n41_I_5_0_0),
    .I_6_0_0(n41_I_6_0_0),
    .I_7_0_0(n41_I_7_0_0),
    .O_0_0_0(n41_O_0_0_0),
    .O_1_0_0(n41_O_1_0_0),
    .O_2_0_0(n41_O_2_0_0),
    .O_3_0_0(n41_O_3_0_0),
    .O_4_0_0(n41_O_4_0_0),
    .O_5_0_0(n41_O_5_0_0),
    .O_6_0_0(n41_O_6_0_0),
    .O_7_0_0(n41_O_7_0_0)
  );
  ShiftTS_2 n42 ( // @[Top.scala 73:21]
    .clock(n42_clock),
    .valid_up(n42_valid_up),
    .valid_down(n42_valid_down),
    .I_0_0_0(n42_I_0_0_0),
    .I_1_0_0(n42_I_1_0_0),
    .I_2_0_0(n42_I_2_0_0),
    .I_3_0_0(n42_I_3_0_0),
    .I_4_0_0(n42_I_4_0_0),
    .I_5_0_0(n42_I_5_0_0),
    .I_6_0_0(n42_I_6_0_0),
    .I_7_0_0(n42_I_7_0_0),
    .O_0_0_0(n42_O_0_0_0),
    .O_1_0_0(n42_O_1_0_0),
    .O_2_0_0(n42_O_2_0_0),
    .O_3_0_0(n42_O_3_0_0),
    .O_4_0_0(n42_O_4_0_0),
    .O_5_0_0(n42_O_5_0_0),
    .O_6_0_0(n42_O_6_0_0),
    .O_7_0_0(n42_O_7_0_0)
  );
  Map2T n43 ( // @[Top.scala 76:21]
    .valid_up(n43_valid_up),
    .valid_down(n43_valid_down),
    .I0_0_0_0(n43_I0_0_0_0),
    .I0_1_0_0(n43_I0_1_0_0),
    .I0_2_0_0(n43_I0_2_0_0),
    .I0_3_0_0(n43_I0_3_0_0),
    .I0_4_0_0(n43_I0_4_0_0),
    .I0_5_0_0(n43_I0_5_0_0),
    .I0_6_0_0(n43_I0_6_0_0),
    .I0_7_0_0(n43_I0_7_0_0),
    .I1_0_0_0(n43_I1_0_0_0),
    .I1_1_0_0(n43_I1_1_0_0),
    .I1_2_0_0(n43_I1_2_0_0),
    .I1_3_0_0(n43_I1_3_0_0),
    .I1_4_0_0(n43_I1_4_0_0),
    .I1_5_0_0(n43_I1_5_0_0),
    .I1_6_0_0(n43_I1_6_0_0),
    .I1_7_0_0(n43_I1_7_0_0),
    .O_0_0_0_0(n43_O_0_0_0_0),
    .O_0_0_0_1(n43_O_0_0_0_1),
    .O_1_0_0_0(n43_O_1_0_0_0),
    .O_1_0_0_1(n43_O_1_0_0_1),
    .O_2_0_0_0(n43_O_2_0_0_0),
    .O_2_0_0_1(n43_O_2_0_0_1),
    .O_3_0_0_0(n43_O_3_0_0_0),
    .O_3_0_0_1(n43_O_3_0_0_1),
    .O_4_0_0_0(n43_O_4_0_0_0),
    .O_4_0_0_1(n43_O_4_0_0_1),
    .O_5_0_0_0(n43_O_5_0_0_0),
    .O_5_0_0_1(n43_O_5_0_0_1),
    .O_6_0_0_0(n43_O_6_0_0_0),
    .O_6_0_0_1(n43_O_6_0_0_1),
    .O_7_0_0_0(n43_O_7_0_0_0),
    .O_7_0_0_1(n43_O_7_0_0_1)
  );
  Map2T_1 n56 ( // @[Top.scala 80:21]
    .valid_up(n56_valid_up),
    .valid_down(n56_valid_down),
    .I0_0_0_0_0(n56_I0_0_0_0_0),
    .I0_0_0_0_1(n56_I0_0_0_0_1),
    .I0_1_0_0_0(n56_I0_1_0_0_0),
    .I0_1_0_0_1(n56_I0_1_0_0_1),
    .I0_2_0_0_0(n56_I0_2_0_0_0),
    .I0_2_0_0_1(n56_I0_2_0_0_1),
    .I0_3_0_0_0(n56_I0_3_0_0_0),
    .I0_3_0_0_1(n56_I0_3_0_0_1),
    .I0_4_0_0_0(n56_I0_4_0_0_0),
    .I0_4_0_0_1(n56_I0_4_0_0_1),
    .I0_5_0_0_0(n56_I0_5_0_0_0),
    .I0_5_0_0_1(n56_I0_5_0_0_1),
    .I0_6_0_0_0(n56_I0_6_0_0_0),
    .I0_6_0_0_1(n56_I0_6_0_0_1),
    .I0_7_0_0_0(n56_I0_7_0_0_0),
    .I0_7_0_0_1(n56_I0_7_0_0_1),
    .I1_0_0_0(n56_I1_0_0_0),
    .I1_1_0_0(n56_I1_1_0_0),
    .I1_2_0_0(n56_I1_2_0_0),
    .I1_3_0_0(n56_I1_3_0_0),
    .I1_4_0_0(n56_I1_4_0_0),
    .I1_5_0_0(n56_I1_5_0_0),
    .I1_6_0_0(n56_I1_6_0_0),
    .I1_7_0_0(n56_I1_7_0_0),
    .O_0_0_0_0(n56_O_0_0_0_0),
    .O_0_0_0_1(n56_O_0_0_0_1),
    .O_0_0_0_2(n56_O_0_0_0_2),
    .O_1_0_0_0(n56_O_1_0_0_0),
    .O_1_0_0_1(n56_O_1_0_0_1),
    .O_1_0_0_2(n56_O_1_0_0_2),
    .O_2_0_0_0(n56_O_2_0_0_0),
    .O_2_0_0_1(n56_O_2_0_0_1),
    .O_2_0_0_2(n56_O_2_0_0_2),
    .O_3_0_0_0(n56_O_3_0_0_0),
    .O_3_0_0_1(n56_O_3_0_0_1),
    .O_3_0_0_2(n56_O_3_0_0_2),
    .O_4_0_0_0(n56_O_4_0_0_0),
    .O_4_0_0_1(n56_O_4_0_0_1),
    .O_4_0_0_2(n56_O_4_0_0_2),
    .O_5_0_0_0(n56_O_5_0_0_0),
    .O_5_0_0_1(n56_O_5_0_0_1),
    .O_5_0_0_2(n56_O_5_0_0_2),
    .O_6_0_0_0(n56_O_6_0_0_0),
    .O_6_0_0_1(n56_O_6_0_0_1),
    .O_6_0_0_2(n56_O_6_0_0_2),
    .O_7_0_0_0(n56_O_7_0_0_0),
    .O_7_0_0_1(n56_O_7_0_0_1),
    .O_7_0_0_2(n56_O_7_0_0_2)
  );
  MapT n77 ( // @[Top.scala 84:21]
    .valid_up(n77_valid_up),
    .valid_down(n77_valid_down),
    .I_0_0_0_0(n77_I_0_0_0_0),
    .I_0_0_0_1(n77_I_0_0_0_1),
    .I_0_0_0_2(n77_I_0_0_0_2),
    .I_1_0_0_0(n77_I_1_0_0_0),
    .I_1_0_0_1(n77_I_1_0_0_1),
    .I_1_0_0_2(n77_I_1_0_0_2),
    .I_2_0_0_0(n77_I_2_0_0_0),
    .I_2_0_0_1(n77_I_2_0_0_1),
    .I_2_0_0_2(n77_I_2_0_0_2),
    .I_3_0_0_0(n77_I_3_0_0_0),
    .I_3_0_0_1(n77_I_3_0_0_1),
    .I_3_0_0_2(n77_I_3_0_0_2),
    .I_4_0_0_0(n77_I_4_0_0_0),
    .I_4_0_0_1(n77_I_4_0_0_1),
    .I_4_0_0_2(n77_I_4_0_0_2),
    .I_5_0_0_0(n77_I_5_0_0_0),
    .I_5_0_0_1(n77_I_5_0_0_1),
    .I_5_0_0_2(n77_I_5_0_0_2),
    .I_6_0_0_0(n77_I_6_0_0_0),
    .I_6_0_0_1(n77_I_6_0_0_1),
    .I_6_0_0_2(n77_I_6_0_0_2),
    .I_7_0_0_0(n77_I_7_0_0_0),
    .I_7_0_0_1(n77_I_7_0_0_1),
    .I_7_0_0_2(n77_I_7_0_0_2),
    .O_0_0_0(n77_O_0_0_0),
    .O_0_0_1(n77_O_0_0_1),
    .O_0_0_2(n77_O_0_0_2),
    .O_1_0_0(n77_O_1_0_0),
    .O_1_0_1(n77_O_1_0_1),
    .O_1_0_2(n77_O_1_0_2),
    .O_2_0_0(n77_O_2_0_0),
    .O_2_0_1(n77_O_2_0_1),
    .O_2_0_2(n77_O_2_0_2),
    .O_3_0_0(n77_O_3_0_0),
    .O_3_0_1(n77_O_3_0_1),
    .O_3_0_2(n77_O_3_0_2),
    .O_4_0_0(n77_O_4_0_0),
    .O_4_0_1(n77_O_4_0_1),
    .O_4_0_2(n77_O_4_0_2),
    .O_5_0_0(n77_O_5_0_0),
    .O_5_0_1(n77_O_5_0_1),
    .O_5_0_2(n77_O_5_0_2),
    .O_6_0_0(n77_O_6_0_0),
    .O_6_0_1(n77_O_6_0_1),
    .O_6_0_2(n77_O_6_0_2),
    .O_7_0_0(n77_O_7_0_0),
    .O_7_0_1(n77_O_7_0_1),
    .O_7_0_2(n77_O_7_0_2)
  );
  Map2T_4 n78 ( // @[Top.scala 87:21]
    .valid_up(n78_valid_up),
    .valid_down(n78_valid_down),
    .I0_0_0_0(n78_I0_0_0_0),
    .I0_0_0_1(n78_I0_0_0_1),
    .I0_0_0_2(n78_I0_0_0_2),
    .I0_1_0_0(n78_I0_1_0_0),
    .I0_1_0_1(n78_I0_1_0_1),
    .I0_1_0_2(n78_I0_1_0_2),
    .I0_2_0_0(n78_I0_2_0_0),
    .I0_2_0_1(n78_I0_2_0_1),
    .I0_2_0_2(n78_I0_2_0_2),
    .I0_3_0_0(n78_I0_3_0_0),
    .I0_3_0_1(n78_I0_3_0_1),
    .I0_3_0_2(n78_I0_3_0_2),
    .I0_4_0_0(n78_I0_4_0_0),
    .I0_4_0_1(n78_I0_4_0_1),
    .I0_4_0_2(n78_I0_4_0_2),
    .I0_5_0_0(n78_I0_5_0_0),
    .I0_5_0_1(n78_I0_5_0_1),
    .I0_5_0_2(n78_I0_5_0_2),
    .I0_6_0_0(n78_I0_6_0_0),
    .I0_6_0_1(n78_I0_6_0_1),
    .I0_6_0_2(n78_I0_6_0_2),
    .I0_7_0_0(n78_I0_7_0_0),
    .I0_7_0_1(n78_I0_7_0_1),
    .I0_7_0_2(n78_I0_7_0_2),
    .I1_0_0_0(n78_I1_0_0_0),
    .I1_0_0_1(n78_I1_0_0_1),
    .I1_0_0_2(n78_I1_0_0_2),
    .I1_1_0_0(n78_I1_1_0_0),
    .I1_1_0_1(n78_I1_1_0_1),
    .I1_1_0_2(n78_I1_1_0_2),
    .I1_2_0_0(n78_I1_2_0_0),
    .I1_2_0_1(n78_I1_2_0_1),
    .I1_2_0_2(n78_I1_2_0_2),
    .I1_3_0_0(n78_I1_3_0_0),
    .I1_3_0_1(n78_I1_3_0_1),
    .I1_3_0_2(n78_I1_3_0_2),
    .I1_4_0_0(n78_I1_4_0_0),
    .I1_4_0_1(n78_I1_4_0_1),
    .I1_4_0_2(n78_I1_4_0_2),
    .I1_5_0_0(n78_I1_5_0_0),
    .I1_5_0_1(n78_I1_5_0_1),
    .I1_5_0_2(n78_I1_5_0_2),
    .I1_6_0_0(n78_I1_6_0_0),
    .I1_6_0_1(n78_I1_6_0_1),
    .I1_6_0_2(n78_I1_6_0_2),
    .I1_7_0_0(n78_I1_7_0_0),
    .I1_7_0_1(n78_I1_7_0_1),
    .I1_7_0_2(n78_I1_7_0_2),
    .O_0_0_0_0(n78_O_0_0_0_0),
    .O_0_0_0_1(n78_O_0_0_0_1),
    .O_0_0_0_2(n78_O_0_0_0_2),
    .O_0_0_1_0(n78_O_0_0_1_0),
    .O_0_0_1_1(n78_O_0_0_1_1),
    .O_0_0_1_2(n78_O_0_0_1_2),
    .O_1_0_0_0(n78_O_1_0_0_0),
    .O_1_0_0_1(n78_O_1_0_0_1),
    .O_1_0_0_2(n78_O_1_0_0_2),
    .O_1_0_1_0(n78_O_1_0_1_0),
    .O_1_0_1_1(n78_O_1_0_1_1),
    .O_1_0_1_2(n78_O_1_0_1_2),
    .O_2_0_0_0(n78_O_2_0_0_0),
    .O_2_0_0_1(n78_O_2_0_0_1),
    .O_2_0_0_2(n78_O_2_0_0_2),
    .O_2_0_1_0(n78_O_2_0_1_0),
    .O_2_0_1_1(n78_O_2_0_1_1),
    .O_2_0_1_2(n78_O_2_0_1_2),
    .O_3_0_0_0(n78_O_3_0_0_0),
    .O_3_0_0_1(n78_O_3_0_0_1),
    .O_3_0_0_2(n78_O_3_0_0_2),
    .O_3_0_1_0(n78_O_3_0_1_0),
    .O_3_0_1_1(n78_O_3_0_1_1),
    .O_3_0_1_2(n78_O_3_0_1_2),
    .O_4_0_0_0(n78_O_4_0_0_0),
    .O_4_0_0_1(n78_O_4_0_0_1),
    .O_4_0_0_2(n78_O_4_0_0_2),
    .O_4_0_1_0(n78_O_4_0_1_0),
    .O_4_0_1_1(n78_O_4_0_1_1),
    .O_4_0_1_2(n78_O_4_0_1_2),
    .O_5_0_0_0(n78_O_5_0_0_0),
    .O_5_0_0_1(n78_O_5_0_0_1),
    .O_5_0_0_2(n78_O_5_0_0_2),
    .O_5_0_1_0(n78_O_5_0_1_0),
    .O_5_0_1_1(n78_O_5_0_1_1),
    .O_5_0_1_2(n78_O_5_0_1_2),
    .O_6_0_0_0(n78_O_6_0_0_0),
    .O_6_0_0_1(n78_O_6_0_0_1),
    .O_6_0_0_2(n78_O_6_0_0_2),
    .O_6_0_1_0(n78_O_6_0_1_0),
    .O_6_0_1_1(n78_O_6_0_1_1),
    .O_6_0_1_2(n78_O_6_0_1_2),
    .O_7_0_0_0(n78_O_7_0_0_0),
    .O_7_0_0_1(n78_O_7_0_0_1),
    .O_7_0_0_2(n78_O_7_0_0_2),
    .O_7_0_1_0(n78_O_7_0_1_0),
    .O_7_0_1_1(n78_O_7_0_1_1),
    .O_7_0_1_2(n78_O_7_0_1_2)
  );
  ShiftTS_2 n88 ( // @[Top.scala 91:21]
    .clock(n88_clock),
    .valid_up(n88_valid_up),
    .valid_down(n88_valid_down),
    .I_0_0_0(n88_I_0_0_0),
    .I_1_0_0(n88_I_1_0_0),
    .I_2_0_0(n88_I_2_0_0),
    .I_3_0_0(n88_I_3_0_0),
    .I_4_0_0(n88_I_4_0_0),
    .I_5_0_0(n88_I_5_0_0),
    .I_6_0_0(n88_I_6_0_0),
    .I_7_0_0(n88_I_7_0_0),
    .O_0_0_0(n88_O_0_0_0),
    .O_1_0_0(n88_O_1_0_0),
    .O_2_0_0(n88_O_2_0_0),
    .O_3_0_0(n88_O_3_0_0),
    .O_4_0_0(n88_O_4_0_0),
    .O_5_0_0(n88_O_5_0_0),
    .O_6_0_0(n88_O_6_0_0),
    .O_7_0_0(n88_O_7_0_0)
  );
  ShiftTS_2 n89 ( // @[Top.scala 94:21]
    .clock(n89_clock),
    .valid_up(n89_valid_up),
    .valid_down(n89_valid_down),
    .I_0_0_0(n89_I_0_0_0),
    .I_1_0_0(n89_I_1_0_0),
    .I_2_0_0(n89_I_2_0_0),
    .I_3_0_0(n89_I_3_0_0),
    .I_4_0_0(n89_I_4_0_0),
    .I_5_0_0(n89_I_5_0_0),
    .I_6_0_0(n89_I_6_0_0),
    .I_7_0_0(n89_I_7_0_0),
    .O_0_0_0(n89_O_0_0_0),
    .O_1_0_0(n89_O_1_0_0),
    .O_2_0_0(n89_O_2_0_0),
    .O_3_0_0(n89_O_3_0_0),
    .O_4_0_0(n89_O_4_0_0),
    .O_5_0_0(n89_O_5_0_0),
    .O_6_0_0(n89_O_6_0_0),
    .O_7_0_0(n89_O_7_0_0)
  );
  Map2T n90 ( // @[Top.scala 97:21]
    .valid_up(n90_valid_up),
    .valid_down(n90_valid_down),
    .I0_0_0_0(n90_I0_0_0_0),
    .I0_1_0_0(n90_I0_1_0_0),
    .I0_2_0_0(n90_I0_2_0_0),
    .I0_3_0_0(n90_I0_3_0_0),
    .I0_4_0_0(n90_I0_4_0_0),
    .I0_5_0_0(n90_I0_5_0_0),
    .I0_6_0_0(n90_I0_6_0_0),
    .I0_7_0_0(n90_I0_7_0_0),
    .I1_0_0_0(n90_I1_0_0_0),
    .I1_1_0_0(n90_I1_1_0_0),
    .I1_2_0_0(n90_I1_2_0_0),
    .I1_3_0_0(n90_I1_3_0_0),
    .I1_4_0_0(n90_I1_4_0_0),
    .I1_5_0_0(n90_I1_5_0_0),
    .I1_6_0_0(n90_I1_6_0_0),
    .I1_7_0_0(n90_I1_7_0_0),
    .O_0_0_0_0(n90_O_0_0_0_0),
    .O_0_0_0_1(n90_O_0_0_0_1),
    .O_1_0_0_0(n90_O_1_0_0_0),
    .O_1_0_0_1(n90_O_1_0_0_1),
    .O_2_0_0_0(n90_O_2_0_0_0),
    .O_2_0_0_1(n90_O_2_0_0_1),
    .O_3_0_0_0(n90_O_3_0_0_0),
    .O_3_0_0_1(n90_O_3_0_0_1),
    .O_4_0_0_0(n90_O_4_0_0_0),
    .O_4_0_0_1(n90_O_4_0_0_1),
    .O_5_0_0_0(n90_O_5_0_0_0),
    .O_5_0_0_1(n90_O_5_0_0_1),
    .O_6_0_0_0(n90_O_6_0_0_0),
    .O_6_0_0_1(n90_O_6_0_0_1),
    .O_7_0_0_0(n90_O_7_0_0_0),
    .O_7_0_0_1(n90_O_7_0_0_1)
  );
  Map2T_1 n103 ( // @[Top.scala 101:22]
    .valid_up(n103_valid_up),
    .valid_down(n103_valid_down),
    .I0_0_0_0_0(n103_I0_0_0_0_0),
    .I0_0_0_0_1(n103_I0_0_0_0_1),
    .I0_1_0_0_0(n103_I0_1_0_0_0),
    .I0_1_0_0_1(n103_I0_1_0_0_1),
    .I0_2_0_0_0(n103_I0_2_0_0_0),
    .I0_2_0_0_1(n103_I0_2_0_0_1),
    .I0_3_0_0_0(n103_I0_3_0_0_0),
    .I0_3_0_0_1(n103_I0_3_0_0_1),
    .I0_4_0_0_0(n103_I0_4_0_0_0),
    .I0_4_0_0_1(n103_I0_4_0_0_1),
    .I0_5_0_0_0(n103_I0_5_0_0_0),
    .I0_5_0_0_1(n103_I0_5_0_0_1),
    .I0_6_0_0_0(n103_I0_6_0_0_0),
    .I0_6_0_0_1(n103_I0_6_0_0_1),
    .I0_7_0_0_0(n103_I0_7_0_0_0),
    .I0_7_0_0_1(n103_I0_7_0_0_1),
    .I1_0_0_0(n103_I1_0_0_0),
    .I1_1_0_0(n103_I1_1_0_0),
    .I1_2_0_0(n103_I1_2_0_0),
    .I1_3_0_0(n103_I1_3_0_0),
    .I1_4_0_0(n103_I1_4_0_0),
    .I1_5_0_0(n103_I1_5_0_0),
    .I1_6_0_0(n103_I1_6_0_0),
    .I1_7_0_0(n103_I1_7_0_0),
    .O_0_0_0_0(n103_O_0_0_0_0),
    .O_0_0_0_1(n103_O_0_0_0_1),
    .O_0_0_0_2(n103_O_0_0_0_2),
    .O_1_0_0_0(n103_O_1_0_0_0),
    .O_1_0_0_1(n103_O_1_0_0_1),
    .O_1_0_0_2(n103_O_1_0_0_2),
    .O_2_0_0_0(n103_O_2_0_0_0),
    .O_2_0_0_1(n103_O_2_0_0_1),
    .O_2_0_0_2(n103_O_2_0_0_2),
    .O_3_0_0_0(n103_O_3_0_0_0),
    .O_3_0_0_1(n103_O_3_0_0_1),
    .O_3_0_0_2(n103_O_3_0_0_2),
    .O_4_0_0_0(n103_O_4_0_0_0),
    .O_4_0_0_1(n103_O_4_0_0_1),
    .O_4_0_0_2(n103_O_4_0_0_2),
    .O_5_0_0_0(n103_O_5_0_0_0),
    .O_5_0_0_1(n103_O_5_0_0_1),
    .O_5_0_0_2(n103_O_5_0_0_2),
    .O_6_0_0_0(n103_O_6_0_0_0),
    .O_6_0_0_1(n103_O_6_0_0_1),
    .O_6_0_0_2(n103_O_6_0_0_2),
    .O_7_0_0_0(n103_O_7_0_0_0),
    .O_7_0_0_1(n103_O_7_0_0_1),
    .O_7_0_0_2(n103_O_7_0_0_2)
  );
  MapT n124 ( // @[Top.scala 105:22]
    .valid_up(n124_valid_up),
    .valid_down(n124_valid_down),
    .I_0_0_0_0(n124_I_0_0_0_0),
    .I_0_0_0_1(n124_I_0_0_0_1),
    .I_0_0_0_2(n124_I_0_0_0_2),
    .I_1_0_0_0(n124_I_1_0_0_0),
    .I_1_0_0_1(n124_I_1_0_0_1),
    .I_1_0_0_2(n124_I_1_0_0_2),
    .I_2_0_0_0(n124_I_2_0_0_0),
    .I_2_0_0_1(n124_I_2_0_0_1),
    .I_2_0_0_2(n124_I_2_0_0_2),
    .I_3_0_0_0(n124_I_3_0_0_0),
    .I_3_0_0_1(n124_I_3_0_0_1),
    .I_3_0_0_2(n124_I_3_0_0_2),
    .I_4_0_0_0(n124_I_4_0_0_0),
    .I_4_0_0_1(n124_I_4_0_0_1),
    .I_4_0_0_2(n124_I_4_0_0_2),
    .I_5_0_0_0(n124_I_5_0_0_0),
    .I_5_0_0_1(n124_I_5_0_0_1),
    .I_5_0_0_2(n124_I_5_0_0_2),
    .I_6_0_0_0(n124_I_6_0_0_0),
    .I_6_0_0_1(n124_I_6_0_0_1),
    .I_6_0_0_2(n124_I_6_0_0_2),
    .I_7_0_0_0(n124_I_7_0_0_0),
    .I_7_0_0_1(n124_I_7_0_0_1),
    .I_7_0_0_2(n124_I_7_0_0_2),
    .O_0_0_0(n124_O_0_0_0),
    .O_0_0_1(n124_O_0_0_1),
    .O_0_0_2(n124_O_0_0_2),
    .O_1_0_0(n124_O_1_0_0),
    .O_1_0_1(n124_O_1_0_1),
    .O_1_0_2(n124_O_1_0_2),
    .O_2_0_0(n124_O_2_0_0),
    .O_2_0_1(n124_O_2_0_1),
    .O_2_0_2(n124_O_2_0_2),
    .O_3_0_0(n124_O_3_0_0),
    .O_3_0_1(n124_O_3_0_1),
    .O_3_0_2(n124_O_3_0_2),
    .O_4_0_0(n124_O_4_0_0),
    .O_4_0_1(n124_O_4_0_1),
    .O_4_0_2(n124_O_4_0_2),
    .O_5_0_0(n124_O_5_0_0),
    .O_5_0_1(n124_O_5_0_1),
    .O_5_0_2(n124_O_5_0_2),
    .O_6_0_0(n124_O_6_0_0),
    .O_6_0_1(n124_O_6_0_1),
    .O_6_0_2(n124_O_6_0_2),
    .O_7_0_0(n124_O_7_0_0),
    .O_7_0_1(n124_O_7_0_1),
    .O_7_0_2(n124_O_7_0_2)
  );
  Map2T_7 n125 ( // @[Top.scala 108:22]
    .valid_up(n125_valid_up),
    .valid_down(n125_valid_down),
    .I0_0_0_0_0(n125_I0_0_0_0_0),
    .I0_0_0_0_1(n125_I0_0_0_0_1),
    .I0_0_0_0_2(n125_I0_0_0_0_2),
    .I0_0_0_1_0(n125_I0_0_0_1_0),
    .I0_0_0_1_1(n125_I0_0_0_1_1),
    .I0_0_0_1_2(n125_I0_0_0_1_2),
    .I0_1_0_0_0(n125_I0_1_0_0_0),
    .I0_1_0_0_1(n125_I0_1_0_0_1),
    .I0_1_0_0_2(n125_I0_1_0_0_2),
    .I0_1_0_1_0(n125_I0_1_0_1_0),
    .I0_1_0_1_1(n125_I0_1_0_1_1),
    .I0_1_0_1_2(n125_I0_1_0_1_2),
    .I0_2_0_0_0(n125_I0_2_0_0_0),
    .I0_2_0_0_1(n125_I0_2_0_0_1),
    .I0_2_0_0_2(n125_I0_2_0_0_2),
    .I0_2_0_1_0(n125_I0_2_0_1_0),
    .I0_2_0_1_1(n125_I0_2_0_1_1),
    .I0_2_0_1_2(n125_I0_2_0_1_2),
    .I0_3_0_0_0(n125_I0_3_0_0_0),
    .I0_3_0_0_1(n125_I0_3_0_0_1),
    .I0_3_0_0_2(n125_I0_3_0_0_2),
    .I0_3_0_1_0(n125_I0_3_0_1_0),
    .I0_3_0_1_1(n125_I0_3_0_1_1),
    .I0_3_0_1_2(n125_I0_3_0_1_2),
    .I0_4_0_0_0(n125_I0_4_0_0_0),
    .I0_4_0_0_1(n125_I0_4_0_0_1),
    .I0_4_0_0_2(n125_I0_4_0_0_2),
    .I0_4_0_1_0(n125_I0_4_0_1_0),
    .I0_4_0_1_1(n125_I0_4_0_1_1),
    .I0_4_0_1_2(n125_I0_4_0_1_2),
    .I0_5_0_0_0(n125_I0_5_0_0_0),
    .I0_5_0_0_1(n125_I0_5_0_0_1),
    .I0_5_0_0_2(n125_I0_5_0_0_2),
    .I0_5_0_1_0(n125_I0_5_0_1_0),
    .I0_5_0_1_1(n125_I0_5_0_1_1),
    .I0_5_0_1_2(n125_I0_5_0_1_2),
    .I0_6_0_0_0(n125_I0_6_0_0_0),
    .I0_6_0_0_1(n125_I0_6_0_0_1),
    .I0_6_0_0_2(n125_I0_6_0_0_2),
    .I0_6_0_1_0(n125_I0_6_0_1_0),
    .I0_6_0_1_1(n125_I0_6_0_1_1),
    .I0_6_0_1_2(n125_I0_6_0_1_2),
    .I0_7_0_0_0(n125_I0_7_0_0_0),
    .I0_7_0_0_1(n125_I0_7_0_0_1),
    .I0_7_0_0_2(n125_I0_7_0_0_2),
    .I0_7_0_1_0(n125_I0_7_0_1_0),
    .I0_7_0_1_1(n125_I0_7_0_1_1),
    .I0_7_0_1_2(n125_I0_7_0_1_2),
    .I1_0_0_0(n125_I1_0_0_0),
    .I1_0_0_1(n125_I1_0_0_1),
    .I1_0_0_2(n125_I1_0_0_2),
    .I1_1_0_0(n125_I1_1_0_0),
    .I1_1_0_1(n125_I1_1_0_1),
    .I1_1_0_2(n125_I1_1_0_2),
    .I1_2_0_0(n125_I1_2_0_0),
    .I1_2_0_1(n125_I1_2_0_1),
    .I1_2_0_2(n125_I1_2_0_2),
    .I1_3_0_0(n125_I1_3_0_0),
    .I1_3_0_1(n125_I1_3_0_1),
    .I1_3_0_2(n125_I1_3_0_2),
    .I1_4_0_0(n125_I1_4_0_0),
    .I1_4_0_1(n125_I1_4_0_1),
    .I1_4_0_2(n125_I1_4_0_2),
    .I1_5_0_0(n125_I1_5_0_0),
    .I1_5_0_1(n125_I1_5_0_1),
    .I1_5_0_2(n125_I1_5_0_2),
    .I1_6_0_0(n125_I1_6_0_0),
    .I1_6_0_1(n125_I1_6_0_1),
    .I1_6_0_2(n125_I1_6_0_2),
    .I1_7_0_0(n125_I1_7_0_0),
    .I1_7_0_1(n125_I1_7_0_1),
    .I1_7_0_2(n125_I1_7_0_2),
    .O_0_0_0_0(n125_O_0_0_0_0),
    .O_0_0_0_1(n125_O_0_0_0_1),
    .O_0_0_0_2(n125_O_0_0_0_2),
    .O_0_0_1_0(n125_O_0_0_1_0),
    .O_0_0_1_1(n125_O_0_0_1_1),
    .O_0_0_1_2(n125_O_0_0_1_2),
    .O_0_0_2_0(n125_O_0_0_2_0),
    .O_0_0_2_1(n125_O_0_0_2_1),
    .O_0_0_2_2(n125_O_0_0_2_2),
    .O_1_0_0_0(n125_O_1_0_0_0),
    .O_1_0_0_1(n125_O_1_0_0_1),
    .O_1_0_0_2(n125_O_1_0_0_2),
    .O_1_0_1_0(n125_O_1_0_1_0),
    .O_1_0_1_1(n125_O_1_0_1_1),
    .O_1_0_1_2(n125_O_1_0_1_2),
    .O_1_0_2_0(n125_O_1_0_2_0),
    .O_1_0_2_1(n125_O_1_0_2_1),
    .O_1_0_2_2(n125_O_1_0_2_2),
    .O_2_0_0_0(n125_O_2_0_0_0),
    .O_2_0_0_1(n125_O_2_0_0_1),
    .O_2_0_0_2(n125_O_2_0_0_2),
    .O_2_0_1_0(n125_O_2_0_1_0),
    .O_2_0_1_1(n125_O_2_0_1_1),
    .O_2_0_1_2(n125_O_2_0_1_2),
    .O_2_0_2_0(n125_O_2_0_2_0),
    .O_2_0_2_1(n125_O_2_0_2_1),
    .O_2_0_2_2(n125_O_2_0_2_2),
    .O_3_0_0_0(n125_O_3_0_0_0),
    .O_3_0_0_1(n125_O_3_0_0_1),
    .O_3_0_0_2(n125_O_3_0_0_2),
    .O_3_0_1_0(n125_O_3_0_1_0),
    .O_3_0_1_1(n125_O_3_0_1_1),
    .O_3_0_1_2(n125_O_3_0_1_2),
    .O_3_0_2_0(n125_O_3_0_2_0),
    .O_3_0_2_1(n125_O_3_0_2_1),
    .O_3_0_2_2(n125_O_3_0_2_2),
    .O_4_0_0_0(n125_O_4_0_0_0),
    .O_4_0_0_1(n125_O_4_0_0_1),
    .O_4_0_0_2(n125_O_4_0_0_2),
    .O_4_0_1_0(n125_O_4_0_1_0),
    .O_4_0_1_1(n125_O_4_0_1_1),
    .O_4_0_1_2(n125_O_4_0_1_2),
    .O_4_0_2_0(n125_O_4_0_2_0),
    .O_4_0_2_1(n125_O_4_0_2_1),
    .O_4_0_2_2(n125_O_4_0_2_2),
    .O_5_0_0_0(n125_O_5_0_0_0),
    .O_5_0_0_1(n125_O_5_0_0_1),
    .O_5_0_0_2(n125_O_5_0_0_2),
    .O_5_0_1_0(n125_O_5_0_1_0),
    .O_5_0_1_1(n125_O_5_0_1_1),
    .O_5_0_1_2(n125_O_5_0_1_2),
    .O_5_0_2_0(n125_O_5_0_2_0),
    .O_5_0_2_1(n125_O_5_0_2_1),
    .O_5_0_2_2(n125_O_5_0_2_2),
    .O_6_0_0_0(n125_O_6_0_0_0),
    .O_6_0_0_1(n125_O_6_0_0_1),
    .O_6_0_0_2(n125_O_6_0_0_2),
    .O_6_0_1_0(n125_O_6_0_1_0),
    .O_6_0_1_1(n125_O_6_0_1_1),
    .O_6_0_1_2(n125_O_6_0_1_2),
    .O_6_0_2_0(n125_O_6_0_2_0),
    .O_6_0_2_1(n125_O_6_0_2_1),
    .O_6_0_2_2(n125_O_6_0_2_2),
    .O_7_0_0_0(n125_O_7_0_0_0),
    .O_7_0_0_1(n125_O_7_0_0_1),
    .O_7_0_0_2(n125_O_7_0_0_2),
    .O_7_0_1_0(n125_O_7_0_1_0),
    .O_7_0_1_1(n125_O_7_0_1_1),
    .O_7_0_1_2(n125_O_7_0_1_2),
    .O_7_0_2_0(n125_O_7_0_2_0),
    .O_7_0_2_1(n125_O_7_0_2_1),
    .O_7_0_2_2(n125_O_7_0_2_2)
  );
  MapT_3 n141 ( // @[Top.scala 112:22]
    .valid_up(n141_valid_up),
    .valid_down(n141_valid_down),
    .I_0_0_0_0(n141_I_0_0_0_0),
    .I_0_0_0_1(n141_I_0_0_0_1),
    .I_0_0_0_2(n141_I_0_0_0_2),
    .I_0_0_1_0(n141_I_0_0_1_0),
    .I_0_0_1_1(n141_I_0_0_1_1),
    .I_0_0_1_2(n141_I_0_0_1_2),
    .I_0_0_2_0(n141_I_0_0_2_0),
    .I_0_0_2_1(n141_I_0_0_2_1),
    .I_0_0_2_2(n141_I_0_0_2_2),
    .I_1_0_0_0(n141_I_1_0_0_0),
    .I_1_0_0_1(n141_I_1_0_0_1),
    .I_1_0_0_2(n141_I_1_0_0_2),
    .I_1_0_1_0(n141_I_1_0_1_0),
    .I_1_0_1_1(n141_I_1_0_1_1),
    .I_1_0_1_2(n141_I_1_0_1_2),
    .I_1_0_2_0(n141_I_1_0_2_0),
    .I_1_0_2_1(n141_I_1_0_2_1),
    .I_1_0_2_2(n141_I_1_0_2_2),
    .I_2_0_0_0(n141_I_2_0_0_0),
    .I_2_0_0_1(n141_I_2_0_0_1),
    .I_2_0_0_2(n141_I_2_0_0_2),
    .I_2_0_1_0(n141_I_2_0_1_0),
    .I_2_0_1_1(n141_I_2_0_1_1),
    .I_2_0_1_2(n141_I_2_0_1_2),
    .I_2_0_2_0(n141_I_2_0_2_0),
    .I_2_0_2_1(n141_I_2_0_2_1),
    .I_2_0_2_2(n141_I_2_0_2_2),
    .I_3_0_0_0(n141_I_3_0_0_0),
    .I_3_0_0_1(n141_I_3_0_0_1),
    .I_3_0_0_2(n141_I_3_0_0_2),
    .I_3_0_1_0(n141_I_3_0_1_0),
    .I_3_0_1_1(n141_I_3_0_1_1),
    .I_3_0_1_2(n141_I_3_0_1_2),
    .I_3_0_2_0(n141_I_3_0_2_0),
    .I_3_0_2_1(n141_I_3_0_2_1),
    .I_3_0_2_2(n141_I_3_0_2_2),
    .I_4_0_0_0(n141_I_4_0_0_0),
    .I_4_0_0_1(n141_I_4_0_0_1),
    .I_4_0_0_2(n141_I_4_0_0_2),
    .I_4_0_1_0(n141_I_4_0_1_0),
    .I_4_0_1_1(n141_I_4_0_1_1),
    .I_4_0_1_2(n141_I_4_0_1_2),
    .I_4_0_2_0(n141_I_4_0_2_0),
    .I_4_0_2_1(n141_I_4_0_2_1),
    .I_4_0_2_2(n141_I_4_0_2_2),
    .I_5_0_0_0(n141_I_5_0_0_0),
    .I_5_0_0_1(n141_I_5_0_0_1),
    .I_5_0_0_2(n141_I_5_0_0_2),
    .I_5_0_1_0(n141_I_5_0_1_0),
    .I_5_0_1_1(n141_I_5_0_1_1),
    .I_5_0_1_2(n141_I_5_0_1_2),
    .I_5_0_2_0(n141_I_5_0_2_0),
    .I_5_0_2_1(n141_I_5_0_2_1),
    .I_5_0_2_2(n141_I_5_0_2_2),
    .I_6_0_0_0(n141_I_6_0_0_0),
    .I_6_0_0_1(n141_I_6_0_0_1),
    .I_6_0_0_2(n141_I_6_0_0_2),
    .I_6_0_1_0(n141_I_6_0_1_0),
    .I_6_0_1_1(n141_I_6_0_1_1),
    .I_6_0_1_2(n141_I_6_0_1_2),
    .I_6_0_2_0(n141_I_6_0_2_0),
    .I_6_0_2_1(n141_I_6_0_2_1),
    .I_6_0_2_2(n141_I_6_0_2_2),
    .I_7_0_0_0(n141_I_7_0_0_0),
    .I_7_0_0_1(n141_I_7_0_0_1),
    .I_7_0_0_2(n141_I_7_0_0_2),
    .I_7_0_1_0(n141_I_7_0_1_0),
    .I_7_0_1_1(n141_I_7_0_1_1),
    .I_7_0_1_2(n141_I_7_0_1_2),
    .I_7_0_2_0(n141_I_7_0_2_0),
    .I_7_0_2_1(n141_I_7_0_2_1),
    .I_7_0_2_2(n141_I_7_0_2_2),
    .O_0_0_0(n141_O_0_0_0),
    .O_0_0_1(n141_O_0_0_1),
    .O_0_0_2(n141_O_0_0_2),
    .O_0_1_0(n141_O_0_1_0),
    .O_0_1_1(n141_O_0_1_1),
    .O_0_1_2(n141_O_0_1_2),
    .O_0_2_0(n141_O_0_2_0),
    .O_0_2_1(n141_O_0_2_1),
    .O_0_2_2(n141_O_0_2_2),
    .O_1_0_0(n141_O_1_0_0),
    .O_1_0_1(n141_O_1_0_1),
    .O_1_0_2(n141_O_1_0_2),
    .O_1_1_0(n141_O_1_1_0),
    .O_1_1_1(n141_O_1_1_1),
    .O_1_1_2(n141_O_1_1_2),
    .O_1_2_0(n141_O_1_2_0),
    .O_1_2_1(n141_O_1_2_1),
    .O_1_2_2(n141_O_1_2_2),
    .O_2_0_0(n141_O_2_0_0),
    .O_2_0_1(n141_O_2_0_1),
    .O_2_0_2(n141_O_2_0_2),
    .O_2_1_0(n141_O_2_1_0),
    .O_2_1_1(n141_O_2_1_1),
    .O_2_1_2(n141_O_2_1_2),
    .O_2_2_0(n141_O_2_2_0),
    .O_2_2_1(n141_O_2_2_1),
    .O_2_2_2(n141_O_2_2_2),
    .O_3_0_0(n141_O_3_0_0),
    .O_3_0_1(n141_O_3_0_1),
    .O_3_0_2(n141_O_3_0_2),
    .O_3_1_0(n141_O_3_1_0),
    .O_3_1_1(n141_O_3_1_1),
    .O_3_1_2(n141_O_3_1_2),
    .O_3_2_0(n141_O_3_2_0),
    .O_3_2_1(n141_O_3_2_1),
    .O_3_2_2(n141_O_3_2_2),
    .O_4_0_0(n141_O_4_0_0),
    .O_4_0_1(n141_O_4_0_1),
    .O_4_0_2(n141_O_4_0_2),
    .O_4_1_0(n141_O_4_1_0),
    .O_4_1_1(n141_O_4_1_1),
    .O_4_1_2(n141_O_4_1_2),
    .O_4_2_0(n141_O_4_2_0),
    .O_4_2_1(n141_O_4_2_1),
    .O_4_2_2(n141_O_4_2_2),
    .O_5_0_0(n141_O_5_0_0),
    .O_5_0_1(n141_O_5_0_1),
    .O_5_0_2(n141_O_5_0_2),
    .O_5_1_0(n141_O_5_1_0),
    .O_5_1_1(n141_O_5_1_1),
    .O_5_1_2(n141_O_5_1_2),
    .O_5_2_0(n141_O_5_2_0),
    .O_5_2_1(n141_O_5_2_1),
    .O_5_2_2(n141_O_5_2_2),
    .O_6_0_0(n141_O_6_0_0),
    .O_6_0_1(n141_O_6_0_1),
    .O_6_0_2(n141_O_6_0_2),
    .O_6_1_0(n141_O_6_1_0),
    .O_6_1_1(n141_O_6_1_1),
    .O_6_1_2(n141_O_6_1_2),
    .O_6_2_0(n141_O_6_2_0),
    .O_6_2_1(n141_O_6_2_1),
    .O_6_2_2(n141_O_6_2_2),
    .O_7_0_0(n141_O_7_0_0),
    .O_7_0_1(n141_O_7_0_1),
    .O_7_0_2(n141_O_7_0_2),
    .O_7_1_0(n141_O_7_1_0),
    .O_7_1_1(n141_O_7_1_1),
    .O_7_1_2(n141_O_7_1_2),
    .O_7_2_0(n141_O_7_2_0),
    .O_7_2_1(n141_O_7_2_1),
    .O_7_2_2(n141_O_7_2_2)
  );
  MapT_4 n183 ( // @[Top.scala 115:22]
    .clock(n183_clock),
    .reset(n183_reset),
    .valid_up(n183_valid_up),
    .valid_down(n183_valid_down),
    .I_0_0_0(n183_I_0_0_0),
    .I_0_0_1(n183_I_0_0_1),
    .I_0_0_2(n183_I_0_0_2),
    .I_0_1_0(n183_I_0_1_0),
    .I_0_1_1(n183_I_0_1_1),
    .I_0_1_2(n183_I_0_1_2),
    .I_0_2_0(n183_I_0_2_0),
    .I_0_2_1(n183_I_0_2_1),
    .I_0_2_2(n183_I_0_2_2),
    .I_1_0_0(n183_I_1_0_0),
    .I_1_0_1(n183_I_1_0_1),
    .I_1_0_2(n183_I_1_0_2),
    .I_1_1_0(n183_I_1_1_0),
    .I_1_1_1(n183_I_1_1_1),
    .I_1_1_2(n183_I_1_1_2),
    .I_1_2_0(n183_I_1_2_0),
    .I_1_2_1(n183_I_1_2_1),
    .I_1_2_2(n183_I_1_2_2),
    .I_2_0_0(n183_I_2_0_0),
    .I_2_0_1(n183_I_2_0_1),
    .I_2_0_2(n183_I_2_0_2),
    .I_2_1_0(n183_I_2_1_0),
    .I_2_1_1(n183_I_2_1_1),
    .I_2_1_2(n183_I_2_1_2),
    .I_2_2_0(n183_I_2_2_0),
    .I_2_2_1(n183_I_2_2_1),
    .I_2_2_2(n183_I_2_2_2),
    .I_3_0_0(n183_I_3_0_0),
    .I_3_0_1(n183_I_3_0_1),
    .I_3_0_2(n183_I_3_0_2),
    .I_3_1_0(n183_I_3_1_0),
    .I_3_1_1(n183_I_3_1_1),
    .I_3_1_2(n183_I_3_1_2),
    .I_3_2_0(n183_I_3_2_0),
    .I_3_2_1(n183_I_3_2_1),
    .I_3_2_2(n183_I_3_2_2),
    .I_4_0_0(n183_I_4_0_0),
    .I_4_0_1(n183_I_4_0_1),
    .I_4_0_2(n183_I_4_0_2),
    .I_4_1_0(n183_I_4_1_0),
    .I_4_1_1(n183_I_4_1_1),
    .I_4_1_2(n183_I_4_1_2),
    .I_4_2_0(n183_I_4_2_0),
    .I_4_2_1(n183_I_4_2_1),
    .I_4_2_2(n183_I_4_2_2),
    .I_5_0_0(n183_I_5_0_0),
    .I_5_0_1(n183_I_5_0_1),
    .I_5_0_2(n183_I_5_0_2),
    .I_5_1_0(n183_I_5_1_0),
    .I_5_1_1(n183_I_5_1_1),
    .I_5_1_2(n183_I_5_1_2),
    .I_5_2_0(n183_I_5_2_0),
    .I_5_2_1(n183_I_5_2_1),
    .I_5_2_2(n183_I_5_2_2),
    .I_6_0_0(n183_I_6_0_0),
    .I_6_0_1(n183_I_6_0_1),
    .I_6_0_2(n183_I_6_0_2),
    .I_6_1_0(n183_I_6_1_0),
    .I_6_1_1(n183_I_6_1_1),
    .I_6_1_2(n183_I_6_1_2),
    .I_6_2_0(n183_I_6_2_0),
    .I_6_2_1(n183_I_6_2_1),
    .I_6_2_2(n183_I_6_2_2),
    .I_7_0_0(n183_I_7_0_0),
    .I_7_0_1(n183_I_7_0_1),
    .I_7_0_2(n183_I_7_0_2),
    .I_7_1_0(n183_I_7_1_0),
    .I_7_1_1(n183_I_7_1_1),
    .I_7_1_2(n183_I_7_1_2),
    .I_7_2_0(n183_I_7_2_0),
    .I_7_2_1(n183_I_7_2_1),
    .I_7_2_2(n183_I_7_2_2),
    .O_0_0_0(n183_O_0_0_0),
    .O_1_0_0(n183_O_1_0_0),
    .O_2_0_0(n183_O_2_0_0),
    .O_3_0_0(n183_O_3_0_0),
    .O_4_0_0(n183_O_4_0_0),
    .O_5_0_0(n183_O_5_0_0),
    .O_6_0_0(n183_O_6_0_0),
    .O_7_0_0(n183_O_7_0_0)
  );
  FIFO n184 ( // @[Top.scala 118:22]
    .clock(n184_clock),
    .valid_up(n184_valid_up),
    .valid_down(n184_valid_down),
    .I_0_0_0(n184_I_0_0_0),
    .I_1_0_0(n184_I_1_0_0),
    .I_2_0_0(n184_I_2_0_0),
    .I_3_0_0(n184_I_3_0_0),
    .I_4_0_0(n184_I_4_0_0),
    .I_5_0_0(n184_I_5_0_0),
    .I_6_0_0(n184_I_6_0_0),
    .I_7_0_0(n184_I_7_0_0),
    .O_0_0_0(n184_O_0_0_0),
    .O_1_0_0(n184_O_1_0_0),
    .O_2_0_0(n184_O_2_0_0),
    .O_3_0_0(n184_O_3_0_0),
    .O_4_0_0(n184_O_4_0_0),
    .O_5_0_0(n184_O_5_0_0),
    .O_6_0_0(n184_O_6_0_0),
    .O_7_0_0(n184_O_7_0_0)
  );
  FIFO n185 ( // @[Top.scala 121:22]
    .clock(n185_clock),
    .valid_up(n185_valid_up),
    .valid_down(n185_valid_down),
    .I_0_0_0(n185_I_0_0_0),
    .I_1_0_0(n185_I_1_0_0),
    .I_2_0_0(n185_I_2_0_0),
    .I_3_0_0(n185_I_3_0_0),
    .I_4_0_0(n185_I_4_0_0),
    .I_5_0_0(n185_I_5_0_0),
    .I_6_0_0(n185_I_6_0_0),
    .I_7_0_0(n185_I_7_0_0),
    .O_0_0_0(n185_O_0_0_0),
    .O_1_0_0(n185_O_1_0_0),
    .O_2_0_0(n185_O_2_0_0),
    .O_3_0_0(n185_O_3_0_0),
    .O_4_0_0(n185_O_4_0_0),
    .O_5_0_0(n185_O_5_0_0),
    .O_6_0_0(n185_O_6_0_0),
    .O_7_0_0(n185_O_7_0_0)
  );
  FIFO n186 ( // @[Top.scala 124:22]
    .clock(n186_clock),
    .valid_up(n186_valid_up),
    .valid_down(n186_valid_down),
    .I_0_0_0(n186_I_0_0_0),
    .I_1_0_0(n186_I_1_0_0),
    .I_2_0_0(n186_I_2_0_0),
    .I_3_0_0(n186_I_3_0_0),
    .I_4_0_0(n186_I_4_0_0),
    .I_5_0_0(n186_I_5_0_0),
    .I_6_0_0(n186_I_6_0_0),
    .I_7_0_0(n186_I_7_0_0),
    .O_0_0_0(n186_O_0_0_0),
    .O_1_0_0(n186_O_1_0_0),
    .O_2_0_0(n186_O_2_0_0),
    .O_3_0_0(n186_O_3_0_0),
    .O_4_0_0(n186_O_4_0_0),
    .O_5_0_0(n186_O_5_0_0),
    .O_6_0_0(n186_O_6_0_0),
    .O_7_0_0(n186_O_7_0_0)
  );
  assign valid_down = n186_valid_down; // @[Top.scala 128:16]
  assign O_0_0_0 = n186_O_0_0_0; // @[Top.scala 127:7]
  assign O_1_0_0 = n186_O_1_0_0; // @[Top.scala 127:7]
  assign O_2_0_0 = n186_O_2_0_0; // @[Top.scala 127:7]
  assign O_3_0_0 = n186_O_3_0_0; // @[Top.scala 127:7]
  assign O_4_0_0 = n186_O_4_0_0; // @[Top.scala 127:7]
  assign O_5_0_0 = n186_O_5_0_0; // @[Top.scala 127:7]
  assign O_6_0_0 = n186_O_6_0_0; // @[Top.scala 127:7]
  assign O_7_0_0 = n186_O_7_0_0; // @[Top.scala 127:7]
  assign n1_clock = clock;
  assign n1_valid_up = valid_up; // @[Top.scala 46:17]
  assign n1_I_0_0_0 = I_0_0_0; // @[Top.scala 45:10]
  assign n1_I_1_0_0 = I_1_0_0; // @[Top.scala 45:10]
  assign n1_I_2_0_0 = I_2_0_0; // @[Top.scala 45:10]
  assign n1_I_3_0_0 = I_3_0_0; // @[Top.scala 45:10]
  assign n1_I_4_0_0 = I_4_0_0; // @[Top.scala 45:10]
  assign n1_I_5_0_0 = I_5_0_0; // @[Top.scala 45:10]
  assign n1_I_6_0_0 = I_6_0_0; // @[Top.scala 45:10]
  assign n1_I_7_0_0 = I_7_0_0; // @[Top.scala 45:10]
  assign n2_clock = clock;
  assign n2_reset = reset;
  assign n2_valid_up = n1_valid_down; // @[Top.scala 49:17]
  assign n2_I_0_0_0 = n1_O_0_0_0; // @[Top.scala 48:10]
  assign n2_I_1_0_0 = n1_O_1_0_0; // @[Top.scala 48:10]
  assign n2_I_2_0_0 = n1_O_2_0_0; // @[Top.scala 48:10]
  assign n2_I_3_0_0 = n1_O_3_0_0; // @[Top.scala 48:10]
  assign n2_I_4_0_0 = n1_O_4_0_0; // @[Top.scala 48:10]
  assign n2_I_5_0_0 = n1_O_5_0_0; // @[Top.scala 48:10]
  assign n2_I_6_0_0 = n1_O_6_0_0; // @[Top.scala 48:10]
  assign n2_I_7_0_0 = n1_O_7_0_0; // @[Top.scala 48:10]
  assign n3_clock = clock;
  assign n3_reset = reset;
  assign n3_valid_up = n2_valid_down; // @[Top.scala 52:17]
  assign n3_I_0_0_0 = n2_O_0_0_0; // @[Top.scala 51:10]
  assign n3_I_1_0_0 = n2_O_1_0_0; // @[Top.scala 51:10]
  assign n3_I_2_0_0 = n2_O_2_0_0; // @[Top.scala 51:10]
  assign n3_I_3_0_0 = n2_O_3_0_0; // @[Top.scala 51:10]
  assign n3_I_4_0_0 = n2_O_4_0_0; // @[Top.scala 51:10]
  assign n3_I_5_0_0 = n2_O_5_0_0; // @[Top.scala 51:10]
  assign n3_I_6_0_0 = n2_O_6_0_0; // @[Top.scala 51:10]
  assign n3_I_7_0_0 = n2_O_7_0_0; // @[Top.scala 51:10]
  assign n4_clock = clock;
  assign n4_valid_up = n3_valid_down; // @[Top.scala 55:17]
  assign n4_I_0_0_0 = n3_O_0_0_0; // @[Top.scala 54:10]
  assign n4_I_1_0_0 = n3_O_1_0_0; // @[Top.scala 54:10]
  assign n4_I_2_0_0 = n3_O_2_0_0; // @[Top.scala 54:10]
  assign n4_I_3_0_0 = n3_O_3_0_0; // @[Top.scala 54:10]
  assign n4_I_4_0_0 = n3_O_4_0_0; // @[Top.scala 54:10]
  assign n4_I_5_0_0 = n3_O_5_0_0; // @[Top.scala 54:10]
  assign n4_I_6_0_0 = n3_O_6_0_0; // @[Top.scala 54:10]
  assign n4_I_7_0_0 = n3_O_7_0_0; // @[Top.scala 54:10]
  assign n5_clock = clock;
  assign n5_valid_up = n4_valid_down; // @[Top.scala 58:17]
  assign n5_I_0_0_0 = n4_O_0_0_0; // @[Top.scala 57:10]
  assign n5_I_1_0_0 = n4_O_1_0_0; // @[Top.scala 57:10]
  assign n5_I_2_0_0 = n4_O_2_0_0; // @[Top.scala 57:10]
  assign n5_I_3_0_0 = n4_O_3_0_0; // @[Top.scala 57:10]
  assign n5_I_4_0_0 = n4_O_4_0_0; // @[Top.scala 57:10]
  assign n5_I_5_0_0 = n4_O_5_0_0; // @[Top.scala 57:10]
  assign n5_I_6_0_0 = n4_O_6_0_0; // @[Top.scala 57:10]
  assign n5_I_7_0_0 = n4_O_7_0_0; // @[Top.scala 57:10]
  assign n6_valid_up = n5_valid_down & n4_valid_down; // @[Top.scala 62:17]
  assign n6_I0_0_0_0 = n5_O_0_0_0; // @[Top.scala 60:11]
  assign n6_I0_1_0_0 = n5_O_1_0_0; // @[Top.scala 60:11]
  assign n6_I0_2_0_0 = n5_O_2_0_0; // @[Top.scala 60:11]
  assign n6_I0_3_0_0 = n5_O_3_0_0; // @[Top.scala 60:11]
  assign n6_I0_4_0_0 = n5_O_4_0_0; // @[Top.scala 60:11]
  assign n6_I0_5_0_0 = n5_O_5_0_0; // @[Top.scala 60:11]
  assign n6_I0_6_0_0 = n5_O_6_0_0; // @[Top.scala 60:11]
  assign n6_I0_7_0_0 = n5_O_7_0_0; // @[Top.scala 60:11]
  assign n6_I1_0_0_0 = n4_O_0_0_0; // @[Top.scala 61:11]
  assign n6_I1_1_0_0 = n4_O_1_0_0; // @[Top.scala 61:11]
  assign n6_I1_2_0_0 = n4_O_2_0_0; // @[Top.scala 61:11]
  assign n6_I1_3_0_0 = n4_O_3_0_0; // @[Top.scala 61:11]
  assign n6_I1_4_0_0 = n4_O_4_0_0; // @[Top.scala 61:11]
  assign n6_I1_5_0_0 = n4_O_5_0_0; // @[Top.scala 61:11]
  assign n6_I1_6_0_0 = n4_O_6_0_0; // @[Top.scala 61:11]
  assign n6_I1_7_0_0 = n4_O_7_0_0; // @[Top.scala 61:11]
  assign n19_valid_up = n6_valid_down & n3_valid_down; // @[Top.scala 66:18]
  assign n19_I0_0_0_0_0 = n6_O_0_0_0_0; // @[Top.scala 64:12]
  assign n19_I0_0_0_0_1 = n6_O_0_0_0_1; // @[Top.scala 64:12]
  assign n19_I0_1_0_0_0 = n6_O_1_0_0_0; // @[Top.scala 64:12]
  assign n19_I0_1_0_0_1 = n6_O_1_0_0_1; // @[Top.scala 64:12]
  assign n19_I0_2_0_0_0 = n6_O_2_0_0_0; // @[Top.scala 64:12]
  assign n19_I0_2_0_0_1 = n6_O_2_0_0_1; // @[Top.scala 64:12]
  assign n19_I0_3_0_0_0 = n6_O_3_0_0_0; // @[Top.scala 64:12]
  assign n19_I0_3_0_0_1 = n6_O_3_0_0_1; // @[Top.scala 64:12]
  assign n19_I0_4_0_0_0 = n6_O_4_0_0_0; // @[Top.scala 64:12]
  assign n19_I0_4_0_0_1 = n6_O_4_0_0_1; // @[Top.scala 64:12]
  assign n19_I0_5_0_0_0 = n6_O_5_0_0_0; // @[Top.scala 64:12]
  assign n19_I0_5_0_0_1 = n6_O_5_0_0_1; // @[Top.scala 64:12]
  assign n19_I0_6_0_0_0 = n6_O_6_0_0_0; // @[Top.scala 64:12]
  assign n19_I0_6_0_0_1 = n6_O_6_0_0_1; // @[Top.scala 64:12]
  assign n19_I0_7_0_0_0 = n6_O_7_0_0_0; // @[Top.scala 64:12]
  assign n19_I0_7_0_0_1 = n6_O_7_0_0_1; // @[Top.scala 64:12]
  assign n19_I1_0_0_0 = n3_O_0_0_0; // @[Top.scala 65:12]
  assign n19_I1_1_0_0 = n3_O_1_0_0; // @[Top.scala 65:12]
  assign n19_I1_2_0_0 = n3_O_2_0_0; // @[Top.scala 65:12]
  assign n19_I1_3_0_0 = n3_O_3_0_0; // @[Top.scala 65:12]
  assign n19_I1_4_0_0 = n3_O_4_0_0; // @[Top.scala 65:12]
  assign n19_I1_5_0_0 = n3_O_5_0_0; // @[Top.scala 65:12]
  assign n19_I1_6_0_0 = n3_O_6_0_0; // @[Top.scala 65:12]
  assign n19_I1_7_0_0 = n3_O_7_0_0; // @[Top.scala 65:12]
  assign n40_valid_up = n19_valid_down; // @[Top.scala 69:18]
  assign n40_I_0_0_0_0 = n19_O_0_0_0_0; // @[Top.scala 68:11]
  assign n40_I_0_0_0_1 = n19_O_0_0_0_1; // @[Top.scala 68:11]
  assign n40_I_0_0_0_2 = n19_O_0_0_0_2; // @[Top.scala 68:11]
  assign n40_I_1_0_0_0 = n19_O_1_0_0_0; // @[Top.scala 68:11]
  assign n40_I_1_0_0_1 = n19_O_1_0_0_1; // @[Top.scala 68:11]
  assign n40_I_1_0_0_2 = n19_O_1_0_0_2; // @[Top.scala 68:11]
  assign n40_I_2_0_0_0 = n19_O_2_0_0_0; // @[Top.scala 68:11]
  assign n40_I_2_0_0_1 = n19_O_2_0_0_1; // @[Top.scala 68:11]
  assign n40_I_2_0_0_2 = n19_O_2_0_0_2; // @[Top.scala 68:11]
  assign n40_I_3_0_0_0 = n19_O_3_0_0_0; // @[Top.scala 68:11]
  assign n40_I_3_0_0_1 = n19_O_3_0_0_1; // @[Top.scala 68:11]
  assign n40_I_3_0_0_2 = n19_O_3_0_0_2; // @[Top.scala 68:11]
  assign n40_I_4_0_0_0 = n19_O_4_0_0_0; // @[Top.scala 68:11]
  assign n40_I_4_0_0_1 = n19_O_4_0_0_1; // @[Top.scala 68:11]
  assign n40_I_4_0_0_2 = n19_O_4_0_0_2; // @[Top.scala 68:11]
  assign n40_I_5_0_0_0 = n19_O_5_0_0_0; // @[Top.scala 68:11]
  assign n40_I_5_0_0_1 = n19_O_5_0_0_1; // @[Top.scala 68:11]
  assign n40_I_5_0_0_2 = n19_O_5_0_0_2; // @[Top.scala 68:11]
  assign n40_I_6_0_0_0 = n19_O_6_0_0_0; // @[Top.scala 68:11]
  assign n40_I_6_0_0_1 = n19_O_6_0_0_1; // @[Top.scala 68:11]
  assign n40_I_6_0_0_2 = n19_O_6_0_0_2; // @[Top.scala 68:11]
  assign n40_I_7_0_0_0 = n19_O_7_0_0_0; // @[Top.scala 68:11]
  assign n40_I_7_0_0_1 = n19_O_7_0_0_1; // @[Top.scala 68:11]
  assign n40_I_7_0_0_2 = n19_O_7_0_0_2; // @[Top.scala 68:11]
  assign n41_clock = clock;
  assign n41_valid_up = n2_valid_down; // @[Top.scala 72:18]
  assign n41_I_0_0_0 = n2_O_0_0_0; // @[Top.scala 71:11]
  assign n41_I_1_0_0 = n2_O_1_0_0; // @[Top.scala 71:11]
  assign n41_I_2_0_0 = n2_O_2_0_0; // @[Top.scala 71:11]
  assign n41_I_3_0_0 = n2_O_3_0_0; // @[Top.scala 71:11]
  assign n41_I_4_0_0 = n2_O_4_0_0; // @[Top.scala 71:11]
  assign n41_I_5_0_0 = n2_O_5_0_0; // @[Top.scala 71:11]
  assign n41_I_6_0_0 = n2_O_6_0_0; // @[Top.scala 71:11]
  assign n41_I_7_0_0 = n2_O_7_0_0; // @[Top.scala 71:11]
  assign n42_clock = clock;
  assign n42_valid_up = n41_valid_down; // @[Top.scala 75:18]
  assign n42_I_0_0_0 = n41_O_0_0_0; // @[Top.scala 74:11]
  assign n42_I_1_0_0 = n41_O_1_0_0; // @[Top.scala 74:11]
  assign n42_I_2_0_0 = n41_O_2_0_0; // @[Top.scala 74:11]
  assign n42_I_3_0_0 = n41_O_3_0_0; // @[Top.scala 74:11]
  assign n42_I_4_0_0 = n41_O_4_0_0; // @[Top.scala 74:11]
  assign n42_I_5_0_0 = n41_O_5_0_0; // @[Top.scala 74:11]
  assign n42_I_6_0_0 = n41_O_6_0_0; // @[Top.scala 74:11]
  assign n42_I_7_0_0 = n41_O_7_0_0; // @[Top.scala 74:11]
  assign n43_valid_up = n42_valid_down & n41_valid_down; // @[Top.scala 79:18]
  assign n43_I0_0_0_0 = n42_O_0_0_0; // @[Top.scala 77:12]
  assign n43_I0_1_0_0 = n42_O_1_0_0; // @[Top.scala 77:12]
  assign n43_I0_2_0_0 = n42_O_2_0_0; // @[Top.scala 77:12]
  assign n43_I0_3_0_0 = n42_O_3_0_0; // @[Top.scala 77:12]
  assign n43_I0_4_0_0 = n42_O_4_0_0; // @[Top.scala 77:12]
  assign n43_I0_5_0_0 = n42_O_5_0_0; // @[Top.scala 77:12]
  assign n43_I0_6_0_0 = n42_O_6_0_0; // @[Top.scala 77:12]
  assign n43_I0_7_0_0 = n42_O_7_0_0; // @[Top.scala 77:12]
  assign n43_I1_0_0_0 = n41_O_0_0_0; // @[Top.scala 78:12]
  assign n43_I1_1_0_0 = n41_O_1_0_0; // @[Top.scala 78:12]
  assign n43_I1_2_0_0 = n41_O_2_0_0; // @[Top.scala 78:12]
  assign n43_I1_3_0_0 = n41_O_3_0_0; // @[Top.scala 78:12]
  assign n43_I1_4_0_0 = n41_O_4_0_0; // @[Top.scala 78:12]
  assign n43_I1_5_0_0 = n41_O_5_0_0; // @[Top.scala 78:12]
  assign n43_I1_6_0_0 = n41_O_6_0_0; // @[Top.scala 78:12]
  assign n43_I1_7_0_0 = n41_O_7_0_0; // @[Top.scala 78:12]
  assign n56_valid_up = n43_valid_down & n2_valid_down; // @[Top.scala 83:18]
  assign n56_I0_0_0_0_0 = n43_O_0_0_0_0; // @[Top.scala 81:12]
  assign n56_I0_0_0_0_1 = n43_O_0_0_0_1; // @[Top.scala 81:12]
  assign n56_I0_1_0_0_0 = n43_O_1_0_0_0; // @[Top.scala 81:12]
  assign n56_I0_1_0_0_1 = n43_O_1_0_0_1; // @[Top.scala 81:12]
  assign n56_I0_2_0_0_0 = n43_O_2_0_0_0; // @[Top.scala 81:12]
  assign n56_I0_2_0_0_1 = n43_O_2_0_0_1; // @[Top.scala 81:12]
  assign n56_I0_3_0_0_0 = n43_O_3_0_0_0; // @[Top.scala 81:12]
  assign n56_I0_3_0_0_1 = n43_O_3_0_0_1; // @[Top.scala 81:12]
  assign n56_I0_4_0_0_0 = n43_O_4_0_0_0; // @[Top.scala 81:12]
  assign n56_I0_4_0_0_1 = n43_O_4_0_0_1; // @[Top.scala 81:12]
  assign n56_I0_5_0_0_0 = n43_O_5_0_0_0; // @[Top.scala 81:12]
  assign n56_I0_5_0_0_1 = n43_O_5_0_0_1; // @[Top.scala 81:12]
  assign n56_I0_6_0_0_0 = n43_O_6_0_0_0; // @[Top.scala 81:12]
  assign n56_I0_6_0_0_1 = n43_O_6_0_0_1; // @[Top.scala 81:12]
  assign n56_I0_7_0_0_0 = n43_O_7_0_0_0; // @[Top.scala 81:12]
  assign n56_I0_7_0_0_1 = n43_O_7_0_0_1; // @[Top.scala 81:12]
  assign n56_I1_0_0_0 = n2_O_0_0_0; // @[Top.scala 82:12]
  assign n56_I1_1_0_0 = n2_O_1_0_0; // @[Top.scala 82:12]
  assign n56_I1_2_0_0 = n2_O_2_0_0; // @[Top.scala 82:12]
  assign n56_I1_3_0_0 = n2_O_3_0_0; // @[Top.scala 82:12]
  assign n56_I1_4_0_0 = n2_O_4_0_0; // @[Top.scala 82:12]
  assign n56_I1_5_0_0 = n2_O_5_0_0; // @[Top.scala 82:12]
  assign n56_I1_6_0_0 = n2_O_6_0_0; // @[Top.scala 82:12]
  assign n56_I1_7_0_0 = n2_O_7_0_0; // @[Top.scala 82:12]
  assign n77_valid_up = n56_valid_down; // @[Top.scala 86:18]
  assign n77_I_0_0_0_0 = n56_O_0_0_0_0; // @[Top.scala 85:11]
  assign n77_I_0_0_0_1 = n56_O_0_0_0_1; // @[Top.scala 85:11]
  assign n77_I_0_0_0_2 = n56_O_0_0_0_2; // @[Top.scala 85:11]
  assign n77_I_1_0_0_0 = n56_O_1_0_0_0; // @[Top.scala 85:11]
  assign n77_I_1_0_0_1 = n56_O_1_0_0_1; // @[Top.scala 85:11]
  assign n77_I_1_0_0_2 = n56_O_1_0_0_2; // @[Top.scala 85:11]
  assign n77_I_2_0_0_0 = n56_O_2_0_0_0; // @[Top.scala 85:11]
  assign n77_I_2_0_0_1 = n56_O_2_0_0_1; // @[Top.scala 85:11]
  assign n77_I_2_0_0_2 = n56_O_2_0_0_2; // @[Top.scala 85:11]
  assign n77_I_3_0_0_0 = n56_O_3_0_0_0; // @[Top.scala 85:11]
  assign n77_I_3_0_0_1 = n56_O_3_0_0_1; // @[Top.scala 85:11]
  assign n77_I_3_0_0_2 = n56_O_3_0_0_2; // @[Top.scala 85:11]
  assign n77_I_4_0_0_0 = n56_O_4_0_0_0; // @[Top.scala 85:11]
  assign n77_I_4_0_0_1 = n56_O_4_0_0_1; // @[Top.scala 85:11]
  assign n77_I_4_0_0_2 = n56_O_4_0_0_2; // @[Top.scala 85:11]
  assign n77_I_5_0_0_0 = n56_O_5_0_0_0; // @[Top.scala 85:11]
  assign n77_I_5_0_0_1 = n56_O_5_0_0_1; // @[Top.scala 85:11]
  assign n77_I_5_0_0_2 = n56_O_5_0_0_2; // @[Top.scala 85:11]
  assign n77_I_6_0_0_0 = n56_O_6_0_0_0; // @[Top.scala 85:11]
  assign n77_I_6_0_0_1 = n56_O_6_0_0_1; // @[Top.scala 85:11]
  assign n77_I_6_0_0_2 = n56_O_6_0_0_2; // @[Top.scala 85:11]
  assign n77_I_7_0_0_0 = n56_O_7_0_0_0; // @[Top.scala 85:11]
  assign n77_I_7_0_0_1 = n56_O_7_0_0_1; // @[Top.scala 85:11]
  assign n77_I_7_0_0_2 = n56_O_7_0_0_2; // @[Top.scala 85:11]
  assign n78_valid_up = n40_valid_down & n77_valid_down; // @[Top.scala 90:18]
  assign n78_I0_0_0_0 = n40_O_0_0_0; // @[Top.scala 88:12]
  assign n78_I0_0_0_1 = n40_O_0_0_1; // @[Top.scala 88:12]
  assign n78_I0_0_0_2 = n40_O_0_0_2; // @[Top.scala 88:12]
  assign n78_I0_1_0_0 = n40_O_1_0_0; // @[Top.scala 88:12]
  assign n78_I0_1_0_1 = n40_O_1_0_1; // @[Top.scala 88:12]
  assign n78_I0_1_0_2 = n40_O_1_0_2; // @[Top.scala 88:12]
  assign n78_I0_2_0_0 = n40_O_2_0_0; // @[Top.scala 88:12]
  assign n78_I0_2_0_1 = n40_O_2_0_1; // @[Top.scala 88:12]
  assign n78_I0_2_0_2 = n40_O_2_0_2; // @[Top.scala 88:12]
  assign n78_I0_3_0_0 = n40_O_3_0_0; // @[Top.scala 88:12]
  assign n78_I0_3_0_1 = n40_O_3_0_1; // @[Top.scala 88:12]
  assign n78_I0_3_0_2 = n40_O_3_0_2; // @[Top.scala 88:12]
  assign n78_I0_4_0_0 = n40_O_4_0_0; // @[Top.scala 88:12]
  assign n78_I0_4_0_1 = n40_O_4_0_1; // @[Top.scala 88:12]
  assign n78_I0_4_0_2 = n40_O_4_0_2; // @[Top.scala 88:12]
  assign n78_I0_5_0_0 = n40_O_5_0_0; // @[Top.scala 88:12]
  assign n78_I0_5_0_1 = n40_O_5_0_1; // @[Top.scala 88:12]
  assign n78_I0_5_0_2 = n40_O_5_0_2; // @[Top.scala 88:12]
  assign n78_I0_6_0_0 = n40_O_6_0_0; // @[Top.scala 88:12]
  assign n78_I0_6_0_1 = n40_O_6_0_1; // @[Top.scala 88:12]
  assign n78_I0_6_0_2 = n40_O_6_0_2; // @[Top.scala 88:12]
  assign n78_I0_7_0_0 = n40_O_7_0_0; // @[Top.scala 88:12]
  assign n78_I0_7_0_1 = n40_O_7_0_1; // @[Top.scala 88:12]
  assign n78_I0_7_0_2 = n40_O_7_0_2; // @[Top.scala 88:12]
  assign n78_I1_0_0_0 = n77_O_0_0_0; // @[Top.scala 89:12]
  assign n78_I1_0_0_1 = n77_O_0_0_1; // @[Top.scala 89:12]
  assign n78_I1_0_0_2 = n77_O_0_0_2; // @[Top.scala 89:12]
  assign n78_I1_1_0_0 = n77_O_1_0_0; // @[Top.scala 89:12]
  assign n78_I1_1_0_1 = n77_O_1_0_1; // @[Top.scala 89:12]
  assign n78_I1_1_0_2 = n77_O_1_0_2; // @[Top.scala 89:12]
  assign n78_I1_2_0_0 = n77_O_2_0_0; // @[Top.scala 89:12]
  assign n78_I1_2_0_1 = n77_O_2_0_1; // @[Top.scala 89:12]
  assign n78_I1_2_0_2 = n77_O_2_0_2; // @[Top.scala 89:12]
  assign n78_I1_3_0_0 = n77_O_3_0_0; // @[Top.scala 89:12]
  assign n78_I1_3_0_1 = n77_O_3_0_1; // @[Top.scala 89:12]
  assign n78_I1_3_0_2 = n77_O_3_0_2; // @[Top.scala 89:12]
  assign n78_I1_4_0_0 = n77_O_4_0_0; // @[Top.scala 89:12]
  assign n78_I1_4_0_1 = n77_O_4_0_1; // @[Top.scala 89:12]
  assign n78_I1_4_0_2 = n77_O_4_0_2; // @[Top.scala 89:12]
  assign n78_I1_5_0_0 = n77_O_5_0_0; // @[Top.scala 89:12]
  assign n78_I1_5_0_1 = n77_O_5_0_1; // @[Top.scala 89:12]
  assign n78_I1_5_0_2 = n77_O_5_0_2; // @[Top.scala 89:12]
  assign n78_I1_6_0_0 = n77_O_6_0_0; // @[Top.scala 89:12]
  assign n78_I1_6_0_1 = n77_O_6_0_1; // @[Top.scala 89:12]
  assign n78_I1_6_0_2 = n77_O_6_0_2; // @[Top.scala 89:12]
  assign n78_I1_7_0_0 = n77_O_7_0_0; // @[Top.scala 89:12]
  assign n78_I1_7_0_1 = n77_O_7_0_1; // @[Top.scala 89:12]
  assign n78_I1_7_0_2 = n77_O_7_0_2; // @[Top.scala 89:12]
  assign n88_clock = clock;
  assign n88_valid_up = n1_valid_down; // @[Top.scala 93:18]
  assign n88_I_0_0_0 = n1_O_0_0_0; // @[Top.scala 92:11]
  assign n88_I_1_0_0 = n1_O_1_0_0; // @[Top.scala 92:11]
  assign n88_I_2_0_0 = n1_O_2_0_0; // @[Top.scala 92:11]
  assign n88_I_3_0_0 = n1_O_3_0_0; // @[Top.scala 92:11]
  assign n88_I_4_0_0 = n1_O_4_0_0; // @[Top.scala 92:11]
  assign n88_I_5_0_0 = n1_O_5_0_0; // @[Top.scala 92:11]
  assign n88_I_6_0_0 = n1_O_6_0_0; // @[Top.scala 92:11]
  assign n88_I_7_0_0 = n1_O_7_0_0; // @[Top.scala 92:11]
  assign n89_clock = clock;
  assign n89_valid_up = n88_valid_down; // @[Top.scala 96:18]
  assign n89_I_0_0_0 = n88_O_0_0_0; // @[Top.scala 95:11]
  assign n89_I_1_0_0 = n88_O_1_0_0; // @[Top.scala 95:11]
  assign n89_I_2_0_0 = n88_O_2_0_0; // @[Top.scala 95:11]
  assign n89_I_3_0_0 = n88_O_3_0_0; // @[Top.scala 95:11]
  assign n89_I_4_0_0 = n88_O_4_0_0; // @[Top.scala 95:11]
  assign n89_I_5_0_0 = n88_O_5_0_0; // @[Top.scala 95:11]
  assign n89_I_6_0_0 = n88_O_6_0_0; // @[Top.scala 95:11]
  assign n89_I_7_0_0 = n88_O_7_0_0; // @[Top.scala 95:11]
  assign n90_valid_up = n89_valid_down & n88_valid_down; // @[Top.scala 100:18]
  assign n90_I0_0_0_0 = n89_O_0_0_0; // @[Top.scala 98:12]
  assign n90_I0_1_0_0 = n89_O_1_0_0; // @[Top.scala 98:12]
  assign n90_I0_2_0_0 = n89_O_2_0_0; // @[Top.scala 98:12]
  assign n90_I0_3_0_0 = n89_O_3_0_0; // @[Top.scala 98:12]
  assign n90_I0_4_0_0 = n89_O_4_0_0; // @[Top.scala 98:12]
  assign n90_I0_5_0_0 = n89_O_5_0_0; // @[Top.scala 98:12]
  assign n90_I0_6_0_0 = n89_O_6_0_0; // @[Top.scala 98:12]
  assign n90_I0_7_0_0 = n89_O_7_0_0; // @[Top.scala 98:12]
  assign n90_I1_0_0_0 = n88_O_0_0_0; // @[Top.scala 99:12]
  assign n90_I1_1_0_0 = n88_O_1_0_0; // @[Top.scala 99:12]
  assign n90_I1_2_0_0 = n88_O_2_0_0; // @[Top.scala 99:12]
  assign n90_I1_3_0_0 = n88_O_3_0_0; // @[Top.scala 99:12]
  assign n90_I1_4_0_0 = n88_O_4_0_0; // @[Top.scala 99:12]
  assign n90_I1_5_0_0 = n88_O_5_0_0; // @[Top.scala 99:12]
  assign n90_I1_6_0_0 = n88_O_6_0_0; // @[Top.scala 99:12]
  assign n90_I1_7_0_0 = n88_O_7_0_0; // @[Top.scala 99:12]
  assign n103_valid_up = n90_valid_down & n1_valid_down; // @[Top.scala 104:19]
  assign n103_I0_0_0_0_0 = n90_O_0_0_0_0; // @[Top.scala 102:13]
  assign n103_I0_0_0_0_1 = n90_O_0_0_0_1; // @[Top.scala 102:13]
  assign n103_I0_1_0_0_0 = n90_O_1_0_0_0; // @[Top.scala 102:13]
  assign n103_I0_1_0_0_1 = n90_O_1_0_0_1; // @[Top.scala 102:13]
  assign n103_I0_2_0_0_0 = n90_O_2_0_0_0; // @[Top.scala 102:13]
  assign n103_I0_2_0_0_1 = n90_O_2_0_0_1; // @[Top.scala 102:13]
  assign n103_I0_3_0_0_0 = n90_O_3_0_0_0; // @[Top.scala 102:13]
  assign n103_I0_3_0_0_1 = n90_O_3_0_0_1; // @[Top.scala 102:13]
  assign n103_I0_4_0_0_0 = n90_O_4_0_0_0; // @[Top.scala 102:13]
  assign n103_I0_4_0_0_1 = n90_O_4_0_0_1; // @[Top.scala 102:13]
  assign n103_I0_5_0_0_0 = n90_O_5_0_0_0; // @[Top.scala 102:13]
  assign n103_I0_5_0_0_1 = n90_O_5_0_0_1; // @[Top.scala 102:13]
  assign n103_I0_6_0_0_0 = n90_O_6_0_0_0; // @[Top.scala 102:13]
  assign n103_I0_6_0_0_1 = n90_O_6_0_0_1; // @[Top.scala 102:13]
  assign n103_I0_7_0_0_0 = n90_O_7_0_0_0; // @[Top.scala 102:13]
  assign n103_I0_7_0_0_1 = n90_O_7_0_0_1; // @[Top.scala 102:13]
  assign n103_I1_0_0_0 = n1_O_0_0_0; // @[Top.scala 103:13]
  assign n103_I1_1_0_0 = n1_O_1_0_0; // @[Top.scala 103:13]
  assign n103_I1_2_0_0 = n1_O_2_0_0; // @[Top.scala 103:13]
  assign n103_I1_3_0_0 = n1_O_3_0_0; // @[Top.scala 103:13]
  assign n103_I1_4_0_0 = n1_O_4_0_0; // @[Top.scala 103:13]
  assign n103_I1_5_0_0 = n1_O_5_0_0; // @[Top.scala 103:13]
  assign n103_I1_6_0_0 = n1_O_6_0_0; // @[Top.scala 103:13]
  assign n103_I1_7_0_0 = n1_O_7_0_0; // @[Top.scala 103:13]
  assign n124_valid_up = n103_valid_down; // @[Top.scala 107:19]
  assign n124_I_0_0_0_0 = n103_O_0_0_0_0; // @[Top.scala 106:12]
  assign n124_I_0_0_0_1 = n103_O_0_0_0_1; // @[Top.scala 106:12]
  assign n124_I_0_0_0_2 = n103_O_0_0_0_2; // @[Top.scala 106:12]
  assign n124_I_1_0_0_0 = n103_O_1_0_0_0; // @[Top.scala 106:12]
  assign n124_I_1_0_0_1 = n103_O_1_0_0_1; // @[Top.scala 106:12]
  assign n124_I_1_0_0_2 = n103_O_1_0_0_2; // @[Top.scala 106:12]
  assign n124_I_2_0_0_0 = n103_O_2_0_0_0; // @[Top.scala 106:12]
  assign n124_I_2_0_0_1 = n103_O_2_0_0_1; // @[Top.scala 106:12]
  assign n124_I_2_0_0_2 = n103_O_2_0_0_2; // @[Top.scala 106:12]
  assign n124_I_3_0_0_0 = n103_O_3_0_0_0; // @[Top.scala 106:12]
  assign n124_I_3_0_0_1 = n103_O_3_0_0_1; // @[Top.scala 106:12]
  assign n124_I_3_0_0_2 = n103_O_3_0_0_2; // @[Top.scala 106:12]
  assign n124_I_4_0_0_0 = n103_O_4_0_0_0; // @[Top.scala 106:12]
  assign n124_I_4_0_0_1 = n103_O_4_0_0_1; // @[Top.scala 106:12]
  assign n124_I_4_0_0_2 = n103_O_4_0_0_2; // @[Top.scala 106:12]
  assign n124_I_5_0_0_0 = n103_O_5_0_0_0; // @[Top.scala 106:12]
  assign n124_I_5_0_0_1 = n103_O_5_0_0_1; // @[Top.scala 106:12]
  assign n124_I_5_0_0_2 = n103_O_5_0_0_2; // @[Top.scala 106:12]
  assign n124_I_6_0_0_0 = n103_O_6_0_0_0; // @[Top.scala 106:12]
  assign n124_I_6_0_0_1 = n103_O_6_0_0_1; // @[Top.scala 106:12]
  assign n124_I_6_0_0_2 = n103_O_6_0_0_2; // @[Top.scala 106:12]
  assign n124_I_7_0_0_0 = n103_O_7_0_0_0; // @[Top.scala 106:12]
  assign n124_I_7_0_0_1 = n103_O_7_0_0_1; // @[Top.scala 106:12]
  assign n124_I_7_0_0_2 = n103_O_7_0_0_2; // @[Top.scala 106:12]
  assign n125_valid_up = n78_valid_down & n124_valid_down; // @[Top.scala 111:19]
  assign n125_I0_0_0_0_0 = n78_O_0_0_0_0; // @[Top.scala 109:13]
  assign n125_I0_0_0_0_1 = n78_O_0_0_0_1; // @[Top.scala 109:13]
  assign n125_I0_0_0_0_2 = n78_O_0_0_0_2; // @[Top.scala 109:13]
  assign n125_I0_0_0_1_0 = n78_O_0_0_1_0; // @[Top.scala 109:13]
  assign n125_I0_0_0_1_1 = n78_O_0_0_1_1; // @[Top.scala 109:13]
  assign n125_I0_0_0_1_2 = n78_O_0_0_1_2; // @[Top.scala 109:13]
  assign n125_I0_1_0_0_0 = n78_O_1_0_0_0; // @[Top.scala 109:13]
  assign n125_I0_1_0_0_1 = n78_O_1_0_0_1; // @[Top.scala 109:13]
  assign n125_I0_1_0_0_2 = n78_O_1_0_0_2; // @[Top.scala 109:13]
  assign n125_I0_1_0_1_0 = n78_O_1_0_1_0; // @[Top.scala 109:13]
  assign n125_I0_1_0_1_1 = n78_O_1_0_1_1; // @[Top.scala 109:13]
  assign n125_I0_1_0_1_2 = n78_O_1_0_1_2; // @[Top.scala 109:13]
  assign n125_I0_2_0_0_0 = n78_O_2_0_0_0; // @[Top.scala 109:13]
  assign n125_I0_2_0_0_1 = n78_O_2_0_0_1; // @[Top.scala 109:13]
  assign n125_I0_2_0_0_2 = n78_O_2_0_0_2; // @[Top.scala 109:13]
  assign n125_I0_2_0_1_0 = n78_O_2_0_1_0; // @[Top.scala 109:13]
  assign n125_I0_2_0_1_1 = n78_O_2_0_1_1; // @[Top.scala 109:13]
  assign n125_I0_2_0_1_2 = n78_O_2_0_1_2; // @[Top.scala 109:13]
  assign n125_I0_3_0_0_0 = n78_O_3_0_0_0; // @[Top.scala 109:13]
  assign n125_I0_3_0_0_1 = n78_O_3_0_0_1; // @[Top.scala 109:13]
  assign n125_I0_3_0_0_2 = n78_O_3_0_0_2; // @[Top.scala 109:13]
  assign n125_I0_3_0_1_0 = n78_O_3_0_1_0; // @[Top.scala 109:13]
  assign n125_I0_3_0_1_1 = n78_O_3_0_1_1; // @[Top.scala 109:13]
  assign n125_I0_3_0_1_2 = n78_O_3_0_1_2; // @[Top.scala 109:13]
  assign n125_I0_4_0_0_0 = n78_O_4_0_0_0; // @[Top.scala 109:13]
  assign n125_I0_4_0_0_1 = n78_O_4_0_0_1; // @[Top.scala 109:13]
  assign n125_I0_4_0_0_2 = n78_O_4_0_0_2; // @[Top.scala 109:13]
  assign n125_I0_4_0_1_0 = n78_O_4_0_1_0; // @[Top.scala 109:13]
  assign n125_I0_4_0_1_1 = n78_O_4_0_1_1; // @[Top.scala 109:13]
  assign n125_I0_4_0_1_2 = n78_O_4_0_1_2; // @[Top.scala 109:13]
  assign n125_I0_5_0_0_0 = n78_O_5_0_0_0; // @[Top.scala 109:13]
  assign n125_I0_5_0_0_1 = n78_O_5_0_0_1; // @[Top.scala 109:13]
  assign n125_I0_5_0_0_2 = n78_O_5_0_0_2; // @[Top.scala 109:13]
  assign n125_I0_5_0_1_0 = n78_O_5_0_1_0; // @[Top.scala 109:13]
  assign n125_I0_5_0_1_1 = n78_O_5_0_1_1; // @[Top.scala 109:13]
  assign n125_I0_5_0_1_2 = n78_O_5_0_1_2; // @[Top.scala 109:13]
  assign n125_I0_6_0_0_0 = n78_O_6_0_0_0; // @[Top.scala 109:13]
  assign n125_I0_6_0_0_1 = n78_O_6_0_0_1; // @[Top.scala 109:13]
  assign n125_I0_6_0_0_2 = n78_O_6_0_0_2; // @[Top.scala 109:13]
  assign n125_I0_6_0_1_0 = n78_O_6_0_1_0; // @[Top.scala 109:13]
  assign n125_I0_6_0_1_1 = n78_O_6_0_1_1; // @[Top.scala 109:13]
  assign n125_I0_6_0_1_2 = n78_O_6_0_1_2; // @[Top.scala 109:13]
  assign n125_I0_7_0_0_0 = n78_O_7_0_0_0; // @[Top.scala 109:13]
  assign n125_I0_7_0_0_1 = n78_O_7_0_0_1; // @[Top.scala 109:13]
  assign n125_I0_7_0_0_2 = n78_O_7_0_0_2; // @[Top.scala 109:13]
  assign n125_I0_7_0_1_0 = n78_O_7_0_1_0; // @[Top.scala 109:13]
  assign n125_I0_7_0_1_1 = n78_O_7_0_1_1; // @[Top.scala 109:13]
  assign n125_I0_7_0_1_2 = n78_O_7_0_1_2; // @[Top.scala 109:13]
  assign n125_I1_0_0_0 = n124_O_0_0_0; // @[Top.scala 110:13]
  assign n125_I1_0_0_1 = n124_O_0_0_1; // @[Top.scala 110:13]
  assign n125_I1_0_0_2 = n124_O_0_0_2; // @[Top.scala 110:13]
  assign n125_I1_1_0_0 = n124_O_1_0_0; // @[Top.scala 110:13]
  assign n125_I1_1_0_1 = n124_O_1_0_1; // @[Top.scala 110:13]
  assign n125_I1_1_0_2 = n124_O_1_0_2; // @[Top.scala 110:13]
  assign n125_I1_2_0_0 = n124_O_2_0_0; // @[Top.scala 110:13]
  assign n125_I1_2_0_1 = n124_O_2_0_1; // @[Top.scala 110:13]
  assign n125_I1_2_0_2 = n124_O_2_0_2; // @[Top.scala 110:13]
  assign n125_I1_3_0_0 = n124_O_3_0_0; // @[Top.scala 110:13]
  assign n125_I1_3_0_1 = n124_O_3_0_1; // @[Top.scala 110:13]
  assign n125_I1_3_0_2 = n124_O_3_0_2; // @[Top.scala 110:13]
  assign n125_I1_4_0_0 = n124_O_4_0_0; // @[Top.scala 110:13]
  assign n125_I1_4_0_1 = n124_O_4_0_1; // @[Top.scala 110:13]
  assign n125_I1_4_0_2 = n124_O_4_0_2; // @[Top.scala 110:13]
  assign n125_I1_5_0_0 = n124_O_5_0_0; // @[Top.scala 110:13]
  assign n125_I1_5_0_1 = n124_O_5_0_1; // @[Top.scala 110:13]
  assign n125_I1_5_0_2 = n124_O_5_0_2; // @[Top.scala 110:13]
  assign n125_I1_6_0_0 = n124_O_6_0_0; // @[Top.scala 110:13]
  assign n125_I1_6_0_1 = n124_O_6_0_1; // @[Top.scala 110:13]
  assign n125_I1_6_0_2 = n124_O_6_0_2; // @[Top.scala 110:13]
  assign n125_I1_7_0_0 = n124_O_7_0_0; // @[Top.scala 110:13]
  assign n125_I1_7_0_1 = n124_O_7_0_1; // @[Top.scala 110:13]
  assign n125_I1_7_0_2 = n124_O_7_0_2; // @[Top.scala 110:13]
  assign n141_valid_up = n125_valid_down; // @[Top.scala 114:19]
  assign n141_I_0_0_0_0 = n125_O_0_0_0_0; // @[Top.scala 113:12]
  assign n141_I_0_0_0_1 = n125_O_0_0_0_1; // @[Top.scala 113:12]
  assign n141_I_0_0_0_2 = n125_O_0_0_0_2; // @[Top.scala 113:12]
  assign n141_I_0_0_1_0 = n125_O_0_0_1_0; // @[Top.scala 113:12]
  assign n141_I_0_0_1_1 = n125_O_0_0_1_1; // @[Top.scala 113:12]
  assign n141_I_0_0_1_2 = n125_O_0_0_1_2; // @[Top.scala 113:12]
  assign n141_I_0_0_2_0 = n125_O_0_0_2_0; // @[Top.scala 113:12]
  assign n141_I_0_0_2_1 = n125_O_0_0_2_1; // @[Top.scala 113:12]
  assign n141_I_0_0_2_2 = n125_O_0_0_2_2; // @[Top.scala 113:12]
  assign n141_I_1_0_0_0 = n125_O_1_0_0_0; // @[Top.scala 113:12]
  assign n141_I_1_0_0_1 = n125_O_1_0_0_1; // @[Top.scala 113:12]
  assign n141_I_1_0_0_2 = n125_O_1_0_0_2; // @[Top.scala 113:12]
  assign n141_I_1_0_1_0 = n125_O_1_0_1_0; // @[Top.scala 113:12]
  assign n141_I_1_0_1_1 = n125_O_1_0_1_1; // @[Top.scala 113:12]
  assign n141_I_1_0_1_2 = n125_O_1_0_1_2; // @[Top.scala 113:12]
  assign n141_I_1_0_2_0 = n125_O_1_0_2_0; // @[Top.scala 113:12]
  assign n141_I_1_0_2_1 = n125_O_1_0_2_1; // @[Top.scala 113:12]
  assign n141_I_1_0_2_2 = n125_O_1_0_2_2; // @[Top.scala 113:12]
  assign n141_I_2_0_0_0 = n125_O_2_0_0_0; // @[Top.scala 113:12]
  assign n141_I_2_0_0_1 = n125_O_2_0_0_1; // @[Top.scala 113:12]
  assign n141_I_2_0_0_2 = n125_O_2_0_0_2; // @[Top.scala 113:12]
  assign n141_I_2_0_1_0 = n125_O_2_0_1_0; // @[Top.scala 113:12]
  assign n141_I_2_0_1_1 = n125_O_2_0_1_1; // @[Top.scala 113:12]
  assign n141_I_2_0_1_2 = n125_O_2_0_1_2; // @[Top.scala 113:12]
  assign n141_I_2_0_2_0 = n125_O_2_0_2_0; // @[Top.scala 113:12]
  assign n141_I_2_0_2_1 = n125_O_2_0_2_1; // @[Top.scala 113:12]
  assign n141_I_2_0_2_2 = n125_O_2_0_2_2; // @[Top.scala 113:12]
  assign n141_I_3_0_0_0 = n125_O_3_0_0_0; // @[Top.scala 113:12]
  assign n141_I_3_0_0_1 = n125_O_3_0_0_1; // @[Top.scala 113:12]
  assign n141_I_3_0_0_2 = n125_O_3_0_0_2; // @[Top.scala 113:12]
  assign n141_I_3_0_1_0 = n125_O_3_0_1_0; // @[Top.scala 113:12]
  assign n141_I_3_0_1_1 = n125_O_3_0_1_1; // @[Top.scala 113:12]
  assign n141_I_3_0_1_2 = n125_O_3_0_1_2; // @[Top.scala 113:12]
  assign n141_I_3_0_2_0 = n125_O_3_0_2_0; // @[Top.scala 113:12]
  assign n141_I_3_0_2_1 = n125_O_3_0_2_1; // @[Top.scala 113:12]
  assign n141_I_3_0_2_2 = n125_O_3_0_2_2; // @[Top.scala 113:12]
  assign n141_I_4_0_0_0 = n125_O_4_0_0_0; // @[Top.scala 113:12]
  assign n141_I_4_0_0_1 = n125_O_4_0_0_1; // @[Top.scala 113:12]
  assign n141_I_4_0_0_2 = n125_O_4_0_0_2; // @[Top.scala 113:12]
  assign n141_I_4_0_1_0 = n125_O_4_0_1_0; // @[Top.scala 113:12]
  assign n141_I_4_0_1_1 = n125_O_4_0_1_1; // @[Top.scala 113:12]
  assign n141_I_4_0_1_2 = n125_O_4_0_1_2; // @[Top.scala 113:12]
  assign n141_I_4_0_2_0 = n125_O_4_0_2_0; // @[Top.scala 113:12]
  assign n141_I_4_0_2_1 = n125_O_4_0_2_1; // @[Top.scala 113:12]
  assign n141_I_4_0_2_2 = n125_O_4_0_2_2; // @[Top.scala 113:12]
  assign n141_I_5_0_0_0 = n125_O_5_0_0_0; // @[Top.scala 113:12]
  assign n141_I_5_0_0_1 = n125_O_5_0_0_1; // @[Top.scala 113:12]
  assign n141_I_5_0_0_2 = n125_O_5_0_0_2; // @[Top.scala 113:12]
  assign n141_I_5_0_1_0 = n125_O_5_0_1_0; // @[Top.scala 113:12]
  assign n141_I_5_0_1_1 = n125_O_5_0_1_1; // @[Top.scala 113:12]
  assign n141_I_5_0_1_2 = n125_O_5_0_1_2; // @[Top.scala 113:12]
  assign n141_I_5_0_2_0 = n125_O_5_0_2_0; // @[Top.scala 113:12]
  assign n141_I_5_0_2_1 = n125_O_5_0_2_1; // @[Top.scala 113:12]
  assign n141_I_5_0_2_2 = n125_O_5_0_2_2; // @[Top.scala 113:12]
  assign n141_I_6_0_0_0 = n125_O_6_0_0_0; // @[Top.scala 113:12]
  assign n141_I_6_0_0_1 = n125_O_6_0_0_1; // @[Top.scala 113:12]
  assign n141_I_6_0_0_2 = n125_O_6_0_0_2; // @[Top.scala 113:12]
  assign n141_I_6_0_1_0 = n125_O_6_0_1_0; // @[Top.scala 113:12]
  assign n141_I_6_0_1_1 = n125_O_6_0_1_1; // @[Top.scala 113:12]
  assign n141_I_6_0_1_2 = n125_O_6_0_1_2; // @[Top.scala 113:12]
  assign n141_I_6_0_2_0 = n125_O_6_0_2_0; // @[Top.scala 113:12]
  assign n141_I_6_0_2_1 = n125_O_6_0_2_1; // @[Top.scala 113:12]
  assign n141_I_6_0_2_2 = n125_O_6_0_2_2; // @[Top.scala 113:12]
  assign n141_I_7_0_0_0 = n125_O_7_0_0_0; // @[Top.scala 113:12]
  assign n141_I_7_0_0_1 = n125_O_7_0_0_1; // @[Top.scala 113:12]
  assign n141_I_7_0_0_2 = n125_O_7_0_0_2; // @[Top.scala 113:12]
  assign n141_I_7_0_1_0 = n125_O_7_0_1_0; // @[Top.scala 113:12]
  assign n141_I_7_0_1_1 = n125_O_7_0_1_1; // @[Top.scala 113:12]
  assign n141_I_7_0_1_2 = n125_O_7_0_1_2; // @[Top.scala 113:12]
  assign n141_I_7_0_2_0 = n125_O_7_0_2_0; // @[Top.scala 113:12]
  assign n141_I_7_0_2_1 = n125_O_7_0_2_1; // @[Top.scala 113:12]
  assign n141_I_7_0_2_2 = n125_O_7_0_2_2; // @[Top.scala 113:12]
  assign n183_clock = clock;
  assign n183_reset = reset;
  assign n183_valid_up = n141_valid_down; // @[Top.scala 117:19]
  assign n183_I_0_0_0 = n141_O_0_0_0; // @[Top.scala 116:12]
  assign n183_I_0_0_1 = n141_O_0_0_1; // @[Top.scala 116:12]
  assign n183_I_0_0_2 = n141_O_0_0_2; // @[Top.scala 116:12]
  assign n183_I_0_1_0 = n141_O_0_1_0; // @[Top.scala 116:12]
  assign n183_I_0_1_1 = n141_O_0_1_1; // @[Top.scala 116:12]
  assign n183_I_0_1_2 = n141_O_0_1_2; // @[Top.scala 116:12]
  assign n183_I_0_2_0 = n141_O_0_2_0; // @[Top.scala 116:12]
  assign n183_I_0_2_1 = n141_O_0_2_1; // @[Top.scala 116:12]
  assign n183_I_0_2_2 = n141_O_0_2_2; // @[Top.scala 116:12]
  assign n183_I_1_0_0 = n141_O_1_0_0; // @[Top.scala 116:12]
  assign n183_I_1_0_1 = n141_O_1_0_1; // @[Top.scala 116:12]
  assign n183_I_1_0_2 = n141_O_1_0_2; // @[Top.scala 116:12]
  assign n183_I_1_1_0 = n141_O_1_1_0; // @[Top.scala 116:12]
  assign n183_I_1_1_1 = n141_O_1_1_1; // @[Top.scala 116:12]
  assign n183_I_1_1_2 = n141_O_1_1_2; // @[Top.scala 116:12]
  assign n183_I_1_2_0 = n141_O_1_2_0; // @[Top.scala 116:12]
  assign n183_I_1_2_1 = n141_O_1_2_1; // @[Top.scala 116:12]
  assign n183_I_1_2_2 = n141_O_1_2_2; // @[Top.scala 116:12]
  assign n183_I_2_0_0 = n141_O_2_0_0; // @[Top.scala 116:12]
  assign n183_I_2_0_1 = n141_O_2_0_1; // @[Top.scala 116:12]
  assign n183_I_2_0_2 = n141_O_2_0_2; // @[Top.scala 116:12]
  assign n183_I_2_1_0 = n141_O_2_1_0; // @[Top.scala 116:12]
  assign n183_I_2_1_1 = n141_O_2_1_1; // @[Top.scala 116:12]
  assign n183_I_2_1_2 = n141_O_2_1_2; // @[Top.scala 116:12]
  assign n183_I_2_2_0 = n141_O_2_2_0; // @[Top.scala 116:12]
  assign n183_I_2_2_1 = n141_O_2_2_1; // @[Top.scala 116:12]
  assign n183_I_2_2_2 = n141_O_2_2_2; // @[Top.scala 116:12]
  assign n183_I_3_0_0 = n141_O_3_0_0; // @[Top.scala 116:12]
  assign n183_I_3_0_1 = n141_O_3_0_1; // @[Top.scala 116:12]
  assign n183_I_3_0_2 = n141_O_3_0_2; // @[Top.scala 116:12]
  assign n183_I_3_1_0 = n141_O_3_1_0; // @[Top.scala 116:12]
  assign n183_I_3_1_1 = n141_O_3_1_1; // @[Top.scala 116:12]
  assign n183_I_3_1_2 = n141_O_3_1_2; // @[Top.scala 116:12]
  assign n183_I_3_2_0 = n141_O_3_2_0; // @[Top.scala 116:12]
  assign n183_I_3_2_1 = n141_O_3_2_1; // @[Top.scala 116:12]
  assign n183_I_3_2_2 = n141_O_3_2_2; // @[Top.scala 116:12]
  assign n183_I_4_0_0 = n141_O_4_0_0; // @[Top.scala 116:12]
  assign n183_I_4_0_1 = n141_O_4_0_1; // @[Top.scala 116:12]
  assign n183_I_4_0_2 = n141_O_4_0_2; // @[Top.scala 116:12]
  assign n183_I_4_1_0 = n141_O_4_1_0; // @[Top.scala 116:12]
  assign n183_I_4_1_1 = n141_O_4_1_1; // @[Top.scala 116:12]
  assign n183_I_4_1_2 = n141_O_4_1_2; // @[Top.scala 116:12]
  assign n183_I_4_2_0 = n141_O_4_2_0; // @[Top.scala 116:12]
  assign n183_I_4_2_1 = n141_O_4_2_1; // @[Top.scala 116:12]
  assign n183_I_4_2_2 = n141_O_4_2_2; // @[Top.scala 116:12]
  assign n183_I_5_0_0 = n141_O_5_0_0; // @[Top.scala 116:12]
  assign n183_I_5_0_1 = n141_O_5_0_1; // @[Top.scala 116:12]
  assign n183_I_5_0_2 = n141_O_5_0_2; // @[Top.scala 116:12]
  assign n183_I_5_1_0 = n141_O_5_1_0; // @[Top.scala 116:12]
  assign n183_I_5_1_1 = n141_O_5_1_1; // @[Top.scala 116:12]
  assign n183_I_5_1_2 = n141_O_5_1_2; // @[Top.scala 116:12]
  assign n183_I_5_2_0 = n141_O_5_2_0; // @[Top.scala 116:12]
  assign n183_I_5_2_1 = n141_O_5_2_1; // @[Top.scala 116:12]
  assign n183_I_5_2_2 = n141_O_5_2_2; // @[Top.scala 116:12]
  assign n183_I_6_0_0 = n141_O_6_0_0; // @[Top.scala 116:12]
  assign n183_I_6_0_1 = n141_O_6_0_1; // @[Top.scala 116:12]
  assign n183_I_6_0_2 = n141_O_6_0_2; // @[Top.scala 116:12]
  assign n183_I_6_1_0 = n141_O_6_1_0; // @[Top.scala 116:12]
  assign n183_I_6_1_1 = n141_O_6_1_1; // @[Top.scala 116:12]
  assign n183_I_6_1_2 = n141_O_6_1_2; // @[Top.scala 116:12]
  assign n183_I_6_2_0 = n141_O_6_2_0; // @[Top.scala 116:12]
  assign n183_I_6_2_1 = n141_O_6_2_1; // @[Top.scala 116:12]
  assign n183_I_6_2_2 = n141_O_6_2_2; // @[Top.scala 116:12]
  assign n183_I_7_0_0 = n141_O_7_0_0; // @[Top.scala 116:12]
  assign n183_I_7_0_1 = n141_O_7_0_1; // @[Top.scala 116:12]
  assign n183_I_7_0_2 = n141_O_7_0_2; // @[Top.scala 116:12]
  assign n183_I_7_1_0 = n141_O_7_1_0; // @[Top.scala 116:12]
  assign n183_I_7_1_1 = n141_O_7_1_1; // @[Top.scala 116:12]
  assign n183_I_7_1_2 = n141_O_7_1_2; // @[Top.scala 116:12]
  assign n183_I_7_2_0 = n141_O_7_2_0; // @[Top.scala 116:12]
  assign n183_I_7_2_1 = n141_O_7_2_1; // @[Top.scala 116:12]
  assign n183_I_7_2_2 = n141_O_7_2_2; // @[Top.scala 116:12]
  assign n184_clock = clock;
  assign n184_valid_up = n183_valid_down; // @[Top.scala 120:19]
  assign n184_I_0_0_0 = n183_O_0_0_0; // @[Top.scala 119:12]
  assign n184_I_1_0_0 = n183_O_1_0_0; // @[Top.scala 119:12]
  assign n184_I_2_0_0 = n183_O_2_0_0; // @[Top.scala 119:12]
  assign n184_I_3_0_0 = n183_O_3_0_0; // @[Top.scala 119:12]
  assign n184_I_4_0_0 = n183_O_4_0_0; // @[Top.scala 119:12]
  assign n184_I_5_0_0 = n183_O_5_0_0; // @[Top.scala 119:12]
  assign n184_I_6_0_0 = n183_O_6_0_0; // @[Top.scala 119:12]
  assign n184_I_7_0_0 = n183_O_7_0_0; // @[Top.scala 119:12]
  assign n185_clock = clock;
  assign n185_valid_up = n184_valid_down; // @[Top.scala 123:19]
  assign n185_I_0_0_0 = n184_O_0_0_0; // @[Top.scala 122:12]
  assign n185_I_1_0_0 = n184_O_1_0_0; // @[Top.scala 122:12]
  assign n185_I_2_0_0 = n184_O_2_0_0; // @[Top.scala 122:12]
  assign n185_I_3_0_0 = n184_O_3_0_0; // @[Top.scala 122:12]
  assign n185_I_4_0_0 = n184_O_4_0_0; // @[Top.scala 122:12]
  assign n185_I_5_0_0 = n184_O_5_0_0; // @[Top.scala 122:12]
  assign n185_I_6_0_0 = n184_O_6_0_0; // @[Top.scala 122:12]
  assign n185_I_7_0_0 = n184_O_7_0_0; // @[Top.scala 122:12]
  assign n186_clock = clock;
  assign n186_valid_up = n185_valid_down; // @[Top.scala 126:19]
  assign n186_I_0_0_0 = n185_O_0_0_0; // @[Top.scala 125:12]
  assign n186_I_1_0_0 = n185_O_1_0_0; // @[Top.scala 125:12]
  assign n186_I_2_0_0 = n185_O_2_0_0; // @[Top.scala 125:12]
  assign n186_I_3_0_0 = n185_O_3_0_0; // @[Top.scala 125:12]
  assign n186_I_4_0_0 = n185_O_4_0_0; // @[Top.scala 125:12]
  assign n186_I_5_0_0 = n185_O_5_0_0; // @[Top.scala 125:12]
  assign n186_I_6_0_0 = n185_O_6_0_0; // @[Top.scala 125:12]
  assign n186_I_7_0_0 = n185_O_7_0_0; // @[Top.scala 125:12]
endmodule
