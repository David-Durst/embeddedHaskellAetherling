// Latency = 4
module top(
  input CLK/*verilator public*/, 
  input [7:0] I_0_0_0/*verilator public*/, 
  output [7:0] O_0_0_0/*verilator public*/, 
  input [7:0] I_1_0_0/*verilator public*/, 
  output [7:0] O_1_0_0/*verilator public*/, 
  input [7:0] I_2_0_0/*verilator public*/, 
  output [7:0] O_2_0_0/*verilator public*/, 
  input [7:0] I_3_0_0/*verilator public*/, 
  output [7:0] O_3_0_0/*verilator public*/, 
  input [7:0] I_4_0_0/*verilator public*/, 
  output [7:0] O_4_0_0/*verilator public*/, 
  input [7:0] I_5_0_0/*verilator public*/, 
  output [7:0] O_5_0_0/*verilator public*/, 
  input [7:0] I_6_0_0/*verilator public*/, 
  output [7:0] O_6_0_0/*verilator public*/, 
  input [7:0] I_7_0_0/*verilator public*/, 
  output [7:0] O_7_0_0/*verilator public*/, 
  output valid_down/*verilator public*/, 
  input valid_up/*verilator public*/
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(CLK), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x511_TREADY(dontcare), // @[:@1298.4]
    .io_in_x511_TDATA({I_0_0_0,I_1_0_0,I_2_0_0,I_3_0_0,I_4_0_0,I_5_0_0,I_6_0_0,I_7_0_0}), // @[:@1298.4]
    .io_in_x511_TID(8'h0),
    .io_in_x511_TDEST(8'h0),
    .io_in_x512_TVALID(valid_down), // @[:@1298.4]
    .io_in_x512_TDATA({O_0_0_0,O_1_0_0,O_2_0_0,O_3_0_0,O_4_0_0,O_5_0_0,O_6_0_0,O_7_0_0}), // @[:@1298.4]
    .io_in_x512_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x519_ctrchain cchain ( // @[:@2879.2]
    .clock(CLK), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule



module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@104.4]
  wire  _T_57; // @[Counter.scala 285:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@118.4]
  FF bases_0 ( // @[Counter.scala 253:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh1d); // @[Counter.scala 285:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh1d); // @[Counter.scala 325:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 276:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 256:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_133 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = io_rst | done_0_io_output; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = done_0_io_output & _T_166; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module x996_outr_UnitPipe_sm( // @[:@2389.2]
  input   clock, // @[:@2390.4]
  input   reset, // @[:@2391.4]
  input   io_enable, // @[:@2392.4]
  output  io_done, // @[:@2392.4]
  input   io_parentAck, // @[:@2392.4]
  input   io_doneIn_0, // @[:@2392.4]
  output  io_enableOut_0, // @[:@2392.4]
  output  io_childAck_0, // @[:@2392.4]
  input   io_ctrCopyDone_0 // @[:@2392.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@2395.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@2398.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@2415.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2532.4]
  wire  _T_105; // @[Controllers.scala 165:35:@2430.4]
  wire  _T_107; // @[Controllers.scala 165:60:@2431.4]
  wire  _T_108; // @[Controllers.scala 165:58:@2432.4]
  wire  _T_110; // @[Controllers.scala 165:76:@2433.4]
  wire  _T_111; // @[Controllers.scala 165:74:@2434.4]
  wire  _T_115; // @[Controllers.scala 165:109:@2437.4]
  wire  _T_118; // @[Controllers.scala 165:141:@2439.4]
  wire  _T_126; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  wire  _T_130; // @[Controllers.scala 167:54:@2454.4]
  wire  _T_131; // @[Controllers.scala 167:52:@2455.4]
  wire  _T_138; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  wire  _T_156; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  wire  _T_160; // @[Controllers.scala 169:67:@2486.4]
  wire  _T_161; // @[Controllers.scala 169:86:@2487.4]
  wire  _T_174; // @[Controllers.scala 213:68:@2501.4]
  wire  _T_176; // @[Controllers.scala 213:90:@2503.4]
  wire  _T_178; // @[Controllers.scala 213:132:@2505.4]
  reg  _T_186; // @[package.scala 48:56:@2511.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@2513.4]
  reg  _T_200; // @[package.scala 48:56:@2529.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@2395.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@2398.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@2415.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2446.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2460.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2478.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2515.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2532.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@2430.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@2431.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@2432.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@2433.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@2434.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@2437.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@2439.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@2454.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@2455.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@2486.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@2487.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@2501.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@2503.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@2505.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@2513.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@2539.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@2509.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@2500.4]
  assign active_0_clock = clock; // @[:@2396.4]
  assign active_0_reset = reset; // @[:@2397.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@2441.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@2445.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@2403.4]
  assign done_0_clock = clock; // @[:@2399.4]
  assign done_0_reset = reset; // @[:@2400.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@2491.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@2413.4 Controllers.scala 170:32:@2498.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@2404.4]
  assign iterDone_0_clock = clock; // @[:@2416.4]
  assign iterDone_0_reset = reset; // @[:@2417.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@2459.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@2427.4 Controllers.scala 168:36:@2475.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@2418.4]
  assign RetimeWrapper_clock = clock; // @[:@2447.4]
  assign RetimeWrapper_reset = reset; // @[:@2448.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2450.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@2449.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2461.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2462.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2464.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@2463.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2479.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2480.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2482.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@2481.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2516.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2517.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2519.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@2518.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2533.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2534.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@2536.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@2535.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module SingleCounter_1( // @[:@2659.2]
  input         clock, // @[:@2660.4]
  input         reset, // @[:@2661.4]
  input         io_input_reset, // @[:@2662.4]
  input         io_input_enable, // @[:@2662.4]
  output [31:0] io_output_count_0, // @[:@2662.4]
  output        io_output_oobs_0, // @[:@2662.4]
  output        io_output_done, // @[:@2662.4]
  output        io_output_saturated // @[:@2662.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2675.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2675.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2691.4]
  wire  _T_36; // @[Counter.scala 256:45:@2694.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@2719.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@2720.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@2721.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@2722.4]
  wire  _T_57; // @[Counter.scala 285:18:@2724.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@2732.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@2735.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@2736.4]
  wire  _T_75; // @[Counter.scala 314:102:@2740.4]
  wire  _T_77; // @[Counter.scala 314:130:@2741.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2675.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2691.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2694.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2719.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh2); // @[Counter.scala 283:33:@2720.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh2); // @[Counter.scala 283:33:@2721.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2722.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@2724.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2732.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2735.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@2736.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2740.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh4); // @[Counter.scala 314:130:@2741.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2739.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2743.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2745.4]
  assign io_output_saturated = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 332:25:@2748.4]
  assign bases_0_clock = clock; // @[:@2676.4]
  assign bases_0_reset = reset; // @[:@2677.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2738.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2717.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2718.4]
  assign SRFF_clock = clock; // @[:@2692.4]
  assign SRFF_reset = reset; // @[:@2693.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2696.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2698.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2699.4]
endmodule
module SingleCounter_2( // @[:@2788.2]
  input         clock, // @[:@2789.4]
  input         reset, // @[:@2790.4]
  input         io_setup_saturate, // @[:@2791.4]
  input         io_input_reset, // @[:@2791.4]
  input         io_input_enable, // @[:@2791.4]
  output [31:0] io_output_count_0, // @[:@2791.4]
  output        io_output_oobs_0, // @[:@2791.4]
  output        io_output_done // @[:@2791.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2804.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2804.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2804.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2820.4]
  wire  _T_36; // @[Counter.scala 256:45:@2823.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@2848.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@2849.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@2850.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@2851.4]
  wire  _T_57; // @[Counter.scala 285:18:@2853.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@2861.4]
  wire [31:0] _T_70; // @[Counter.scala 291:85:@2863.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@2864.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@2865.4]
  wire  _T_75; // @[Counter.scala 314:102:@2869.4]
  wire  _T_77; // @[Counter.scala 314:130:@2870.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2804.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2820.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2823.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2848.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh4); // @[Counter.scala 283:33:@2849.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh4); // @[Counter.scala 283:33:@2850.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2851.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@2853.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2861.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 32'h0; // @[Counter.scala 291:85:@2863.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2864.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 291:74:@2865.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2869.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh4); // @[Counter.scala 314:130:@2870.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2868.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2872.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2874.4]
  assign bases_0_clock = clock; // @[:@2805.4]
  assign bases_0_reset = reset; // @[:@2806.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2867.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2846.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2847.4]
  assign SRFF_clock = clock; // @[:@2821.4]
  assign SRFF_reset = reset; // @[:@2822.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2825.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2827.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2828.4]
endmodule
module x519_ctrchain( // @[:@2879.2]
  input         clock, // @[:@2880.4]
  input         reset, // @[:@2881.4]
  input         io_input_reset, // @[:@2882.4]
  input         io_input_enable, // @[:@2882.4]
  output [31:0] io_output_counts_1, // @[:@2882.4]
  output [31:0] io_output_counts_0, // @[:@2882.4]
  output        io_output_oobs_0, // @[:@2882.4]
  output        io_output_oobs_1, // @[:@2882.4]
  output        io_output_done // @[:@2882.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 505:46:@2884.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_1_clock; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 505:46:@2887.4]
  wire [31:0] ctrs_1_io_output_count_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 505:46:@2887.4]
  wire  isDone; // @[Counter.scala 533:51:@2904.4]
  reg  wasDone; // @[Counter.scala 534:24:@2905.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 538:69:@2913.4]
  wire  _T_66; // @[Counter.scala 538:80:@2914.4]
  reg  doneLatch; // @[Counter.scala 542:26:@2919.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 543:48:@2920.4]
  wire  _T_74; // @[Counter.scala 543:19:@2921.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 505:46:@2884.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 505:46:@2887.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 533:51:@2904.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 538:69:@2913.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 538:80:@2914.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 543:48:@2920.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 543:19:@2921.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 549:32:@2926.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 549:32:@2923.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2925.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2928.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 538:18:@2916.4]
  assign ctrs_0_clock = clock; // @[:@2885.4]
  assign ctrs_0_reset = reset; // @[:@2886.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2893.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 518:29:@2900.4]
  assign ctrs_1_clock = clock; // @[:@2888.4]
  assign ctrs_1_reset = reset; // @[:@2889.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 524:31:@2903.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2897.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 516:33:@2898.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_12( // @[:@2968.2]
  input   clock, // @[:@2969.4]
  input   reset, // @[:@2970.4]
  input   io_flow, // @[:@2971.4]
  input   io_in, // @[:@2971.4]
  output  io_out // @[:@2971.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(52)) sr ( // @[RetimeShiftRegister.scala 15:20:@2973.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2986.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2985.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2984.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2983.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2982.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2980.4]
endmodule
module RetimeWrapper_16( // @[:@3096.2]
  input   clock, // @[:@3097.4]
  input   reset, // @[:@3098.4]
  input   io_flow, // @[:@3099.4]
  input   io_in, // @[:@3099.4]
  output  io_out // @[:@3099.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(51)) sr ( // @[RetimeShiftRegister.scala 15:20:@3101.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3114.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3113.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3112.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3111.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3110.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3108.4]
endmodule
module x995_inr_Foreach_SAMPLER_BOX_sm( // @[:@3116.2]
  input   clock, // @[:@3117.4]
  input   reset, // @[:@3118.4]
  input   io_enable, // @[:@3119.4]
  output  io_done, // @[:@3119.4]
  output  io_doneLatch, // @[:@3119.4]
  input   io_ctrDone, // @[:@3119.4]
  output  io_datapathEn, // @[:@3119.4]
  output  io_ctrInc, // @[:@3119.4]
  output  io_ctrRst, // @[:@3119.4]
  input   io_parentAck, // @[:@3119.4]
  input   io_backpressure, // @[:@3119.4]
  input   io_break // @[:@3119.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3121.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3121.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3124.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3124.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3216.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3129.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3130.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3131.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3132.4]
  wire  _T_100; // @[package.scala 100:49:@3149.4]
  reg  _T_103; // @[package.scala 48:56:@3150.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  wire  _T_110; // @[package.scala 100:49:@3165.4]
  reg  _T_113; // @[package.scala 48:56:@3166.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3168.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3173.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3174.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3177.4]
  wire  _T_124; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  wire  _T_126; // @[package.scala 100:49:@3187.4]
  reg  _T_129; // @[package.scala 48:56:@3188.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3210.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3212.4]
  reg  _T_153; // @[package.scala 48:56:@3213.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3223.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3224.4]
  SRFF active ( // @[Controllers.scala 261:22:@3121.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3124.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_12 RetimeWrapper ( // @[package.scala 93:22:@3158.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_1 ( // @[package.scala 93:22:@3180.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3192.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3200.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_4 ( // @[package.scala 93:22:@3216.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3129.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3130.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3131.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3132.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3149.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3165.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3168.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3173.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3174.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3177.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3187.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3212.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3223.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3224.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3191.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3226.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3176.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3179.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3171.4]
  assign active_clock = clock; // @[:@3122.4]
  assign active_reset = reset; // @[:@3123.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3134.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3138.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3139.4]
  assign done_clock = clock; // @[:@3125.4]
  assign done_reset = reset; // @[:@3126.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3154.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3147.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3148.4]
  assign RetimeWrapper_clock = clock; // @[:@3159.4]
  assign RetimeWrapper_reset = reset; // @[:@3160.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3162.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3161.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3181.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3182.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3184.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3183.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3193.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3194.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3196.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3195.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3201.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3202.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3204.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3203.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3217.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3218.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3220.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3219.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3332.2]
  input  [31:0] io_a, // @[:@3335.4]
  output [31:0] io_b // @[:@3335.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3345.4]
endmodule
module _( // @[:@3347.2]
  input  [31:0] io_b, // @[:@3350.4]
  output [31:0] io_result // @[:@3350.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3355.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3355.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3355.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3368.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3363.4]
endmodule
module RetimeWrapper_21( // @[:@3452.2]
  input        clock, // @[:@3453.4]
  input        reset, // @[:@3454.4]
  input        io_flow, // @[:@3455.4]
  input  [7:0] io_in, // @[:@3455.4]
  output [7:0] io_out // @[:@3455.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3457.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3470.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3469.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@3468.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3467.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3466.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3464.4]
endmodule
module Mem1D_4( // @[:@3472.2]
  input        clock, // @[:@3473.4]
  input        reset, // @[:@3474.4]
  input        io_r_ofs_0, // @[:@3475.4]
  input        io_r_backpressure, // @[:@3475.4]
  input        io_w_ofs_0, // @[:@3475.4]
  input  [7:0] io_w_data_0, // @[:@3475.4]
  input        io_w_en_0, // @[:@3475.4]
  output [7:0] io_output // @[:@3475.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@3494.4]
  reg [7:0] _T_127; // @[MemPrimitives.scala 560:26:@3479.4]
  reg [31:0] _RAND_0;
  wire  _T_130; // @[MemPrimitives.scala 561:61:@3481.4]
  wire  _T_131; // @[MemPrimitives.scala 561:44:@3482.4]
  wire [7:0] _T_132; // @[MemPrimitives.scala 561:19:@3483.4]
  wire  _T_135; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  wire  _T_137; // @[Mux.scala 46:19:@3492.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@3485.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3494.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_130 = io_w_ofs_0 == 1'h0; // @[MemPrimitives.scala 561:61:@3481.4]
  assign _T_131 = io_w_en_0 & _T_130; // @[MemPrimitives.scala 561:44:@3482.4]
  assign _T_132 = _T_131 ? io_w_data_0 : _T_127; // @[MemPrimitives.scala 561:19:@3483.4]
  assign _T_135 = RetimeWrapper_io_out; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  assign _T_137 = 1'h0 == _T_135; // @[Mux.scala 46:19:@3492.4]
  assign io_output = RetimeWrapper_1_io_out; // @[MemPrimitives.scala 565:17:@3501.4]
  assign RetimeWrapper_clock = clock; // @[:@3486.4]
  assign RetimeWrapper_reset = reset; // @[:@3487.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@3489.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@3488.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3495.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3496.4]
  assign RetimeWrapper_1_io_flow = io_r_backpressure; // @[package.scala 95:18:@3498.4]
  assign RetimeWrapper_1_io_in = _T_137 ? _T_127 : 8'h0; // @[package.scala 94:16:@3497.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_127 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_127 <= 8'h0;
    end else begin
      if (_T_131) begin
        _T_127 <= io_w_data_0;
      end
    end
  end
endmodule
module StickySelects( // @[:@4928.2]
  input   clock, // @[:@4929.4]
  input   reset, // @[:@4930.4]
  input   io_ins_0, // @[:@4931.4]
  input   io_ins_1, // @[:@4931.4]
  input   io_ins_2, // @[:@4931.4]
  input   io_ins_3, // @[:@4931.4]
  output  io_outs_0, // @[:@4931.4]
  output  io_outs_1, // @[:@4931.4]
  output  io_outs_2, // @[:@4931.4]
  output  io_outs_3 // @[:@4931.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@4933.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@4934.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@4935.4]
  wire  _T_23; // @[StickySelects.scala 24:52:@4936.4]
  wire  _T_24; // @[StickySelects.scala 24:21:@4937.4]
  reg  _T_27; // @[StickySelects.scala 21:22:@4939.4]
  reg [31:0] _RAND_1;
  wire  _T_28; // @[StickySelects.scala 22:54:@4940.4]
  wire  _T_29; // @[StickySelects.scala 22:54:@4941.4]
  wire  _T_31; // @[StickySelects.scala 24:52:@4942.4]
  wire  _T_32; // @[StickySelects.scala 24:21:@4943.4]
  reg  _T_35; // @[StickySelects.scala 21:22:@4945.4]
  reg [31:0] _RAND_2;
  wire  _T_36; // @[StickySelects.scala 22:54:@4946.4]
  wire  _T_37; // @[StickySelects.scala 22:54:@4947.4]
  wire  _T_39; // @[StickySelects.scala 24:52:@4948.4]
  wire  _T_40; // @[StickySelects.scala 24:21:@4949.4]
  reg  _T_43; // @[StickySelects.scala 21:22:@4951.4]
  reg [31:0] _RAND_3;
  wire  _T_45; // @[StickySelects.scala 22:54:@4953.4]
  wire  _T_47; // @[StickySelects.scala 24:52:@4954.4]
  wire  _T_48; // @[StickySelects.scala 24:21:@4955.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@4934.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@4935.4]
  assign _T_23 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@4936.4]
  assign _T_24 = _T_21 ? 1'h0 : _T_23; // @[StickySelects.scala 24:21:@4937.4]
  assign _T_28 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@4940.4]
  assign _T_29 = _T_28 | io_ins_3; // @[StickySelects.scala 22:54:@4941.4]
  assign _T_31 = io_ins_1 | _T_27; // @[StickySelects.scala 24:52:@4942.4]
  assign _T_32 = _T_29 ? 1'h0 : _T_31; // @[StickySelects.scala 24:21:@4943.4]
  assign _T_36 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@4946.4]
  assign _T_37 = _T_36 | io_ins_3; // @[StickySelects.scala 22:54:@4947.4]
  assign _T_39 = io_ins_2 | _T_35; // @[StickySelects.scala 24:52:@4948.4]
  assign _T_40 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 24:21:@4949.4]
  assign _T_45 = _T_36 | io_ins_2; // @[StickySelects.scala 22:54:@4953.4]
  assign _T_47 = io_ins_3 | _T_43; // @[StickySelects.scala 24:52:@4954.4]
  assign _T_48 = _T_45 ? 1'h0 : _T_47; // @[StickySelects.scala 24:21:@4955.4]
  assign io_outs_0 = _T_21 ? 1'h0 : _T_23; // @[StickySelects.scala 28:52:@4957.4]
  assign io_outs_1 = _T_29 ? 1'h0 : _T_31; // @[StickySelects.scala 28:52:@4958.4]
  assign io_outs_2 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 28:52:@4959.4]
  assign io_outs_3 = _T_45 ? 1'h0 : _T_47; // @[StickySelects.scala 28:52:@4960.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_27 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_35 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_43 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_21) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_23;
      end
    end
    if (reset) begin
      _T_27 <= 1'h0;
    end else begin
      if (_T_29) begin
        _T_27 <= 1'h0;
      end else begin
        _T_27 <= _T_31;
      end
    end
    if (reset) begin
      _T_35 <= 1'h0;
    end else begin
      if (_T_37) begin
        _T_35 <= 1'h0;
      end else begin
        _T_35 <= _T_39;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_45) begin
        _T_43 <= 1'h0;
      end else begin
        _T_43 <= _T_47;
      end
    end
  end
endmodule
module StickySelects_2( // @[:@4996.2]
  input   clock, // @[:@4997.4]
  input   reset, // @[:@4998.4]
  input   io_ins_0, // @[:@4999.4]
  input   io_ins_1, // @[:@4999.4]
  input   io_ins_2, // @[:@4999.4]
  input   io_ins_3, // @[:@4999.4]
  input   io_ins_4, // @[:@4999.4]
  input   io_ins_5, // @[:@4999.4]
  input   io_ins_6, // @[:@4999.4]
  input   io_ins_7, // @[:@4999.4]
  output  io_outs_0, // @[:@4999.4]
  output  io_outs_1, // @[:@4999.4]
  output  io_outs_2, // @[:@4999.4]
  output  io_outs_3, // @[:@4999.4]
  output  io_outs_4, // @[:@4999.4]
  output  io_outs_5, // @[:@4999.4]
  output  io_outs_6, // @[:@4999.4]
  output  io_outs_7 // @[:@4999.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@5001.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@5002.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@5003.4]
  wire  _T_22; // @[StickySelects.scala 22:54:@5004.4]
  wire  _T_23; // @[StickySelects.scala 22:54:@5005.4]
  wire  _T_24; // @[StickySelects.scala 22:54:@5006.4]
  wire  _T_25; // @[StickySelects.scala 22:54:@5007.4]
  wire  _T_27; // @[StickySelects.scala 24:52:@5008.4]
  wire  _T_28; // @[StickySelects.scala 24:21:@5009.4]
  reg  _T_31; // @[StickySelects.scala 21:22:@5011.4]
  reg [31:0] _RAND_1;
  wire  _T_32; // @[StickySelects.scala 22:54:@5012.4]
  wire  _T_33; // @[StickySelects.scala 22:54:@5013.4]
  wire  _T_34; // @[StickySelects.scala 22:54:@5014.4]
  wire  _T_35; // @[StickySelects.scala 22:54:@5015.4]
  wire  _T_36; // @[StickySelects.scala 22:54:@5016.4]
  wire  _T_37; // @[StickySelects.scala 22:54:@5017.4]
  wire  _T_39; // @[StickySelects.scala 24:52:@5018.4]
  wire  _T_40; // @[StickySelects.scala 24:21:@5019.4]
  reg  _T_43; // @[StickySelects.scala 21:22:@5021.4]
  reg [31:0] _RAND_2;
  wire  _T_44; // @[StickySelects.scala 22:54:@5022.4]
  wire  _T_45; // @[StickySelects.scala 22:54:@5023.4]
  wire  _T_46; // @[StickySelects.scala 22:54:@5024.4]
  wire  _T_47; // @[StickySelects.scala 22:54:@5025.4]
  wire  _T_48; // @[StickySelects.scala 22:54:@5026.4]
  wire  _T_49; // @[StickySelects.scala 22:54:@5027.4]
  wire  _T_51; // @[StickySelects.scala 24:52:@5028.4]
  wire  _T_52; // @[StickySelects.scala 24:21:@5029.4]
  reg  _T_55; // @[StickySelects.scala 21:22:@5031.4]
  reg [31:0] _RAND_3;
  wire  _T_57; // @[StickySelects.scala 22:54:@5033.4]
  wire  _T_58; // @[StickySelects.scala 22:54:@5034.4]
  wire  _T_59; // @[StickySelects.scala 22:54:@5035.4]
  wire  _T_60; // @[StickySelects.scala 22:54:@5036.4]
  wire  _T_61; // @[StickySelects.scala 22:54:@5037.4]
  wire  _T_63; // @[StickySelects.scala 24:52:@5038.4]
  wire  _T_64; // @[StickySelects.scala 24:21:@5039.4]
  reg  _T_67; // @[StickySelects.scala 21:22:@5041.4]
  reg [31:0] _RAND_4;
  wire  _T_70; // @[StickySelects.scala 22:54:@5044.4]
  wire  _T_71; // @[StickySelects.scala 22:54:@5045.4]
  wire  _T_72; // @[StickySelects.scala 22:54:@5046.4]
  wire  _T_73; // @[StickySelects.scala 22:54:@5047.4]
  wire  _T_75; // @[StickySelects.scala 24:52:@5048.4]
  wire  _T_76; // @[StickySelects.scala 24:21:@5049.4]
  reg  _T_79; // @[StickySelects.scala 21:22:@5051.4]
  reg [31:0] _RAND_5;
  wire  _T_83; // @[StickySelects.scala 22:54:@5055.4]
  wire  _T_84; // @[StickySelects.scala 22:54:@5056.4]
  wire  _T_85; // @[StickySelects.scala 22:54:@5057.4]
  wire  _T_87; // @[StickySelects.scala 24:52:@5058.4]
  wire  _T_88; // @[StickySelects.scala 24:21:@5059.4]
  reg  _T_91; // @[StickySelects.scala 21:22:@5061.4]
  reg [31:0] _RAND_6;
  wire  _T_96; // @[StickySelects.scala 22:54:@5066.4]
  wire  _T_97; // @[StickySelects.scala 22:54:@5067.4]
  wire  _T_99; // @[StickySelects.scala 24:52:@5068.4]
  wire  _T_100; // @[StickySelects.scala 24:21:@5069.4]
  reg  _T_103; // @[StickySelects.scala 21:22:@5071.4]
  reg [31:0] _RAND_7;
  wire  _T_109; // @[StickySelects.scala 22:54:@5077.4]
  wire  _T_111; // @[StickySelects.scala 24:52:@5078.4]
  wire  _T_112; // @[StickySelects.scala 24:21:@5079.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@5002.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@5003.4]
  assign _T_22 = _T_21 | io_ins_4; // @[StickySelects.scala 22:54:@5004.4]
  assign _T_23 = _T_22 | io_ins_5; // @[StickySelects.scala 22:54:@5005.4]
  assign _T_24 = _T_23 | io_ins_6; // @[StickySelects.scala 22:54:@5006.4]
  assign _T_25 = _T_24 | io_ins_7; // @[StickySelects.scala 22:54:@5007.4]
  assign _T_27 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@5008.4]
  assign _T_28 = _T_25 ? 1'h0 : _T_27; // @[StickySelects.scala 24:21:@5009.4]
  assign _T_32 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@5012.4]
  assign _T_33 = _T_32 | io_ins_3; // @[StickySelects.scala 22:54:@5013.4]
  assign _T_34 = _T_33 | io_ins_4; // @[StickySelects.scala 22:54:@5014.4]
  assign _T_35 = _T_34 | io_ins_5; // @[StickySelects.scala 22:54:@5015.4]
  assign _T_36 = _T_35 | io_ins_6; // @[StickySelects.scala 22:54:@5016.4]
  assign _T_37 = _T_36 | io_ins_7; // @[StickySelects.scala 22:54:@5017.4]
  assign _T_39 = io_ins_1 | _T_31; // @[StickySelects.scala 24:52:@5018.4]
  assign _T_40 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 24:21:@5019.4]
  assign _T_44 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@5022.4]
  assign _T_45 = _T_44 | io_ins_3; // @[StickySelects.scala 22:54:@5023.4]
  assign _T_46 = _T_45 | io_ins_4; // @[StickySelects.scala 22:54:@5024.4]
  assign _T_47 = _T_46 | io_ins_5; // @[StickySelects.scala 22:54:@5025.4]
  assign _T_48 = _T_47 | io_ins_6; // @[StickySelects.scala 22:54:@5026.4]
  assign _T_49 = _T_48 | io_ins_7; // @[StickySelects.scala 22:54:@5027.4]
  assign _T_51 = io_ins_2 | _T_43; // @[StickySelects.scala 24:52:@5028.4]
  assign _T_52 = _T_49 ? 1'h0 : _T_51; // @[StickySelects.scala 24:21:@5029.4]
  assign _T_57 = _T_44 | io_ins_2; // @[StickySelects.scala 22:54:@5033.4]
  assign _T_58 = _T_57 | io_ins_4; // @[StickySelects.scala 22:54:@5034.4]
  assign _T_59 = _T_58 | io_ins_5; // @[StickySelects.scala 22:54:@5035.4]
  assign _T_60 = _T_59 | io_ins_6; // @[StickySelects.scala 22:54:@5036.4]
  assign _T_61 = _T_60 | io_ins_7; // @[StickySelects.scala 22:54:@5037.4]
  assign _T_63 = io_ins_3 | _T_55; // @[StickySelects.scala 24:52:@5038.4]
  assign _T_64 = _T_61 ? 1'h0 : _T_63; // @[StickySelects.scala 24:21:@5039.4]
  assign _T_70 = _T_57 | io_ins_3; // @[StickySelects.scala 22:54:@5044.4]
  assign _T_71 = _T_70 | io_ins_5; // @[StickySelects.scala 22:54:@5045.4]
  assign _T_72 = _T_71 | io_ins_6; // @[StickySelects.scala 22:54:@5046.4]
  assign _T_73 = _T_72 | io_ins_7; // @[StickySelects.scala 22:54:@5047.4]
  assign _T_75 = io_ins_4 | _T_67; // @[StickySelects.scala 24:52:@5048.4]
  assign _T_76 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 24:21:@5049.4]
  assign _T_83 = _T_70 | io_ins_4; // @[StickySelects.scala 22:54:@5055.4]
  assign _T_84 = _T_83 | io_ins_6; // @[StickySelects.scala 22:54:@5056.4]
  assign _T_85 = _T_84 | io_ins_7; // @[StickySelects.scala 22:54:@5057.4]
  assign _T_87 = io_ins_5 | _T_79; // @[StickySelects.scala 24:52:@5058.4]
  assign _T_88 = _T_85 ? 1'h0 : _T_87; // @[StickySelects.scala 24:21:@5059.4]
  assign _T_96 = _T_83 | io_ins_5; // @[StickySelects.scala 22:54:@5066.4]
  assign _T_97 = _T_96 | io_ins_7; // @[StickySelects.scala 22:54:@5067.4]
  assign _T_99 = io_ins_6 | _T_91; // @[StickySelects.scala 24:52:@5068.4]
  assign _T_100 = _T_97 ? 1'h0 : _T_99; // @[StickySelects.scala 24:21:@5069.4]
  assign _T_109 = _T_96 | io_ins_6; // @[StickySelects.scala 22:54:@5077.4]
  assign _T_111 = io_ins_7 | _T_103; // @[StickySelects.scala 24:52:@5078.4]
  assign _T_112 = _T_109 ? 1'h0 : _T_111; // @[StickySelects.scala 24:21:@5079.4]
  assign io_outs_0 = _T_25 ? 1'h0 : _T_27; // @[StickySelects.scala 28:52:@5081.4]
  assign io_outs_1 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 28:52:@5082.4]
  assign io_outs_2 = _T_49 ? 1'h0 : _T_51; // @[StickySelects.scala 28:52:@5083.4]
  assign io_outs_3 = _T_61 ? 1'h0 : _T_63; // @[StickySelects.scala 28:52:@5084.4]
  assign io_outs_4 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 28:52:@5085.4]
  assign io_outs_5 = _T_85 ? 1'h0 : _T_87; // @[StickySelects.scala 28:52:@5086.4]
  assign io_outs_6 = _T_97 ? 1'h0 : _T_99; // @[StickySelects.scala 28:52:@5087.4]
  assign io_outs_7 = _T_109 ? 1'h0 : _T_111; // @[StickySelects.scala 28:52:@5088.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_31 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_43 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_55 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_67 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_79 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_91 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_103 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_25) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_27;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_37) begin
        _T_31 <= 1'h0;
      end else begin
        _T_31 <= _T_39;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_49) begin
        _T_43 <= 1'h0;
      end else begin
        _T_43 <= _T_51;
      end
    end
    if (reset) begin
      _T_55 <= 1'h0;
    end else begin
      if (_T_61) begin
        _T_55 <= 1'h0;
      end else begin
        _T_55 <= _T_63;
      end
    end
    if (reset) begin
      _T_67 <= 1'h0;
    end else begin
      if (_T_73) begin
        _T_67 <= 1'h0;
      end else begin
        _T_67 <= _T_75;
      end
    end
    if (reset) begin
      _T_79 <= 1'h0;
    end else begin
      if (_T_85) begin
        _T_79 <= 1'h0;
      end else begin
        _T_79 <= _T_87;
      end
    end
    if (reset) begin
      _T_91 <= 1'h0;
    end else begin
      if (_T_97) begin
        _T_91 <= 1'h0;
      end else begin
        _T_91 <= _T_99;
      end
    end
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      if (_T_109) begin
        _T_103 <= 1'h0;
      end else begin
        _T_103 <= _T_111;
      end
    end
  end
endmodule
module RetimeWrapper_52( // @[:@5964.2]
  input   clock, // @[:@5965.4]
  input   reset, // @[:@5966.4]
  input   io_flow, // @[:@5967.4]
  input   io_in, // @[:@5967.4]
  output  io_out // @[:@5967.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@5969.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@5982.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@5981.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@5980.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@5979.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@5978.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@5976.4]
endmodule
module x524_lb_0( // @[:@9024.2]
  input        clock, // @[:@9025.4]
  input        reset, // @[:@9026.4]
  input  [2:0] io_rPort_23_banks_0, // @[:@9027.4]
  input        io_rPort_23_ofs_0, // @[:@9027.4]
  input        io_rPort_23_en_0, // @[:@9027.4]
  input        io_rPort_23_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_23_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_22_banks_0, // @[:@9027.4]
  input        io_rPort_22_ofs_0, // @[:@9027.4]
  input        io_rPort_22_en_0, // @[:@9027.4]
  input        io_rPort_22_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_22_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_21_banks_0, // @[:@9027.4]
  input        io_rPort_21_ofs_0, // @[:@9027.4]
  input        io_rPort_21_en_0, // @[:@9027.4]
  input        io_rPort_21_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_21_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_20_banks_0, // @[:@9027.4]
  input        io_rPort_20_ofs_0, // @[:@9027.4]
  input        io_rPort_20_en_0, // @[:@9027.4]
  input        io_rPort_20_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_20_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_19_banks_0, // @[:@9027.4]
  input        io_rPort_19_ofs_0, // @[:@9027.4]
  input        io_rPort_19_en_0, // @[:@9027.4]
  input        io_rPort_19_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_19_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_18_banks_0, // @[:@9027.4]
  input        io_rPort_18_ofs_0, // @[:@9027.4]
  input        io_rPort_18_en_0, // @[:@9027.4]
  input        io_rPort_18_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_18_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_17_banks_0, // @[:@9027.4]
  input        io_rPort_17_ofs_0, // @[:@9027.4]
  input        io_rPort_17_en_0, // @[:@9027.4]
  input        io_rPort_17_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_17_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_16_banks_0, // @[:@9027.4]
  input        io_rPort_16_ofs_0, // @[:@9027.4]
  input        io_rPort_16_en_0, // @[:@9027.4]
  input        io_rPort_16_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_16_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_15_banks_0, // @[:@9027.4]
  input        io_rPort_15_ofs_0, // @[:@9027.4]
  input        io_rPort_15_en_0, // @[:@9027.4]
  input        io_rPort_15_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_15_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_14_banks_0, // @[:@9027.4]
  input        io_rPort_14_ofs_0, // @[:@9027.4]
  input        io_rPort_14_en_0, // @[:@9027.4]
  input        io_rPort_14_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_14_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_13_banks_0, // @[:@9027.4]
  input        io_rPort_13_ofs_0, // @[:@9027.4]
  input        io_rPort_13_en_0, // @[:@9027.4]
  input        io_rPort_13_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_13_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_12_banks_0, // @[:@9027.4]
  input        io_rPort_12_ofs_0, // @[:@9027.4]
  input        io_rPort_12_en_0, // @[:@9027.4]
  input        io_rPort_12_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_12_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_11_banks_0, // @[:@9027.4]
  input        io_rPort_11_ofs_0, // @[:@9027.4]
  input        io_rPort_11_en_0, // @[:@9027.4]
  input        io_rPort_11_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_11_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_10_banks_0, // @[:@9027.4]
  input        io_rPort_10_ofs_0, // @[:@9027.4]
  input        io_rPort_10_en_0, // @[:@9027.4]
  input        io_rPort_10_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_10_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_9_banks_0, // @[:@9027.4]
  input        io_rPort_9_ofs_0, // @[:@9027.4]
  input        io_rPort_9_en_0, // @[:@9027.4]
  input        io_rPort_9_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_9_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@9027.4]
  input        io_rPort_8_ofs_0, // @[:@9027.4]
  input        io_rPort_8_en_0, // @[:@9027.4]
  input        io_rPort_8_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_8_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@9027.4]
  input        io_rPort_7_ofs_0, // @[:@9027.4]
  input        io_rPort_7_en_0, // @[:@9027.4]
  input        io_rPort_7_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_7_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@9027.4]
  input        io_rPort_6_ofs_0, // @[:@9027.4]
  input        io_rPort_6_en_0, // @[:@9027.4]
  input        io_rPort_6_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_6_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@9027.4]
  input        io_rPort_5_ofs_0, // @[:@9027.4]
  input        io_rPort_5_en_0, // @[:@9027.4]
  input        io_rPort_5_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_5_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@9027.4]
  input        io_rPort_4_ofs_0, // @[:@9027.4]
  input        io_rPort_4_en_0, // @[:@9027.4]
  input        io_rPort_4_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_4_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@9027.4]
  input        io_rPort_3_ofs_0, // @[:@9027.4]
  input        io_rPort_3_en_0, // @[:@9027.4]
  input        io_rPort_3_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_3_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@9027.4]
  input        io_rPort_2_ofs_0, // @[:@9027.4]
  input        io_rPort_2_en_0, // @[:@9027.4]
  input        io_rPort_2_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_2_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@9027.4]
  input        io_rPort_1_ofs_0, // @[:@9027.4]
  input        io_rPort_1_en_0, // @[:@9027.4]
  input        io_rPort_1_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_1_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@9027.4]
  input        io_rPort_0_ofs_0, // @[:@9027.4]
  input        io_rPort_0_en_0, // @[:@9027.4]
  input        io_rPort_0_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_0_output_0, // @[:@9027.4]
  input  [2:0] io_wPort_7_banks_0, // @[:@9027.4]
  input        io_wPort_7_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_7_data_0, // @[:@9027.4]
  input        io_wPort_7_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_6_banks_0, // @[:@9027.4]
  input        io_wPort_6_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_6_data_0, // @[:@9027.4]
  input        io_wPort_6_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_5_banks_0, // @[:@9027.4]
  input        io_wPort_5_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_5_data_0, // @[:@9027.4]
  input        io_wPort_5_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_4_banks_0, // @[:@9027.4]
  input        io_wPort_4_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_4_data_0, // @[:@9027.4]
  input        io_wPort_4_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_3_banks_0, // @[:@9027.4]
  input        io_wPort_3_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_3_data_0, // @[:@9027.4]
  input        io_wPort_3_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_2_banks_0, // @[:@9027.4]
  input        io_wPort_2_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_2_data_0, // @[:@9027.4]
  input        io_wPort_2_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_1_banks_0, // @[:@9027.4]
  input        io_wPort_1_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_1_data_0, // @[:@9027.4]
  input        io_wPort_1_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@9027.4]
  input        io_wPort_0_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_0_data_0, // @[:@9027.4]
  input        io_wPort_0_en_0 // @[:@9027.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9238.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@9238.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9254.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@9254.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9270.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@9270.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9286.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@9286.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9302.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@9302.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9318.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@9318.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9334.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@9334.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9350.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@9350.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9366.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@9366.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9382.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@9382.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9398.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@9398.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9414.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@9414.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9430.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@9430.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9446.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@9446.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9462.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@9462.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9478.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@9478.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_6; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_7; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_6; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_7; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_6; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_7; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_6; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_7; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@10675.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@10675.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@10675.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@10675.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@10675.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@10683.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@10683.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@10683.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@10683.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@10683.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@10691.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@10691.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@10691.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@10691.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@10691.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@10699.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@10699.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@10699.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@10699.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@10699.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@10723.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@10723.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@10723.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@10723.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@10723.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@10731.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@10731.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@10731.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@10731.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@10731.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@10739.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@10739.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@10739.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@10739.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@10739.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@10771.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@10771.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@10771.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@10771.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@10771.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@10779.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@10779.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@10779.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@10779.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@10779.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@10787.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@10787.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@10787.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@10787.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@10787.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@10795.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@10795.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@10795.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@10795.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@10795.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@10819.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@10819.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@10819.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@10819.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@10819.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@10827.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@10827.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@10827.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@10827.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@10827.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@10835.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@10835.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@10835.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@10835.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@10835.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@10843.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@10843.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@10843.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@10843.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@10843.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@10867.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@10867.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@10867.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@10867.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@10867.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@10875.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@10875.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@10875.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@10875.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@10875.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@10883.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@10883.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@10883.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@10883.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@10883.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@10891.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@10891.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@10891.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@10891.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@10891.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@10915.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@10915.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@10915.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@10915.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@10915.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@10923.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@10923.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@10923.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@10923.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@10923.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@10931.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@10931.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@10931.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@10931.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@10931.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@10939.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@10939.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@10939.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@10939.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@10939.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@10963.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@10963.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@10963.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@10963.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@10963.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@10971.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@10971.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@10971.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@10971.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@10971.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@10979.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@10979.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@10979.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@10979.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@10979.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@10987.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@10987.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@10987.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@10987.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@10987.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@11011.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@11011.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@11011.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@11011.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@11011.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@11019.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@11019.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@11019.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@11019.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@11019.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@11027.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@11027.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@11027.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@11027.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@11027.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@11035.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@11035.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@11035.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@11035.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@11035.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@11059.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@11059.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@11059.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@11059.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@11059.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@11067.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@11067.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@11067.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@11067.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@11067.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@11075.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@11075.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@11075.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@11075.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@11075.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@11083.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@11083.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@11083.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@11083.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@11083.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@11107.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@11107.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@11107.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@11107.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@11107.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@11115.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@11115.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@11115.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@11115.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@11115.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@11123.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@11123.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@11123.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@11123.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@11123.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@11131.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@11131.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@11131.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@11131.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@11131.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@11155.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@11155.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@11155.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@11155.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@11155.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@11163.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@11163.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@11163.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@11163.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@11163.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@11171.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@11171.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@11171.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@11171.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@11171.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@11203.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@11203.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@11203.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@11203.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@11203.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@11211.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@11211.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@11211.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@11211.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@11211.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@11219.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@11219.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@11219.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@11219.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@11219.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@11227.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@11227.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@11227.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@11227.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@11227.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@11251.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@11251.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@11251.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@11251.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@11251.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@11259.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@11259.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@11259.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@11259.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@11259.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@11267.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@11267.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@11267.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@11267.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@11267.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@11275.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@11275.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@11275.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@11275.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@11275.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@11299.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@11299.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@11299.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@11299.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@11299.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@11307.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@11307.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@11307.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@11307.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@11307.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@11315.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@11315.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@11315.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@11315.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@11315.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@11323.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@11323.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@11323.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@11323.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@11323.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@11347.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@11347.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@11347.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@11347.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@11347.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@11355.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@11355.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@11355.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@11355.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@11355.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@11363.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@11363.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@11363.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@11363.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@11363.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@11371.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@11371.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@11371.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@11371.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@11371.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@11395.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@11395.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@11395.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@11395.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@11395.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@11403.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@11403.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@11403.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@11403.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@11403.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@11411.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@11411.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@11411.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@11411.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@11411.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@11419.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@11419.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@11419.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@11419.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@11419.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@11443.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@11443.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@11443.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@11443.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@11443.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@11451.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@11451.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@11451.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@11451.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@11451.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@11459.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@11459.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@11459.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@11459.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@11459.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@11467.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@11467.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@11467.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@11467.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@11467.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@11491.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@11491.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@11491.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@11491.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@11491.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@11499.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@11499.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@11499.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@11499.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@11499.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@11507.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@11507.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@11507.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@11507.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@11507.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@11515.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@11515.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@11515.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@11515.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@11515.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@11539.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@11539.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@11539.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@11539.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@11539.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@11547.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@11547.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@11547.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@11547.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@11547.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@11555.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@11555.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@11555.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@11555.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@11555.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@11563.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@11563.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@11563.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@11563.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@11563.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@11587.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@11587.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@11587.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@11587.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@11587.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@11595.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@11595.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@11595.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@11595.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@11595.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@11603.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@11603.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@11603.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@11603.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@11603.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@11611.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@11611.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@11611.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@11611.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@11611.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@11635.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@11635.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@11635.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@11635.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@11635.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@11643.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@11643.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@11643.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@11643.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@11643.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@11651.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@11651.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@11651.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@11651.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@11651.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@11659.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@11659.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@11659.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@11659.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@11659.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@11683.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@11683.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@11683.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@11683.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@11683.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@11691.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@11691.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@11691.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@11691.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@11691.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@11699.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@11699.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@11699.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@11699.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@11699.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@11707.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@11707.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@11707.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@11707.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@11707.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@11731.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@11731.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@11731.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@11731.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@11731.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@11739.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@11739.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@11739.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@11739.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@11739.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@11747.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@11747.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@11747.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@11747.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@11747.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@11755.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@11755.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@11755.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@11755.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@11755.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@11779.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@11779.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@11779.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@11779.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@11779.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@11787.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@11787.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@11787.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@11787.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@11787.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@11795.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@11795.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@11795.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@11795.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@11795.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@11803.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@11803.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@11803.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@11803.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@11803.4]
  wire  _T_1032; // @[MemPrimitives.scala 82:210:@9494.4]
  wire  _T_1035; // @[MemPrimitives.scala 83:102:@9496.4]
  wire  _T_1037; // @[MemPrimitives.scala 82:210:@9497.4]
  wire  _T_1040; // @[MemPrimitives.scala 83:102:@9499.4]
  wire [9:0] _T_1042; // @[Cat.scala 30:58:@9501.4]
  wire [9:0] _T_1044; // @[Cat.scala 30:58:@9503.4]
  wire [9:0] _T_1045; // @[Mux.scala 31:69:@9504.4]
  wire  _T_1050; // @[MemPrimitives.scala 82:210:@9511.4]
  wire  _T_1053; // @[MemPrimitives.scala 83:102:@9513.4]
  wire  _T_1055; // @[MemPrimitives.scala 82:210:@9514.4]
  wire  _T_1058; // @[MemPrimitives.scala 83:102:@9516.4]
  wire [9:0] _T_1060; // @[Cat.scala 30:58:@9518.4]
  wire [9:0] _T_1062; // @[Cat.scala 30:58:@9520.4]
  wire [9:0] _T_1063; // @[Mux.scala 31:69:@9521.4]
  wire  _T_1068; // @[MemPrimitives.scala 82:210:@9528.4]
  wire  _T_1071; // @[MemPrimitives.scala 83:102:@9530.4]
  wire  _T_1073; // @[MemPrimitives.scala 82:210:@9531.4]
  wire  _T_1076; // @[MemPrimitives.scala 83:102:@9533.4]
  wire [9:0] _T_1078; // @[Cat.scala 30:58:@9535.4]
  wire [9:0] _T_1080; // @[Cat.scala 30:58:@9537.4]
  wire [9:0] _T_1081; // @[Mux.scala 31:69:@9538.4]
  wire  _T_1086; // @[MemPrimitives.scala 82:210:@9545.4]
  wire  _T_1089; // @[MemPrimitives.scala 83:102:@9547.4]
  wire  _T_1091; // @[MemPrimitives.scala 82:210:@9548.4]
  wire  _T_1094; // @[MemPrimitives.scala 83:102:@9550.4]
  wire [9:0] _T_1096; // @[Cat.scala 30:58:@9552.4]
  wire [9:0] _T_1098; // @[Cat.scala 30:58:@9554.4]
  wire [9:0] _T_1099; // @[Mux.scala 31:69:@9555.4]
  wire  _T_1104; // @[MemPrimitives.scala 82:210:@9562.4]
  wire  _T_1107; // @[MemPrimitives.scala 83:102:@9564.4]
  wire  _T_1109; // @[MemPrimitives.scala 82:210:@9565.4]
  wire  _T_1112; // @[MemPrimitives.scala 83:102:@9567.4]
  wire [9:0] _T_1114; // @[Cat.scala 30:58:@9569.4]
  wire [9:0] _T_1116; // @[Cat.scala 30:58:@9571.4]
  wire [9:0] _T_1117; // @[Mux.scala 31:69:@9572.4]
  wire  _T_1122; // @[MemPrimitives.scala 82:210:@9579.4]
  wire  _T_1125; // @[MemPrimitives.scala 83:102:@9581.4]
  wire  _T_1127; // @[MemPrimitives.scala 82:210:@9582.4]
  wire  _T_1130; // @[MemPrimitives.scala 83:102:@9584.4]
  wire [9:0] _T_1132; // @[Cat.scala 30:58:@9586.4]
  wire [9:0] _T_1134; // @[Cat.scala 30:58:@9588.4]
  wire [9:0] _T_1135; // @[Mux.scala 31:69:@9589.4]
  wire  _T_1140; // @[MemPrimitives.scala 82:210:@9596.4]
  wire  _T_1143; // @[MemPrimitives.scala 83:102:@9598.4]
  wire  _T_1145; // @[MemPrimitives.scala 82:210:@9599.4]
  wire  _T_1148; // @[MemPrimitives.scala 83:102:@9601.4]
  wire [9:0] _T_1150; // @[Cat.scala 30:58:@9603.4]
  wire [9:0] _T_1152; // @[Cat.scala 30:58:@9605.4]
  wire [9:0] _T_1153; // @[Mux.scala 31:69:@9606.4]
  wire  _T_1158; // @[MemPrimitives.scala 82:210:@9613.4]
  wire  _T_1161; // @[MemPrimitives.scala 83:102:@9615.4]
  wire  _T_1163; // @[MemPrimitives.scala 82:210:@9616.4]
  wire  _T_1166; // @[MemPrimitives.scala 83:102:@9618.4]
  wire [9:0] _T_1168; // @[Cat.scala 30:58:@9620.4]
  wire [9:0] _T_1170; // @[Cat.scala 30:58:@9622.4]
  wire [9:0] _T_1171; // @[Mux.scala 31:69:@9623.4]
  wire  _T_1176; // @[MemPrimitives.scala 82:210:@9630.4]
  wire  _T_1179; // @[MemPrimitives.scala 83:102:@9632.4]
  wire  _T_1181; // @[MemPrimitives.scala 82:210:@9633.4]
  wire  _T_1184; // @[MemPrimitives.scala 83:102:@9635.4]
  wire [9:0] _T_1186; // @[Cat.scala 30:58:@9637.4]
  wire [9:0] _T_1188; // @[Cat.scala 30:58:@9639.4]
  wire [9:0] _T_1189; // @[Mux.scala 31:69:@9640.4]
  wire  _T_1194; // @[MemPrimitives.scala 82:210:@9647.4]
  wire  _T_1197; // @[MemPrimitives.scala 83:102:@9649.4]
  wire  _T_1199; // @[MemPrimitives.scala 82:210:@9650.4]
  wire  _T_1202; // @[MemPrimitives.scala 83:102:@9652.4]
  wire [9:0] _T_1204; // @[Cat.scala 30:58:@9654.4]
  wire [9:0] _T_1206; // @[Cat.scala 30:58:@9656.4]
  wire [9:0] _T_1207; // @[Mux.scala 31:69:@9657.4]
  wire  _T_1212; // @[MemPrimitives.scala 82:210:@9664.4]
  wire  _T_1215; // @[MemPrimitives.scala 83:102:@9666.4]
  wire  _T_1217; // @[MemPrimitives.scala 82:210:@9667.4]
  wire  _T_1220; // @[MemPrimitives.scala 83:102:@9669.4]
  wire [9:0] _T_1222; // @[Cat.scala 30:58:@9671.4]
  wire [9:0] _T_1224; // @[Cat.scala 30:58:@9673.4]
  wire [9:0] _T_1225; // @[Mux.scala 31:69:@9674.4]
  wire  _T_1230; // @[MemPrimitives.scala 82:210:@9681.4]
  wire  _T_1233; // @[MemPrimitives.scala 83:102:@9683.4]
  wire  _T_1235; // @[MemPrimitives.scala 82:210:@9684.4]
  wire  _T_1238; // @[MemPrimitives.scala 83:102:@9686.4]
  wire [9:0] _T_1240; // @[Cat.scala 30:58:@9688.4]
  wire [9:0] _T_1242; // @[Cat.scala 30:58:@9690.4]
  wire [9:0] _T_1243; // @[Mux.scala 31:69:@9691.4]
  wire  _T_1248; // @[MemPrimitives.scala 82:210:@9698.4]
  wire  _T_1251; // @[MemPrimitives.scala 83:102:@9700.4]
  wire  _T_1253; // @[MemPrimitives.scala 82:210:@9701.4]
  wire  _T_1256; // @[MemPrimitives.scala 83:102:@9703.4]
  wire [9:0] _T_1258; // @[Cat.scala 30:58:@9705.4]
  wire [9:0] _T_1260; // @[Cat.scala 30:58:@9707.4]
  wire [9:0] _T_1261; // @[Mux.scala 31:69:@9708.4]
  wire  _T_1266; // @[MemPrimitives.scala 82:210:@9715.4]
  wire  _T_1269; // @[MemPrimitives.scala 83:102:@9717.4]
  wire  _T_1271; // @[MemPrimitives.scala 82:210:@9718.4]
  wire  _T_1274; // @[MemPrimitives.scala 83:102:@9720.4]
  wire [9:0] _T_1276; // @[Cat.scala 30:58:@9722.4]
  wire [9:0] _T_1278; // @[Cat.scala 30:58:@9724.4]
  wire [9:0] _T_1279; // @[Mux.scala 31:69:@9725.4]
  wire  _T_1284; // @[MemPrimitives.scala 82:210:@9732.4]
  wire  _T_1287; // @[MemPrimitives.scala 83:102:@9734.4]
  wire  _T_1289; // @[MemPrimitives.scala 82:210:@9735.4]
  wire  _T_1292; // @[MemPrimitives.scala 83:102:@9737.4]
  wire [9:0] _T_1294; // @[Cat.scala 30:58:@9739.4]
  wire [9:0] _T_1296; // @[Cat.scala 30:58:@9741.4]
  wire [9:0] _T_1297; // @[Mux.scala 31:69:@9742.4]
  wire  _T_1302; // @[MemPrimitives.scala 82:210:@9749.4]
  wire  _T_1305; // @[MemPrimitives.scala 83:102:@9751.4]
  wire  _T_1307; // @[MemPrimitives.scala 82:210:@9752.4]
  wire  _T_1310; // @[MemPrimitives.scala 83:102:@9754.4]
  wire [9:0] _T_1312; // @[Cat.scala 30:58:@9756.4]
  wire [9:0] _T_1314; // @[Cat.scala 30:58:@9758.4]
  wire [9:0] _T_1315; // @[Mux.scala 31:69:@9759.4]
  wire  _T_1320; // @[MemPrimitives.scala 110:210:@9766.4]
  wire  _T_1325; // @[MemPrimitives.scala 110:210:@9769.4]
  wire  _T_1330; // @[MemPrimitives.scala 110:210:@9772.4]
  wire  _T_1335; // @[MemPrimitives.scala 110:210:@9775.4]
  wire  _T_1339; // @[MemPrimitives.scala 123:41:@9785.4]
  wire  _T_1340; // @[MemPrimitives.scala 123:41:@9786.4]
  wire  _T_1341; // @[MemPrimitives.scala 123:41:@9787.4]
  wire  _T_1342; // @[MemPrimitives.scala 123:41:@9788.4]
  wire [2:0] _T_1344; // @[Cat.scala 30:58:@9790.4]
  wire [2:0] _T_1346; // @[Cat.scala 30:58:@9792.4]
  wire [2:0] _T_1348; // @[Cat.scala 30:58:@9794.4]
  wire [2:0] _T_1350; // @[Cat.scala 30:58:@9796.4]
  wire [2:0] _T_1351; // @[Mux.scala 31:69:@9797.4]
  wire [2:0] _T_1352; // @[Mux.scala 31:69:@9798.4]
  wire [2:0] _T_1353; // @[Mux.scala 31:69:@9799.4]
  wire  _T_1358; // @[MemPrimitives.scala 110:210:@9806.4]
  wire  _T_1363; // @[MemPrimitives.scala 110:210:@9809.4]
  wire  _T_1368; // @[MemPrimitives.scala 110:210:@9812.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:210:@9815.4]
  wire  _T_1377; // @[MemPrimitives.scala 123:41:@9825.4]
  wire  _T_1378; // @[MemPrimitives.scala 123:41:@9826.4]
  wire  _T_1379; // @[MemPrimitives.scala 123:41:@9827.4]
  wire  _T_1380; // @[MemPrimitives.scala 123:41:@9828.4]
  wire [2:0] _T_1382; // @[Cat.scala 30:58:@9830.4]
  wire [2:0] _T_1384; // @[Cat.scala 30:58:@9832.4]
  wire [2:0] _T_1386; // @[Cat.scala 30:58:@9834.4]
  wire [2:0] _T_1388; // @[Cat.scala 30:58:@9836.4]
  wire [2:0] _T_1389; // @[Mux.scala 31:69:@9837.4]
  wire [2:0] _T_1390; // @[Mux.scala 31:69:@9838.4]
  wire [2:0] _T_1391; // @[Mux.scala 31:69:@9839.4]
  wire  _T_1396; // @[MemPrimitives.scala 110:210:@9846.4]
  wire  _T_1401; // @[MemPrimitives.scala 110:210:@9849.4]
  wire  _T_1406; // @[MemPrimitives.scala 110:210:@9852.4]
  wire  _T_1411; // @[MemPrimitives.scala 110:210:@9855.4]
  wire  _T_1416; // @[MemPrimitives.scala 110:210:@9858.4]
  wire  _T_1421; // @[MemPrimitives.scala 110:210:@9861.4]
  wire  _T_1426; // @[MemPrimitives.scala 110:210:@9864.4]
  wire  _T_1431; // @[MemPrimitives.scala 110:210:@9867.4]
  wire  _T_1435; // @[MemPrimitives.scala 123:41:@9881.4]
  wire  _T_1436; // @[MemPrimitives.scala 123:41:@9882.4]
  wire  _T_1437; // @[MemPrimitives.scala 123:41:@9883.4]
  wire  _T_1438; // @[MemPrimitives.scala 123:41:@9884.4]
  wire  _T_1439; // @[MemPrimitives.scala 123:41:@9885.4]
  wire  _T_1440; // @[MemPrimitives.scala 123:41:@9886.4]
  wire  _T_1441; // @[MemPrimitives.scala 123:41:@9887.4]
  wire  _T_1442; // @[MemPrimitives.scala 123:41:@9888.4]
  wire [2:0] _T_1444; // @[Cat.scala 30:58:@9890.4]
  wire [2:0] _T_1446; // @[Cat.scala 30:58:@9892.4]
  wire [2:0] _T_1448; // @[Cat.scala 30:58:@9894.4]
  wire [2:0] _T_1450; // @[Cat.scala 30:58:@9896.4]
  wire [2:0] _T_1452; // @[Cat.scala 30:58:@9898.4]
  wire [2:0] _T_1454; // @[Cat.scala 30:58:@9900.4]
  wire [2:0] _T_1456; // @[Cat.scala 30:58:@9902.4]
  wire [2:0] _T_1458; // @[Cat.scala 30:58:@9904.4]
  wire [2:0] _T_1459; // @[Mux.scala 31:69:@9905.4]
  wire [2:0] _T_1460; // @[Mux.scala 31:69:@9906.4]
  wire [2:0] _T_1461; // @[Mux.scala 31:69:@9907.4]
  wire [2:0] _T_1462; // @[Mux.scala 31:69:@9908.4]
  wire [2:0] _T_1463; // @[Mux.scala 31:69:@9909.4]
  wire [2:0] _T_1464; // @[Mux.scala 31:69:@9910.4]
  wire [2:0] _T_1465; // @[Mux.scala 31:69:@9911.4]
  wire  _T_1470; // @[MemPrimitives.scala 110:210:@9918.4]
  wire  _T_1475; // @[MemPrimitives.scala 110:210:@9921.4]
  wire  _T_1480; // @[MemPrimitives.scala 110:210:@9924.4]
  wire  _T_1485; // @[MemPrimitives.scala 110:210:@9927.4]
  wire  _T_1490; // @[MemPrimitives.scala 110:210:@9930.4]
  wire  _T_1495; // @[MemPrimitives.scala 110:210:@9933.4]
  wire  _T_1500; // @[MemPrimitives.scala 110:210:@9936.4]
  wire  _T_1505; // @[MemPrimitives.scala 110:210:@9939.4]
  wire  _T_1509; // @[MemPrimitives.scala 123:41:@9953.4]
  wire  _T_1510; // @[MemPrimitives.scala 123:41:@9954.4]
  wire  _T_1511; // @[MemPrimitives.scala 123:41:@9955.4]
  wire  _T_1512; // @[MemPrimitives.scala 123:41:@9956.4]
  wire  _T_1513; // @[MemPrimitives.scala 123:41:@9957.4]
  wire  _T_1514; // @[MemPrimitives.scala 123:41:@9958.4]
  wire  _T_1515; // @[MemPrimitives.scala 123:41:@9959.4]
  wire  _T_1516; // @[MemPrimitives.scala 123:41:@9960.4]
  wire [2:0] _T_1518; // @[Cat.scala 30:58:@9962.4]
  wire [2:0] _T_1520; // @[Cat.scala 30:58:@9964.4]
  wire [2:0] _T_1522; // @[Cat.scala 30:58:@9966.4]
  wire [2:0] _T_1524; // @[Cat.scala 30:58:@9968.4]
  wire [2:0] _T_1526; // @[Cat.scala 30:58:@9970.4]
  wire [2:0] _T_1528; // @[Cat.scala 30:58:@9972.4]
  wire [2:0] _T_1530; // @[Cat.scala 30:58:@9974.4]
  wire [2:0] _T_1532; // @[Cat.scala 30:58:@9976.4]
  wire [2:0] _T_1533; // @[Mux.scala 31:69:@9977.4]
  wire [2:0] _T_1534; // @[Mux.scala 31:69:@9978.4]
  wire [2:0] _T_1535; // @[Mux.scala 31:69:@9979.4]
  wire [2:0] _T_1536; // @[Mux.scala 31:69:@9980.4]
  wire [2:0] _T_1537; // @[Mux.scala 31:69:@9981.4]
  wire [2:0] _T_1538; // @[Mux.scala 31:69:@9982.4]
  wire [2:0] _T_1539; // @[Mux.scala 31:69:@9983.4]
  wire  _T_1544; // @[MemPrimitives.scala 110:210:@9990.4]
  wire  _T_1549; // @[MemPrimitives.scala 110:210:@9993.4]
  wire  _T_1554; // @[MemPrimitives.scala 110:210:@9996.4]
  wire  _T_1559; // @[MemPrimitives.scala 110:210:@9999.4]
  wire  _T_1563; // @[MemPrimitives.scala 123:41:@10009.4]
  wire  _T_1564; // @[MemPrimitives.scala 123:41:@10010.4]
  wire  _T_1565; // @[MemPrimitives.scala 123:41:@10011.4]
  wire  _T_1566; // @[MemPrimitives.scala 123:41:@10012.4]
  wire [2:0] _T_1568; // @[Cat.scala 30:58:@10014.4]
  wire [2:0] _T_1570; // @[Cat.scala 30:58:@10016.4]
  wire [2:0] _T_1572; // @[Cat.scala 30:58:@10018.4]
  wire [2:0] _T_1574; // @[Cat.scala 30:58:@10020.4]
  wire [2:0] _T_1575; // @[Mux.scala 31:69:@10021.4]
  wire [2:0] _T_1576; // @[Mux.scala 31:69:@10022.4]
  wire [2:0] _T_1577; // @[Mux.scala 31:69:@10023.4]
  wire  _T_1582; // @[MemPrimitives.scala 110:210:@10030.4]
  wire  _T_1587; // @[MemPrimitives.scala 110:210:@10033.4]
  wire  _T_1592; // @[MemPrimitives.scala 110:210:@10036.4]
  wire  _T_1597; // @[MemPrimitives.scala 110:210:@10039.4]
  wire  _T_1601; // @[MemPrimitives.scala 123:41:@10049.4]
  wire  _T_1602; // @[MemPrimitives.scala 123:41:@10050.4]
  wire  _T_1603; // @[MemPrimitives.scala 123:41:@10051.4]
  wire  _T_1604; // @[MemPrimitives.scala 123:41:@10052.4]
  wire [2:0] _T_1606; // @[Cat.scala 30:58:@10054.4]
  wire [2:0] _T_1608; // @[Cat.scala 30:58:@10056.4]
  wire [2:0] _T_1610; // @[Cat.scala 30:58:@10058.4]
  wire [2:0] _T_1612; // @[Cat.scala 30:58:@10060.4]
  wire [2:0] _T_1613; // @[Mux.scala 31:69:@10061.4]
  wire [2:0] _T_1614; // @[Mux.scala 31:69:@10062.4]
  wire [2:0] _T_1615; // @[Mux.scala 31:69:@10063.4]
  wire  _T_1620; // @[MemPrimitives.scala 110:210:@10070.4]
  wire  _T_1625; // @[MemPrimitives.scala 110:210:@10073.4]
  wire  _T_1630; // @[MemPrimitives.scala 110:210:@10076.4]
  wire  _T_1635; // @[MemPrimitives.scala 110:210:@10079.4]
  wire  _T_1640; // @[MemPrimitives.scala 110:210:@10082.4]
  wire  _T_1645; // @[MemPrimitives.scala 110:210:@10085.4]
  wire  _T_1650; // @[MemPrimitives.scala 110:210:@10088.4]
  wire  _T_1655; // @[MemPrimitives.scala 110:210:@10091.4]
  wire  _T_1659; // @[MemPrimitives.scala 123:41:@10105.4]
  wire  _T_1660; // @[MemPrimitives.scala 123:41:@10106.4]
  wire  _T_1661; // @[MemPrimitives.scala 123:41:@10107.4]
  wire  _T_1662; // @[MemPrimitives.scala 123:41:@10108.4]
  wire  _T_1663; // @[MemPrimitives.scala 123:41:@10109.4]
  wire  _T_1664; // @[MemPrimitives.scala 123:41:@10110.4]
  wire  _T_1665; // @[MemPrimitives.scala 123:41:@10111.4]
  wire  _T_1666; // @[MemPrimitives.scala 123:41:@10112.4]
  wire [2:0] _T_1668; // @[Cat.scala 30:58:@10114.4]
  wire [2:0] _T_1670; // @[Cat.scala 30:58:@10116.4]
  wire [2:0] _T_1672; // @[Cat.scala 30:58:@10118.4]
  wire [2:0] _T_1674; // @[Cat.scala 30:58:@10120.4]
  wire [2:0] _T_1676; // @[Cat.scala 30:58:@10122.4]
  wire [2:0] _T_1678; // @[Cat.scala 30:58:@10124.4]
  wire [2:0] _T_1680; // @[Cat.scala 30:58:@10126.4]
  wire [2:0] _T_1682; // @[Cat.scala 30:58:@10128.4]
  wire [2:0] _T_1683; // @[Mux.scala 31:69:@10129.4]
  wire [2:0] _T_1684; // @[Mux.scala 31:69:@10130.4]
  wire [2:0] _T_1685; // @[Mux.scala 31:69:@10131.4]
  wire [2:0] _T_1686; // @[Mux.scala 31:69:@10132.4]
  wire [2:0] _T_1687; // @[Mux.scala 31:69:@10133.4]
  wire [2:0] _T_1688; // @[Mux.scala 31:69:@10134.4]
  wire [2:0] _T_1689; // @[Mux.scala 31:69:@10135.4]
  wire  _T_1694; // @[MemPrimitives.scala 110:210:@10142.4]
  wire  _T_1699; // @[MemPrimitives.scala 110:210:@10145.4]
  wire  _T_1704; // @[MemPrimitives.scala 110:210:@10148.4]
  wire  _T_1709; // @[MemPrimitives.scala 110:210:@10151.4]
  wire  _T_1714; // @[MemPrimitives.scala 110:210:@10154.4]
  wire  _T_1719; // @[MemPrimitives.scala 110:210:@10157.4]
  wire  _T_1724; // @[MemPrimitives.scala 110:210:@10160.4]
  wire  _T_1729; // @[MemPrimitives.scala 110:210:@10163.4]
  wire  _T_1733; // @[MemPrimitives.scala 123:41:@10177.4]
  wire  _T_1734; // @[MemPrimitives.scala 123:41:@10178.4]
  wire  _T_1735; // @[MemPrimitives.scala 123:41:@10179.4]
  wire  _T_1736; // @[MemPrimitives.scala 123:41:@10180.4]
  wire  _T_1737; // @[MemPrimitives.scala 123:41:@10181.4]
  wire  _T_1738; // @[MemPrimitives.scala 123:41:@10182.4]
  wire  _T_1739; // @[MemPrimitives.scala 123:41:@10183.4]
  wire  _T_1740; // @[MemPrimitives.scala 123:41:@10184.4]
  wire [2:0] _T_1742; // @[Cat.scala 30:58:@10186.4]
  wire [2:0] _T_1744; // @[Cat.scala 30:58:@10188.4]
  wire [2:0] _T_1746; // @[Cat.scala 30:58:@10190.4]
  wire [2:0] _T_1748; // @[Cat.scala 30:58:@10192.4]
  wire [2:0] _T_1750; // @[Cat.scala 30:58:@10194.4]
  wire [2:0] _T_1752; // @[Cat.scala 30:58:@10196.4]
  wire [2:0] _T_1754; // @[Cat.scala 30:58:@10198.4]
  wire [2:0] _T_1756; // @[Cat.scala 30:58:@10200.4]
  wire [2:0] _T_1757; // @[Mux.scala 31:69:@10201.4]
  wire [2:0] _T_1758; // @[Mux.scala 31:69:@10202.4]
  wire [2:0] _T_1759; // @[Mux.scala 31:69:@10203.4]
  wire [2:0] _T_1760; // @[Mux.scala 31:69:@10204.4]
  wire [2:0] _T_1761; // @[Mux.scala 31:69:@10205.4]
  wire [2:0] _T_1762; // @[Mux.scala 31:69:@10206.4]
  wire [2:0] _T_1763; // @[Mux.scala 31:69:@10207.4]
  wire  _T_1768; // @[MemPrimitives.scala 110:210:@10214.4]
  wire  _T_1773; // @[MemPrimitives.scala 110:210:@10217.4]
  wire  _T_1778; // @[MemPrimitives.scala 110:210:@10220.4]
  wire  _T_1783; // @[MemPrimitives.scala 110:210:@10223.4]
  wire  _T_1787; // @[MemPrimitives.scala 123:41:@10233.4]
  wire  _T_1788; // @[MemPrimitives.scala 123:41:@10234.4]
  wire  _T_1789; // @[MemPrimitives.scala 123:41:@10235.4]
  wire  _T_1790; // @[MemPrimitives.scala 123:41:@10236.4]
  wire [2:0] _T_1792; // @[Cat.scala 30:58:@10238.4]
  wire [2:0] _T_1794; // @[Cat.scala 30:58:@10240.4]
  wire [2:0] _T_1796; // @[Cat.scala 30:58:@10242.4]
  wire [2:0] _T_1798; // @[Cat.scala 30:58:@10244.4]
  wire [2:0] _T_1799; // @[Mux.scala 31:69:@10245.4]
  wire [2:0] _T_1800; // @[Mux.scala 31:69:@10246.4]
  wire [2:0] _T_1801; // @[Mux.scala 31:69:@10247.4]
  wire  _T_1806; // @[MemPrimitives.scala 110:210:@10254.4]
  wire  _T_1811; // @[MemPrimitives.scala 110:210:@10257.4]
  wire  _T_1816; // @[MemPrimitives.scala 110:210:@10260.4]
  wire  _T_1821; // @[MemPrimitives.scala 110:210:@10263.4]
  wire  _T_1825; // @[MemPrimitives.scala 123:41:@10273.4]
  wire  _T_1826; // @[MemPrimitives.scala 123:41:@10274.4]
  wire  _T_1827; // @[MemPrimitives.scala 123:41:@10275.4]
  wire  _T_1828; // @[MemPrimitives.scala 123:41:@10276.4]
  wire [2:0] _T_1830; // @[Cat.scala 30:58:@10278.4]
  wire [2:0] _T_1832; // @[Cat.scala 30:58:@10280.4]
  wire [2:0] _T_1834; // @[Cat.scala 30:58:@10282.4]
  wire [2:0] _T_1836; // @[Cat.scala 30:58:@10284.4]
  wire [2:0] _T_1837; // @[Mux.scala 31:69:@10285.4]
  wire [2:0] _T_1838; // @[Mux.scala 31:69:@10286.4]
  wire [2:0] _T_1839; // @[Mux.scala 31:69:@10287.4]
  wire  _T_1844; // @[MemPrimitives.scala 110:210:@10294.4]
  wire  _T_1849; // @[MemPrimitives.scala 110:210:@10297.4]
  wire  _T_1854; // @[MemPrimitives.scala 110:210:@10300.4]
  wire  _T_1859; // @[MemPrimitives.scala 110:210:@10303.4]
  wire  _T_1864; // @[MemPrimitives.scala 110:210:@10306.4]
  wire  _T_1869; // @[MemPrimitives.scala 110:210:@10309.4]
  wire  _T_1874; // @[MemPrimitives.scala 110:210:@10312.4]
  wire  _T_1879; // @[MemPrimitives.scala 110:210:@10315.4]
  wire  _T_1883; // @[MemPrimitives.scala 123:41:@10329.4]
  wire  _T_1884; // @[MemPrimitives.scala 123:41:@10330.4]
  wire  _T_1885; // @[MemPrimitives.scala 123:41:@10331.4]
  wire  _T_1886; // @[MemPrimitives.scala 123:41:@10332.4]
  wire  _T_1887; // @[MemPrimitives.scala 123:41:@10333.4]
  wire  _T_1888; // @[MemPrimitives.scala 123:41:@10334.4]
  wire  _T_1889; // @[MemPrimitives.scala 123:41:@10335.4]
  wire  _T_1890; // @[MemPrimitives.scala 123:41:@10336.4]
  wire [2:0] _T_1892; // @[Cat.scala 30:58:@10338.4]
  wire [2:0] _T_1894; // @[Cat.scala 30:58:@10340.4]
  wire [2:0] _T_1896; // @[Cat.scala 30:58:@10342.4]
  wire [2:0] _T_1898; // @[Cat.scala 30:58:@10344.4]
  wire [2:0] _T_1900; // @[Cat.scala 30:58:@10346.4]
  wire [2:0] _T_1902; // @[Cat.scala 30:58:@10348.4]
  wire [2:0] _T_1904; // @[Cat.scala 30:58:@10350.4]
  wire [2:0] _T_1906; // @[Cat.scala 30:58:@10352.4]
  wire [2:0] _T_1907; // @[Mux.scala 31:69:@10353.4]
  wire [2:0] _T_1908; // @[Mux.scala 31:69:@10354.4]
  wire [2:0] _T_1909; // @[Mux.scala 31:69:@10355.4]
  wire [2:0] _T_1910; // @[Mux.scala 31:69:@10356.4]
  wire [2:0] _T_1911; // @[Mux.scala 31:69:@10357.4]
  wire [2:0] _T_1912; // @[Mux.scala 31:69:@10358.4]
  wire [2:0] _T_1913; // @[Mux.scala 31:69:@10359.4]
  wire  _T_1918; // @[MemPrimitives.scala 110:210:@10366.4]
  wire  _T_1923; // @[MemPrimitives.scala 110:210:@10369.4]
  wire  _T_1928; // @[MemPrimitives.scala 110:210:@10372.4]
  wire  _T_1933; // @[MemPrimitives.scala 110:210:@10375.4]
  wire  _T_1938; // @[MemPrimitives.scala 110:210:@10378.4]
  wire  _T_1943; // @[MemPrimitives.scala 110:210:@10381.4]
  wire  _T_1948; // @[MemPrimitives.scala 110:210:@10384.4]
  wire  _T_1953; // @[MemPrimitives.scala 110:210:@10387.4]
  wire  _T_1957; // @[MemPrimitives.scala 123:41:@10401.4]
  wire  _T_1958; // @[MemPrimitives.scala 123:41:@10402.4]
  wire  _T_1959; // @[MemPrimitives.scala 123:41:@10403.4]
  wire  _T_1960; // @[MemPrimitives.scala 123:41:@10404.4]
  wire  _T_1961; // @[MemPrimitives.scala 123:41:@10405.4]
  wire  _T_1962; // @[MemPrimitives.scala 123:41:@10406.4]
  wire  _T_1963; // @[MemPrimitives.scala 123:41:@10407.4]
  wire  _T_1964; // @[MemPrimitives.scala 123:41:@10408.4]
  wire [2:0] _T_1966; // @[Cat.scala 30:58:@10410.4]
  wire [2:0] _T_1968; // @[Cat.scala 30:58:@10412.4]
  wire [2:0] _T_1970; // @[Cat.scala 30:58:@10414.4]
  wire [2:0] _T_1972; // @[Cat.scala 30:58:@10416.4]
  wire [2:0] _T_1974; // @[Cat.scala 30:58:@10418.4]
  wire [2:0] _T_1976; // @[Cat.scala 30:58:@10420.4]
  wire [2:0] _T_1978; // @[Cat.scala 30:58:@10422.4]
  wire [2:0] _T_1980; // @[Cat.scala 30:58:@10424.4]
  wire [2:0] _T_1981; // @[Mux.scala 31:69:@10425.4]
  wire [2:0] _T_1982; // @[Mux.scala 31:69:@10426.4]
  wire [2:0] _T_1983; // @[Mux.scala 31:69:@10427.4]
  wire [2:0] _T_1984; // @[Mux.scala 31:69:@10428.4]
  wire [2:0] _T_1985; // @[Mux.scala 31:69:@10429.4]
  wire [2:0] _T_1986; // @[Mux.scala 31:69:@10430.4]
  wire [2:0] _T_1987; // @[Mux.scala 31:69:@10431.4]
  wire  _T_1992; // @[MemPrimitives.scala 110:210:@10438.4]
  wire  _T_1997; // @[MemPrimitives.scala 110:210:@10441.4]
  wire  _T_2002; // @[MemPrimitives.scala 110:210:@10444.4]
  wire  _T_2007; // @[MemPrimitives.scala 110:210:@10447.4]
  wire  _T_2011; // @[MemPrimitives.scala 123:41:@10457.4]
  wire  _T_2012; // @[MemPrimitives.scala 123:41:@10458.4]
  wire  _T_2013; // @[MemPrimitives.scala 123:41:@10459.4]
  wire  _T_2014; // @[MemPrimitives.scala 123:41:@10460.4]
  wire [2:0] _T_2016; // @[Cat.scala 30:58:@10462.4]
  wire [2:0] _T_2018; // @[Cat.scala 30:58:@10464.4]
  wire [2:0] _T_2020; // @[Cat.scala 30:58:@10466.4]
  wire [2:0] _T_2022; // @[Cat.scala 30:58:@10468.4]
  wire [2:0] _T_2023; // @[Mux.scala 31:69:@10469.4]
  wire [2:0] _T_2024; // @[Mux.scala 31:69:@10470.4]
  wire [2:0] _T_2025; // @[Mux.scala 31:69:@10471.4]
  wire  _T_2030; // @[MemPrimitives.scala 110:210:@10478.4]
  wire  _T_2035; // @[MemPrimitives.scala 110:210:@10481.4]
  wire  _T_2040; // @[MemPrimitives.scala 110:210:@10484.4]
  wire  _T_2045; // @[MemPrimitives.scala 110:210:@10487.4]
  wire  _T_2049; // @[MemPrimitives.scala 123:41:@10497.4]
  wire  _T_2050; // @[MemPrimitives.scala 123:41:@10498.4]
  wire  _T_2051; // @[MemPrimitives.scala 123:41:@10499.4]
  wire  _T_2052; // @[MemPrimitives.scala 123:41:@10500.4]
  wire [2:0] _T_2054; // @[Cat.scala 30:58:@10502.4]
  wire [2:0] _T_2056; // @[Cat.scala 30:58:@10504.4]
  wire [2:0] _T_2058; // @[Cat.scala 30:58:@10506.4]
  wire [2:0] _T_2060; // @[Cat.scala 30:58:@10508.4]
  wire [2:0] _T_2061; // @[Mux.scala 31:69:@10509.4]
  wire [2:0] _T_2062; // @[Mux.scala 31:69:@10510.4]
  wire [2:0] _T_2063; // @[Mux.scala 31:69:@10511.4]
  wire  _T_2068; // @[MemPrimitives.scala 110:210:@10518.4]
  wire  _T_2073; // @[MemPrimitives.scala 110:210:@10521.4]
  wire  _T_2078; // @[MemPrimitives.scala 110:210:@10524.4]
  wire  _T_2083; // @[MemPrimitives.scala 110:210:@10527.4]
  wire  _T_2088; // @[MemPrimitives.scala 110:210:@10530.4]
  wire  _T_2093; // @[MemPrimitives.scala 110:210:@10533.4]
  wire  _T_2098; // @[MemPrimitives.scala 110:210:@10536.4]
  wire  _T_2103; // @[MemPrimitives.scala 110:210:@10539.4]
  wire  _T_2107; // @[MemPrimitives.scala 123:41:@10553.4]
  wire  _T_2108; // @[MemPrimitives.scala 123:41:@10554.4]
  wire  _T_2109; // @[MemPrimitives.scala 123:41:@10555.4]
  wire  _T_2110; // @[MemPrimitives.scala 123:41:@10556.4]
  wire  _T_2111; // @[MemPrimitives.scala 123:41:@10557.4]
  wire  _T_2112; // @[MemPrimitives.scala 123:41:@10558.4]
  wire  _T_2113; // @[MemPrimitives.scala 123:41:@10559.4]
  wire  _T_2114; // @[MemPrimitives.scala 123:41:@10560.4]
  wire [2:0] _T_2116; // @[Cat.scala 30:58:@10562.4]
  wire [2:0] _T_2118; // @[Cat.scala 30:58:@10564.4]
  wire [2:0] _T_2120; // @[Cat.scala 30:58:@10566.4]
  wire [2:0] _T_2122; // @[Cat.scala 30:58:@10568.4]
  wire [2:0] _T_2124; // @[Cat.scala 30:58:@10570.4]
  wire [2:0] _T_2126; // @[Cat.scala 30:58:@10572.4]
  wire [2:0] _T_2128; // @[Cat.scala 30:58:@10574.4]
  wire [2:0] _T_2130; // @[Cat.scala 30:58:@10576.4]
  wire [2:0] _T_2131; // @[Mux.scala 31:69:@10577.4]
  wire [2:0] _T_2132; // @[Mux.scala 31:69:@10578.4]
  wire [2:0] _T_2133; // @[Mux.scala 31:69:@10579.4]
  wire [2:0] _T_2134; // @[Mux.scala 31:69:@10580.4]
  wire [2:0] _T_2135; // @[Mux.scala 31:69:@10581.4]
  wire [2:0] _T_2136; // @[Mux.scala 31:69:@10582.4]
  wire [2:0] _T_2137; // @[Mux.scala 31:69:@10583.4]
  wire  _T_2142; // @[MemPrimitives.scala 110:210:@10590.4]
  wire  _T_2147; // @[MemPrimitives.scala 110:210:@10593.4]
  wire  _T_2152; // @[MemPrimitives.scala 110:210:@10596.4]
  wire  _T_2157; // @[MemPrimitives.scala 110:210:@10599.4]
  wire  _T_2162; // @[MemPrimitives.scala 110:210:@10602.4]
  wire  _T_2167; // @[MemPrimitives.scala 110:210:@10605.4]
  wire  _T_2172; // @[MemPrimitives.scala 110:210:@10608.4]
  wire  _T_2177; // @[MemPrimitives.scala 110:210:@10611.4]
  wire  _T_2181; // @[MemPrimitives.scala 123:41:@10625.4]
  wire  _T_2182; // @[MemPrimitives.scala 123:41:@10626.4]
  wire  _T_2183; // @[MemPrimitives.scala 123:41:@10627.4]
  wire  _T_2184; // @[MemPrimitives.scala 123:41:@10628.4]
  wire  _T_2185; // @[MemPrimitives.scala 123:41:@10629.4]
  wire  _T_2186; // @[MemPrimitives.scala 123:41:@10630.4]
  wire  _T_2187; // @[MemPrimitives.scala 123:41:@10631.4]
  wire  _T_2188; // @[MemPrimitives.scala 123:41:@10632.4]
  wire [2:0] _T_2190; // @[Cat.scala 30:58:@10634.4]
  wire [2:0] _T_2192; // @[Cat.scala 30:58:@10636.4]
  wire [2:0] _T_2194; // @[Cat.scala 30:58:@10638.4]
  wire [2:0] _T_2196; // @[Cat.scala 30:58:@10640.4]
  wire [2:0] _T_2198; // @[Cat.scala 30:58:@10642.4]
  wire [2:0] _T_2200; // @[Cat.scala 30:58:@10644.4]
  wire [2:0] _T_2202; // @[Cat.scala 30:58:@10646.4]
  wire [2:0] _T_2204; // @[Cat.scala 30:58:@10648.4]
  wire [2:0] _T_2205; // @[Mux.scala 31:69:@10649.4]
  wire [2:0] _T_2206; // @[Mux.scala 31:69:@10650.4]
  wire [2:0] _T_2207; // @[Mux.scala 31:69:@10651.4]
  wire [2:0] _T_2208; // @[Mux.scala 31:69:@10652.4]
  wire [2:0] _T_2209; // @[Mux.scala 31:69:@10653.4]
  wire [2:0] _T_2210; // @[Mux.scala 31:69:@10654.4]
  wire [2:0] _T_2211; // @[Mux.scala 31:69:@10655.4]
  wire  _T_2243; // @[package.scala 96:25:@10696.4 package.scala 96:25:@10697.4]
  wire [7:0] _T_2247; // @[Mux.scala 31:69:@10706.4]
  wire  _T_2240; // @[package.scala 96:25:@10688.4 package.scala 96:25:@10689.4]
  wire [7:0] _T_2248; // @[Mux.scala 31:69:@10707.4]
  wire  _T_2237; // @[package.scala 96:25:@10680.4 package.scala 96:25:@10681.4]
  wire  _T_2278; // @[package.scala 96:25:@10744.4 package.scala 96:25:@10745.4]
  wire [7:0] _T_2282; // @[Mux.scala 31:69:@10754.4]
  wire  _T_2275; // @[package.scala 96:25:@10736.4 package.scala 96:25:@10737.4]
  wire [7:0] _T_2283; // @[Mux.scala 31:69:@10755.4]
  wire  _T_2272; // @[package.scala 96:25:@10728.4 package.scala 96:25:@10729.4]
  wire  _T_2313; // @[package.scala 96:25:@10792.4 package.scala 96:25:@10793.4]
  wire [7:0] _T_2317; // @[Mux.scala 31:69:@10802.4]
  wire  _T_2310; // @[package.scala 96:25:@10784.4 package.scala 96:25:@10785.4]
  wire [7:0] _T_2318; // @[Mux.scala 31:69:@10803.4]
  wire  _T_2307; // @[package.scala 96:25:@10776.4 package.scala 96:25:@10777.4]
  wire  _T_2348; // @[package.scala 96:25:@10840.4 package.scala 96:25:@10841.4]
  wire [7:0] _T_2352; // @[Mux.scala 31:69:@10850.4]
  wire  _T_2345; // @[package.scala 96:25:@10832.4 package.scala 96:25:@10833.4]
  wire [7:0] _T_2353; // @[Mux.scala 31:69:@10851.4]
  wire  _T_2342; // @[package.scala 96:25:@10824.4 package.scala 96:25:@10825.4]
  wire  _T_2383; // @[package.scala 96:25:@10888.4 package.scala 96:25:@10889.4]
  wire [7:0] _T_2387; // @[Mux.scala 31:69:@10898.4]
  wire  _T_2380; // @[package.scala 96:25:@10880.4 package.scala 96:25:@10881.4]
  wire [7:0] _T_2388; // @[Mux.scala 31:69:@10899.4]
  wire  _T_2377; // @[package.scala 96:25:@10872.4 package.scala 96:25:@10873.4]
  wire  _T_2418; // @[package.scala 96:25:@10936.4 package.scala 96:25:@10937.4]
  wire [7:0] _T_2422; // @[Mux.scala 31:69:@10946.4]
  wire  _T_2415; // @[package.scala 96:25:@10928.4 package.scala 96:25:@10929.4]
  wire [7:0] _T_2423; // @[Mux.scala 31:69:@10947.4]
  wire  _T_2412; // @[package.scala 96:25:@10920.4 package.scala 96:25:@10921.4]
  wire  _T_2453; // @[package.scala 96:25:@10984.4 package.scala 96:25:@10985.4]
  wire [7:0] _T_2457; // @[Mux.scala 31:69:@10994.4]
  wire  _T_2450; // @[package.scala 96:25:@10976.4 package.scala 96:25:@10977.4]
  wire [7:0] _T_2458; // @[Mux.scala 31:69:@10995.4]
  wire  _T_2447; // @[package.scala 96:25:@10968.4 package.scala 96:25:@10969.4]
  wire  _T_2488; // @[package.scala 96:25:@11032.4 package.scala 96:25:@11033.4]
  wire [7:0] _T_2492; // @[Mux.scala 31:69:@11042.4]
  wire  _T_2485; // @[package.scala 96:25:@11024.4 package.scala 96:25:@11025.4]
  wire [7:0] _T_2493; // @[Mux.scala 31:69:@11043.4]
  wire  _T_2482; // @[package.scala 96:25:@11016.4 package.scala 96:25:@11017.4]
  wire  _T_2523; // @[package.scala 96:25:@11080.4 package.scala 96:25:@11081.4]
  wire [7:0] _T_2527; // @[Mux.scala 31:69:@11090.4]
  wire  _T_2520; // @[package.scala 96:25:@11072.4 package.scala 96:25:@11073.4]
  wire [7:0] _T_2528; // @[Mux.scala 31:69:@11091.4]
  wire  _T_2517; // @[package.scala 96:25:@11064.4 package.scala 96:25:@11065.4]
  wire  _T_2558; // @[package.scala 96:25:@11128.4 package.scala 96:25:@11129.4]
  wire [7:0] _T_2562; // @[Mux.scala 31:69:@11138.4]
  wire  _T_2555; // @[package.scala 96:25:@11120.4 package.scala 96:25:@11121.4]
  wire [7:0] _T_2563; // @[Mux.scala 31:69:@11139.4]
  wire  _T_2552; // @[package.scala 96:25:@11112.4 package.scala 96:25:@11113.4]
  wire  _T_2593; // @[package.scala 96:25:@11176.4 package.scala 96:25:@11177.4]
  wire [7:0] _T_2597; // @[Mux.scala 31:69:@11186.4]
  wire  _T_2590; // @[package.scala 96:25:@11168.4 package.scala 96:25:@11169.4]
  wire [7:0] _T_2598; // @[Mux.scala 31:69:@11187.4]
  wire  _T_2587; // @[package.scala 96:25:@11160.4 package.scala 96:25:@11161.4]
  wire  _T_2628; // @[package.scala 96:25:@11224.4 package.scala 96:25:@11225.4]
  wire [7:0] _T_2632; // @[Mux.scala 31:69:@11234.4]
  wire  _T_2625; // @[package.scala 96:25:@11216.4 package.scala 96:25:@11217.4]
  wire [7:0] _T_2633; // @[Mux.scala 31:69:@11235.4]
  wire  _T_2622; // @[package.scala 96:25:@11208.4 package.scala 96:25:@11209.4]
  wire  _T_2663; // @[package.scala 96:25:@11272.4 package.scala 96:25:@11273.4]
  wire [7:0] _T_2667; // @[Mux.scala 31:69:@11282.4]
  wire  _T_2660; // @[package.scala 96:25:@11264.4 package.scala 96:25:@11265.4]
  wire [7:0] _T_2668; // @[Mux.scala 31:69:@11283.4]
  wire  _T_2657; // @[package.scala 96:25:@11256.4 package.scala 96:25:@11257.4]
  wire  _T_2698; // @[package.scala 96:25:@11320.4 package.scala 96:25:@11321.4]
  wire [7:0] _T_2702; // @[Mux.scala 31:69:@11330.4]
  wire  _T_2695; // @[package.scala 96:25:@11312.4 package.scala 96:25:@11313.4]
  wire [7:0] _T_2703; // @[Mux.scala 31:69:@11331.4]
  wire  _T_2692; // @[package.scala 96:25:@11304.4 package.scala 96:25:@11305.4]
  wire  _T_2733; // @[package.scala 96:25:@11368.4 package.scala 96:25:@11369.4]
  wire [7:0] _T_2737; // @[Mux.scala 31:69:@11378.4]
  wire  _T_2730; // @[package.scala 96:25:@11360.4 package.scala 96:25:@11361.4]
  wire [7:0] _T_2738; // @[Mux.scala 31:69:@11379.4]
  wire  _T_2727; // @[package.scala 96:25:@11352.4 package.scala 96:25:@11353.4]
  wire  _T_2768; // @[package.scala 96:25:@11416.4 package.scala 96:25:@11417.4]
  wire [7:0] _T_2772; // @[Mux.scala 31:69:@11426.4]
  wire  _T_2765; // @[package.scala 96:25:@11408.4 package.scala 96:25:@11409.4]
  wire [7:0] _T_2773; // @[Mux.scala 31:69:@11427.4]
  wire  _T_2762; // @[package.scala 96:25:@11400.4 package.scala 96:25:@11401.4]
  wire  _T_2803; // @[package.scala 96:25:@11464.4 package.scala 96:25:@11465.4]
  wire [7:0] _T_2807; // @[Mux.scala 31:69:@11474.4]
  wire  _T_2800; // @[package.scala 96:25:@11456.4 package.scala 96:25:@11457.4]
  wire [7:0] _T_2808; // @[Mux.scala 31:69:@11475.4]
  wire  _T_2797; // @[package.scala 96:25:@11448.4 package.scala 96:25:@11449.4]
  wire  _T_2838; // @[package.scala 96:25:@11512.4 package.scala 96:25:@11513.4]
  wire [7:0] _T_2842; // @[Mux.scala 31:69:@11522.4]
  wire  _T_2835; // @[package.scala 96:25:@11504.4 package.scala 96:25:@11505.4]
  wire [7:0] _T_2843; // @[Mux.scala 31:69:@11523.4]
  wire  _T_2832; // @[package.scala 96:25:@11496.4 package.scala 96:25:@11497.4]
  wire  _T_2873; // @[package.scala 96:25:@11560.4 package.scala 96:25:@11561.4]
  wire [7:0] _T_2877; // @[Mux.scala 31:69:@11570.4]
  wire  _T_2870; // @[package.scala 96:25:@11552.4 package.scala 96:25:@11553.4]
  wire [7:0] _T_2878; // @[Mux.scala 31:69:@11571.4]
  wire  _T_2867; // @[package.scala 96:25:@11544.4 package.scala 96:25:@11545.4]
  wire  _T_2908; // @[package.scala 96:25:@11608.4 package.scala 96:25:@11609.4]
  wire [7:0] _T_2912; // @[Mux.scala 31:69:@11618.4]
  wire  _T_2905; // @[package.scala 96:25:@11600.4 package.scala 96:25:@11601.4]
  wire [7:0] _T_2913; // @[Mux.scala 31:69:@11619.4]
  wire  _T_2902; // @[package.scala 96:25:@11592.4 package.scala 96:25:@11593.4]
  wire  _T_2943; // @[package.scala 96:25:@11656.4 package.scala 96:25:@11657.4]
  wire [7:0] _T_2947; // @[Mux.scala 31:69:@11666.4]
  wire  _T_2940; // @[package.scala 96:25:@11648.4 package.scala 96:25:@11649.4]
  wire [7:0] _T_2948; // @[Mux.scala 31:69:@11667.4]
  wire  _T_2937; // @[package.scala 96:25:@11640.4 package.scala 96:25:@11641.4]
  wire  _T_2978; // @[package.scala 96:25:@11704.4 package.scala 96:25:@11705.4]
  wire [7:0] _T_2982; // @[Mux.scala 31:69:@11714.4]
  wire  _T_2975; // @[package.scala 96:25:@11696.4 package.scala 96:25:@11697.4]
  wire [7:0] _T_2983; // @[Mux.scala 31:69:@11715.4]
  wire  _T_2972; // @[package.scala 96:25:@11688.4 package.scala 96:25:@11689.4]
  wire  _T_3013; // @[package.scala 96:25:@11752.4 package.scala 96:25:@11753.4]
  wire [7:0] _T_3017; // @[Mux.scala 31:69:@11762.4]
  wire  _T_3010; // @[package.scala 96:25:@11744.4 package.scala 96:25:@11745.4]
  wire [7:0] _T_3018; // @[Mux.scala 31:69:@11763.4]
  wire  _T_3007; // @[package.scala 96:25:@11736.4 package.scala 96:25:@11737.4]
  wire  _T_3048; // @[package.scala 96:25:@11800.4 package.scala 96:25:@11801.4]
  wire [7:0] _T_3052; // @[Mux.scala 31:69:@11810.4]
  wire  _T_3045; // @[package.scala 96:25:@11792.4 package.scala 96:25:@11793.4]
  wire [7:0] _T_3053; // @[Mux.scala 31:69:@11811.4]
  wire  _T_3042; // @[package.scala 96:25:@11784.4 package.scala 96:25:@11785.4]
  Mem1D_4 Mem1D ( // @[MemPrimitives.scala 64:21:@9238.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_4 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@9254.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_4 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@9270.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_4 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@9286.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_4 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@9302.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_4 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@9318.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_4 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@9334.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_4 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@9350.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_4 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@9366.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_4 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@9382.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_4 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@9398.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_4 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@9414.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_4 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@9430.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_4 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@9446.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_4 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@9462.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_4 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@9478.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@9778.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3)
  );
  StickySelects StickySelects_1 ( // @[MemPrimitives.scala 121:29:@9818.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3)
  );
  StickySelects_2 StickySelects_2 ( // @[MemPrimitives.scala 121:29:@9870.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7)
  );
  StickySelects_2 StickySelects_3 ( // @[MemPrimitives.scala 121:29:@9942.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7)
  );
  StickySelects StickySelects_4 ( // @[MemPrimitives.scala 121:29:@10002.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3)
  );
  StickySelects StickySelects_5 ( // @[MemPrimitives.scala 121:29:@10042.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3)
  );
  StickySelects_2 StickySelects_6 ( // @[MemPrimitives.scala 121:29:@10094.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7)
  );
  StickySelects_2 StickySelects_7 ( // @[MemPrimitives.scala 121:29:@10166.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7)
  );
  StickySelects StickySelects_8 ( // @[MemPrimitives.scala 121:29:@10226.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3)
  );
  StickySelects StickySelects_9 ( // @[MemPrimitives.scala 121:29:@10266.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3)
  );
  StickySelects_2 StickySelects_10 ( // @[MemPrimitives.scala 121:29:@10318.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7)
  );
  StickySelects_2 StickySelects_11 ( // @[MemPrimitives.scala 121:29:@10390.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7)
  );
  StickySelects StickySelects_12 ( // @[MemPrimitives.scala 121:29:@10450.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3)
  );
  StickySelects StickySelects_13 ( // @[MemPrimitives.scala 121:29:@10490.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3)
  );
  StickySelects_2 StickySelects_14 ( // @[MemPrimitives.scala 121:29:@10542.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_ins_6(StickySelects_14_io_ins_6),
    .io_ins_7(StickySelects_14_io_ins_7),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5),
    .io_outs_6(StickySelects_14_io_outs_6),
    .io_outs_7(StickySelects_14_io_outs_7)
  );
  StickySelects_2 StickySelects_15 ( // @[MemPrimitives.scala 121:29:@10614.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_ins_6(StickySelects_15_io_ins_6),
    .io_ins_7(StickySelects_15_io_ins_7),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5),
    .io_outs_6(StickySelects_15_io_outs_6),
    .io_outs_7(StickySelects_15_io_outs_7)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@10675.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_1 ( // @[package.scala 93:22:@10683.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_2 ( // @[package.scala 93:22:@10691.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_3 ( // @[package.scala 93:22:@10699.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_4 ( // @[package.scala 93:22:@10723.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_5 ( // @[package.scala 93:22:@10731.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_6 ( // @[package.scala 93:22:@10739.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_7 ( // @[package.scala 93:22:@10747.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_8 ( // @[package.scala 93:22:@10771.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_9 ( // @[package.scala 93:22:@10779.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_10 ( // @[package.scala 93:22:@10787.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_11 ( // @[package.scala 93:22:@10795.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_12 ( // @[package.scala 93:22:@10819.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_13 ( // @[package.scala 93:22:@10827.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_14 ( // @[package.scala 93:22:@10835.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_15 ( // @[package.scala 93:22:@10843.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_16 ( // @[package.scala 93:22:@10867.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_17 ( // @[package.scala 93:22:@10875.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_18 ( // @[package.scala 93:22:@10883.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_19 ( // @[package.scala 93:22:@10891.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_20 ( // @[package.scala 93:22:@10915.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_21 ( // @[package.scala 93:22:@10923.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_22 ( // @[package.scala 93:22:@10931.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_23 ( // @[package.scala 93:22:@10939.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_24 ( // @[package.scala 93:22:@10963.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_25 ( // @[package.scala 93:22:@10971.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_26 ( // @[package.scala 93:22:@10979.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_27 ( // @[package.scala 93:22:@10987.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_28 ( // @[package.scala 93:22:@11011.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_29 ( // @[package.scala 93:22:@11019.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_30 ( // @[package.scala 93:22:@11027.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_31 ( // @[package.scala 93:22:@11035.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_32 ( // @[package.scala 93:22:@11059.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_33 ( // @[package.scala 93:22:@11067.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_34 ( // @[package.scala 93:22:@11075.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_35 ( // @[package.scala 93:22:@11083.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_36 ( // @[package.scala 93:22:@11107.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_37 ( // @[package.scala 93:22:@11115.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_38 ( // @[package.scala 93:22:@11123.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_39 ( // @[package.scala 93:22:@11131.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_40 ( // @[package.scala 93:22:@11155.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_41 ( // @[package.scala 93:22:@11163.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_42 ( // @[package.scala 93:22:@11171.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_43 ( // @[package.scala 93:22:@11179.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_44 ( // @[package.scala 93:22:@11203.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_45 ( // @[package.scala 93:22:@11211.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_46 ( // @[package.scala 93:22:@11219.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_47 ( // @[package.scala 93:22:@11227.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_48 ( // @[package.scala 93:22:@11251.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_49 ( // @[package.scala 93:22:@11259.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_50 ( // @[package.scala 93:22:@11267.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_51 ( // @[package.scala 93:22:@11275.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_52 ( // @[package.scala 93:22:@11299.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_53 ( // @[package.scala 93:22:@11307.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_54 ( // @[package.scala 93:22:@11315.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_55 ( // @[package.scala 93:22:@11323.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_56 ( // @[package.scala 93:22:@11347.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_57 ( // @[package.scala 93:22:@11355.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_58 ( // @[package.scala 93:22:@11363.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_59 ( // @[package.scala 93:22:@11371.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_60 ( // @[package.scala 93:22:@11395.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_61 ( // @[package.scala 93:22:@11403.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_62 ( // @[package.scala 93:22:@11411.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_63 ( // @[package.scala 93:22:@11419.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_64 ( // @[package.scala 93:22:@11443.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_65 ( // @[package.scala 93:22:@11451.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_66 ( // @[package.scala 93:22:@11459.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_67 ( // @[package.scala 93:22:@11467.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_68 ( // @[package.scala 93:22:@11491.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_69 ( // @[package.scala 93:22:@11499.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_70 ( // @[package.scala 93:22:@11507.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_71 ( // @[package.scala 93:22:@11515.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_72 ( // @[package.scala 93:22:@11539.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_73 ( // @[package.scala 93:22:@11547.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_74 ( // @[package.scala 93:22:@11555.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_75 ( // @[package.scala 93:22:@11563.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_76 ( // @[package.scala 93:22:@11587.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_77 ( // @[package.scala 93:22:@11595.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_78 ( // @[package.scala 93:22:@11603.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_79 ( // @[package.scala 93:22:@11611.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_80 ( // @[package.scala 93:22:@11635.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_81 ( // @[package.scala 93:22:@11643.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_82 ( // @[package.scala 93:22:@11651.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_83 ( // @[package.scala 93:22:@11659.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_84 ( // @[package.scala 93:22:@11683.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_85 ( // @[package.scala 93:22:@11691.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_86 ( // @[package.scala 93:22:@11699.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_87 ( // @[package.scala 93:22:@11707.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_88 ( // @[package.scala 93:22:@11731.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_89 ( // @[package.scala 93:22:@11739.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_90 ( // @[package.scala 93:22:@11747.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_91 ( // @[package.scala 93:22:@11755.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_92 ( // @[package.scala 93:22:@11779.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_93 ( // @[package.scala 93:22:@11787.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_94 ( // @[package.scala 93:22:@11795.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_95 ( // @[package.scala 93:22:@11803.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  assign _T_1032 = io_wPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9494.4]
  assign _T_1035 = io_wPort_3_en_0 & _T_1032; // @[MemPrimitives.scala 83:102:@9496.4]
  assign _T_1037 = io_wPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9497.4]
  assign _T_1040 = io_wPort_4_en_0 & _T_1037; // @[MemPrimitives.scala 83:102:@9499.4]
  assign _T_1042 = {_T_1035,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@9501.4]
  assign _T_1044 = {_T_1040,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@9503.4]
  assign _T_1045 = _T_1035 ? _T_1042 : _T_1044; // @[Mux.scala 31:69:@9504.4]
  assign _T_1050 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9511.4]
  assign _T_1053 = io_wPort_0_en_0 & _T_1050; // @[MemPrimitives.scala 83:102:@9513.4]
  assign _T_1055 = io_wPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9514.4]
  assign _T_1058 = io_wPort_2_en_0 & _T_1055; // @[MemPrimitives.scala 83:102:@9516.4]
  assign _T_1060 = {_T_1053,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9518.4]
  assign _T_1062 = {_T_1058,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@9520.4]
  assign _T_1063 = _T_1053 ? _T_1060 : _T_1062; // @[Mux.scala 31:69:@9521.4]
  assign _T_1068 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9528.4]
  assign _T_1071 = io_wPort_1_en_0 & _T_1068; // @[MemPrimitives.scala 83:102:@9530.4]
  assign _T_1073 = io_wPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9531.4]
  assign _T_1076 = io_wPort_7_en_0 & _T_1073; // @[MemPrimitives.scala 83:102:@9533.4]
  assign _T_1078 = {_T_1071,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9535.4]
  assign _T_1080 = {_T_1076,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@9537.4]
  assign _T_1081 = _T_1071 ? _T_1078 : _T_1080; // @[Mux.scala 31:69:@9538.4]
  assign _T_1086 = io_wPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9545.4]
  assign _T_1089 = io_wPort_5_en_0 & _T_1086; // @[MemPrimitives.scala 83:102:@9547.4]
  assign _T_1091 = io_wPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9548.4]
  assign _T_1094 = io_wPort_6_en_0 & _T_1091; // @[MemPrimitives.scala 83:102:@9550.4]
  assign _T_1096 = {_T_1089,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@9552.4]
  assign _T_1098 = {_T_1094,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@9554.4]
  assign _T_1099 = _T_1089 ? _T_1096 : _T_1098; // @[Mux.scala 31:69:@9555.4]
  assign _T_1104 = io_wPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9562.4]
  assign _T_1107 = io_wPort_3_en_0 & _T_1104; // @[MemPrimitives.scala 83:102:@9564.4]
  assign _T_1109 = io_wPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9565.4]
  assign _T_1112 = io_wPort_4_en_0 & _T_1109; // @[MemPrimitives.scala 83:102:@9567.4]
  assign _T_1114 = {_T_1107,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@9569.4]
  assign _T_1116 = {_T_1112,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@9571.4]
  assign _T_1117 = _T_1107 ? _T_1114 : _T_1116; // @[Mux.scala 31:69:@9572.4]
  assign _T_1122 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9579.4]
  assign _T_1125 = io_wPort_0_en_0 & _T_1122; // @[MemPrimitives.scala 83:102:@9581.4]
  assign _T_1127 = io_wPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9582.4]
  assign _T_1130 = io_wPort_2_en_0 & _T_1127; // @[MemPrimitives.scala 83:102:@9584.4]
  assign _T_1132 = {_T_1125,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9586.4]
  assign _T_1134 = {_T_1130,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@9588.4]
  assign _T_1135 = _T_1125 ? _T_1132 : _T_1134; // @[Mux.scala 31:69:@9589.4]
  assign _T_1140 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9596.4]
  assign _T_1143 = io_wPort_1_en_0 & _T_1140; // @[MemPrimitives.scala 83:102:@9598.4]
  assign _T_1145 = io_wPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9599.4]
  assign _T_1148 = io_wPort_7_en_0 & _T_1145; // @[MemPrimitives.scala 83:102:@9601.4]
  assign _T_1150 = {_T_1143,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9603.4]
  assign _T_1152 = {_T_1148,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@9605.4]
  assign _T_1153 = _T_1143 ? _T_1150 : _T_1152; // @[Mux.scala 31:69:@9606.4]
  assign _T_1158 = io_wPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9613.4]
  assign _T_1161 = io_wPort_5_en_0 & _T_1158; // @[MemPrimitives.scala 83:102:@9615.4]
  assign _T_1163 = io_wPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9616.4]
  assign _T_1166 = io_wPort_6_en_0 & _T_1163; // @[MemPrimitives.scala 83:102:@9618.4]
  assign _T_1168 = {_T_1161,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@9620.4]
  assign _T_1170 = {_T_1166,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@9622.4]
  assign _T_1171 = _T_1161 ? _T_1168 : _T_1170; // @[Mux.scala 31:69:@9623.4]
  assign _T_1176 = io_wPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9630.4]
  assign _T_1179 = io_wPort_3_en_0 & _T_1176; // @[MemPrimitives.scala 83:102:@9632.4]
  assign _T_1181 = io_wPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9633.4]
  assign _T_1184 = io_wPort_4_en_0 & _T_1181; // @[MemPrimitives.scala 83:102:@9635.4]
  assign _T_1186 = {_T_1179,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@9637.4]
  assign _T_1188 = {_T_1184,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@9639.4]
  assign _T_1189 = _T_1179 ? _T_1186 : _T_1188; // @[Mux.scala 31:69:@9640.4]
  assign _T_1194 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9647.4]
  assign _T_1197 = io_wPort_0_en_0 & _T_1194; // @[MemPrimitives.scala 83:102:@9649.4]
  assign _T_1199 = io_wPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9650.4]
  assign _T_1202 = io_wPort_2_en_0 & _T_1199; // @[MemPrimitives.scala 83:102:@9652.4]
  assign _T_1204 = {_T_1197,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9654.4]
  assign _T_1206 = {_T_1202,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@9656.4]
  assign _T_1207 = _T_1197 ? _T_1204 : _T_1206; // @[Mux.scala 31:69:@9657.4]
  assign _T_1212 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9664.4]
  assign _T_1215 = io_wPort_1_en_0 & _T_1212; // @[MemPrimitives.scala 83:102:@9666.4]
  assign _T_1217 = io_wPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9667.4]
  assign _T_1220 = io_wPort_7_en_0 & _T_1217; // @[MemPrimitives.scala 83:102:@9669.4]
  assign _T_1222 = {_T_1215,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9671.4]
  assign _T_1224 = {_T_1220,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@9673.4]
  assign _T_1225 = _T_1215 ? _T_1222 : _T_1224; // @[Mux.scala 31:69:@9674.4]
  assign _T_1230 = io_wPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9681.4]
  assign _T_1233 = io_wPort_5_en_0 & _T_1230; // @[MemPrimitives.scala 83:102:@9683.4]
  assign _T_1235 = io_wPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9684.4]
  assign _T_1238 = io_wPort_6_en_0 & _T_1235; // @[MemPrimitives.scala 83:102:@9686.4]
  assign _T_1240 = {_T_1233,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@9688.4]
  assign _T_1242 = {_T_1238,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@9690.4]
  assign _T_1243 = _T_1233 ? _T_1240 : _T_1242; // @[Mux.scala 31:69:@9691.4]
  assign _T_1248 = io_wPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9698.4]
  assign _T_1251 = io_wPort_3_en_0 & _T_1248; // @[MemPrimitives.scala 83:102:@9700.4]
  assign _T_1253 = io_wPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9701.4]
  assign _T_1256 = io_wPort_4_en_0 & _T_1253; // @[MemPrimitives.scala 83:102:@9703.4]
  assign _T_1258 = {_T_1251,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@9705.4]
  assign _T_1260 = {_T_1256,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@9707.4]
  assign _T_1261 = _T_1251 ? _T_1258 : _T_1260; // @[Mux.scala 31:69:@9708.4]
  assign _T_1266 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9715.4]
  assign _T_1269 = io_wPort_0_en_0 & _T_1266; // @[MemPrimitives.scala 83:102:@9717.4]
  assign _T_1271 = io_wPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9718.4]
  assign _T_1274 = io_wPort_2_en_0 & _T_1271; // @[MemPrimitives.scala 83:102:@9720.4]
  assign _T_1276 = {_T_1269,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9722.4]
  assign _T_1278 = {_T_1274,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@9724.4]
  assign _T_1279 = _T_1269 ? _T_1276 : _T_1278; // @[Mux.scala 31:69:@9725.4]
  assign _T_1284 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9732.4]
  assign _T_1287 = io_wPort_1_en_0 & _T_1284; // @[MemPrimitives.scala 83:102:@9734.4]
  assign _T_1289 = io_wPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9735.4]
  assign _T_1292 = io_wPort_7_en_0 & _T_1289; // @[MemPrimitives.scala 83:102:@9737.4]
  assign _T_1294 = {_T_1287,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9739.4]
  assign _T_1296 = {_T_1292,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@9741.4]
  assign _T_1297 = _T_1287 ? _T_1294 : _T_1296; // @[Mux.scala 31:69:@9742.4]
  assign _T_1302 = io_wPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9749.4]
  assign _T_1305 = io_wPort_5_en_0 & _T_1302; // @[MemPrimitives.scala 83:102:@9751.4]
  assign _T_1307 = io_wPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9752.4]
  assign _T_1310 = io_wPort_6_en_0 & _T_1307; // @[MemPrimitives.scala 83:102:@9754.4]
  assign _T_1312 = {_T_1305,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@9756.4]
  assign _T_1314 = {_T_1310,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@9758.4]
  assign _T_1315 = _T_1305 ? _T_1312 : _T_1314; // @[Mux.scala 31:69:@9759.4]
  assign _T_1320 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9766.4]
  assign _T_1325 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9769.4]
  assign _T_1330 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9772.4]
  assign _T_1335 = io_rPort_20_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9775.4]
  assign _T_1339 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@9785.4]
  assign _T_1340 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@9786.4]
  assign _T_1341 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@9787.4]
  assign _T_1342 = StickySelects_io_outs_3; // @[MemPrimitives.scala 123:41:@9788.4]
  assign _T_1344 = {_T_1339,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9790.4]
  assign _T_1346 = {_T_1340,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9792.4]
  assign _T_1348 = {_T_1341,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9794.4]
  assign _T_1350 = {_T_1342,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@9796.4]
  assign _T_1351 = _T_1341 ? _T_1348 : _T_1350; // @[Mux.scala 31:69:@9797.4]
  assign _T_1352 = _T_1340 ? _T_1346 : _T_1351; // @[Mux.scala 31:69:@9798.4]
  assign _T_1353 = _T_1339 ? _T_1344 : _T_1352; // @[Mux.scala 31:69:@9799.4]
  assign _T_1358 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9806.4]
  assign _T_1363 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9809.4]
  assign _T_1368 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9812.4]
  assign _T_1373 = io_rPort_21_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9815.4]
  assign _T_1377 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@9825.4]
  assign _T_1378 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@9826.4]
  assign _T_1379 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@9827.4]
  assign _T_1380 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 123:41:@9828.4]
  assign _T_1382 = {_T_1377,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9830.4]
  assign _T_1384 = {_T_1378,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9832.4]
  assign _T_1386 = {_T_1379,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9834.4]
  assign _T_1388 = {_T_1380,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@9836.4]
  assign _T_1389 = _T_1379 ? _T_1386 : _T_1388; // @[Mux.scala 31:69:@9837.4]
  assign _T_1390 = _T_1378 ? _T_1384 : _T_1389; // @[Mux.scala 31:69:@9838.4]
  assign _T_1391 = _T_1377 ? _T_1382 : _T_1390; // @[Mux.scala 31:69:@9839.4]
  assign _T_1396 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9846.4]
  assign _T_1401 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9849.4]
  assign _T_1406 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9852.4]
  assign _T_1411 = io_rPort_13_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9855.4]
  assign _T_1416 = io_rPort_15_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9858.4]
  assign _T_1421 = io_rPort_17_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9861.4]
  assign _T_1426 = io_rPort_22_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9864.4]
  assign _T_1431 = io_rPort_23_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9867.4]
  assign _T_1435 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@9881.4]
  assign _T_1436 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@9882.4]
  assign _T_1437 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@9883.4]
  assign _T_1438 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 123:41:@9884.4]
  assign _T_1439 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 123:41:@9885.4]
  assign _T_1440 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 123:41:@9886.4]
  assign _T_1441 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 123:41:@9887.4]
  assign _T_1442 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 123:41:@9888.4]
  assign _T_1444 = {_T_1435,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9890.4]
  assign _T_1446 = {_T_1436,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9892.4]
  assign _T_1448 = {_T_1437,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9894.4]
  assign _T_1450 = {_T_1438,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@9896.4]
  assign _T_1452 = {_T_1439,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@9898.4]
  assign _T_1454 = {_T_1440,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@9900.4]
  assign _T_1456 = {_T_1441,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@9902.4]
  assign _T_1458 = {_T_1442,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@9904.4]
  assign _T_1459 = _T_1441 ? _T_1456 : _T_1458; // @[Mux.scala 31:69:@9905.4]
  assign _T_1460 = _T_1440 ? _T_1454 : _T_1459; // @[Mux.scala 31:69:@9906.4]
  assign _T_1461 = _T_1439 ? _T_1452 : _T_1460; // @[Mux.scala 31:69:@9907.4]
  assign _T_1462 = _T_1438 ? _T_1450 : _T_1461; // @[Mux.scala 31:69:@9908.4]
  assign _T_1463 = _T_1437 ? _T_1448 : _T_1462; // @[Mux.scala 31:69:@9909.4]
  assign _T_1464 = _T_1436 ? _T_1446 : _T_1463; // @[Mux.scala 31:69:@9910.4]
  assign _T_1465 = _T_1435 ? _T_1444 : _T_1464; // @[Mux.scala 31:69:@9911.4]
  assign _T_1470 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9918.4]
  assign _T_1475 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9921.4]
  assign _T_1480 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9924.4]
  assign _T_1485 = io_rPort_12_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9927.4]
  assign _T_1490 = io_rPort_14_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9930.4]
  assign _T_1495 = io_rPort_16_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9933.4]
  assign _T_1500 = io_rPort_18_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9936.4]
  assign _T_1505 = io_rPort_19_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9939.4]
  assign _T_1509 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@9953.4]
  assign _T_1510 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@9954.4]
  assign _T_1511 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@9955.4]
  assign _T_1512 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@9956.4]
  assign _T_1513 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@9957.4]
  assign _T_1514 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@9958.4]
  assign _T_1515 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 123:41:@9959.4]
  assign _T_1516 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 123:41:@9960.4]
  assign _T_1518 = {_T_1509,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9962.4]
  assign _T_1520 = {_T_1510,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9964.4]
  assign _T_1522 = {_T_1511,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9966.4]
  assign _T_1524 = {_T_1512,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@9968.4]
  assign _T_1526 = {_T_1513,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@9970.4]
  assign _T_1528 = {_T_1514,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@9972.4]
  assign _T_1530 = {_T_1515,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@9974.4]
  assign _T_1532 = {_T_1516,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@9976.4]
  assign _T_1533 = _T_1515 ? _T_1530 : _T_1532; // @[Mux.scala 31:69:@9977.4]
  assign _T_1534 = _T_1514 ? _T_1528 : _T_1533; // @[Mux.scala 31:69:@9978.4]
  assign _T_1535 = _T_1513 ? _T_1526 : _T_1534; // @[Mux.scala 31:69:@9979.4]
  assign _T_1536 = _T_1512 ? _T_1524 : _T_1535; // @[Mux.scala 31:69:@9980.4]
  assign _T_1537 = _T_1511 ? _T_1522 : _T_1536; // @[Mux.scala 31:69:@9981.4]
  assign _T_1538 = _T_1510 ? _T_1520 : _T_1537; // @[Mux.scala 31:69:@9982.4]
  assign _T_1539 = _T_1509 ? _T_1518 : _T_1538; // @[Mux.scala 31:69:@9983.4]
  assign _T_1544 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9990.4]
  assign _T_1549 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9993.4]
  assign _T_1554 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9996.4]
  assign _T_1559 = io_rPort_20_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9999.4]
  assign _T_1563 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@10009.4]
  assign _T_1564 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@10010.4]
  assign _T_1565 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@10011.4]
  assign _T_1566 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 123:41:@10012.4]
  assign _T_1568 = {_T_1563,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10014.4]
  assign _T_1570 = {_T_1564,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10016.4]
  assign _T_1572 = {_T_1565,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10018.4]
  assign _T_1574 = {_T_1566,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@10020.4]
  assign _T_1575 = _T_1565 ? _T_1572 : _T_1574; // @[Mux.scala 31:69:@10021.4]
  assign _T_1576 = _T_1564 ? _T_1570 : _T_1575; // @[Mux.scala 31:69:@10022.4]
  assign _T_1577 = _T_1563 ? _T_1568 : _T_1576; // @[Mux.scala 31:69:@10023.4]
  assign _T_1582 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10030.4]
  assign _T_1587 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10033.4]
  assign _T_1592 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10036.4]
  assign _T_1597 = io_rPort_21_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10039.4]
  assign _T_1601 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@10049.4]
  assign _T_1602 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@10050.4]
  assign _T_1603 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@10051.4]
  assign _T_1604 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 123:41:@10052.4]
  assign _T_1606 = {_T_1601,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10054.4]
  assign _T_1608 = {_T_1602,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10056.4]
  assign _T_1610 = {_T_1603,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10058.4]
  assign _T_1612 = {_T_1604,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@10060.4]
  assign _T_1613 = _T_1603 ? _T_1610 : _T_1612; // @[Mux.scala 31:69:@10061.4]
  assign _T_1614 = _T_1602 ? _T_1608 : _T_1613; // @[Mux.scala 31:69:@10062.4]
  assign _T_1615 = _T_1601 ? _T_1606 : _T_1614; // @[Mux.scala 31:69:@10063.4]
  assign _T_1620 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10070.4]
  assign _T_1625 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10073.4]
  assign _T_1630 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10076.4]
  assign _T_1635 = io_rPort_13_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10079.4]
  assign _T_1640 = io_rPort_15_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10082.4]
  assign _T_1645 = io_rPort_17_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10085.4]
  assign _T_1650 = io_rPort_22_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10088.4]
  assign _T_1655 = io_rPort_23_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10091.4]
  assign _T_1659 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@10105.4]
  assign _T_1660 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@10106.4]
  assign _T_1661 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@10107.4]
  assign _T_1662 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 123:41:@10108.4]
  assign _T_1663 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 123:41:@10109.4]
  assign _T_1664 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 123:41:@10110.4]
  assign _T_1665 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 123:41:@10111.4]
  assign _T_1666 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 123:41:@10112.4]
  assign _T_1668 = {_T_1659,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10114.4]
  assign _T_1670 = {_T_1660,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10116.4]
  assign _T_1672 = {_T_1661,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10118.4]
  assign _T_1674 = {_T_1662,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@10120.4]
  assign _T_1676 = {_T_1663,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@10122.4]
  assign _T_1678 = {_T_1664,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@10124.4]
  assign _T_1680 = {_T_1665,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@10126.4]
  assign _T_1682 = {_T_1666,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@10128.4]
  assign _T_1683 = _T_1665 ? _T_1680 : _T_1682; // @[Mux.scala 31:69:@10129.4]
  assign _T_1684 = _T_1664 ? _T_1678 : _T_1683; // @[Mux.scala 31:69:@10130.4]
  assign _T_1685 = _T_1663 ? _T_1676 : _T_1684; // @[Mux.scala 31:69:@10131.4]
  assign _T_1686 = _T_1662 ? _T_1674 : _T_1685; // @[Mux.scala 31:69:@10132.4]
  assign _T_1687 = _T_1661 ? _T_1672 : _T_1686; // @[Mux.scala 31:69:@10133.4]
  assign _T_1688 = _T_1660 ? _T_1670 : _T_1687; // @[Mux.scala 31:69:@10134.4]
  assign _T_1689 = _T_1659 ? _T_1668 : _T_1688; // @[Mux.scala 31:69:@10135.4]
  assign _T_1694 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10142.4]
  assign _T_1699 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10145.4]
  assign _T_1704 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10148.4]
  assign _T_1709 = io_rPort_12_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10151.4]
  assign _T_1714 = io_rPort_14_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10154.4]
  assign _T_1719 = io_rPort_16_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10157.4]
  assign _T_1724 = io_rPort_18_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10160.4]
  assign _T_1729 = io_rPort_19_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10163.4]
  assign _T_1733 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@10177.4]
  assign _T_1734 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@10178.4]
  assign _T_1735 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@10179.4]
  assign _T_1736 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@10180.4]
  assign _T_1737 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@10181.4]
  assign _T_1738 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@10182.4]
  assign _T_1739 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 123:41:@10183.4]
  assign _T_1740 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 123:41:@10184.4]
  assign _T_1742 = {_T_1733,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10186.4]
  assign _T_1744 = {_T_1734,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10188.4]
  assign _T_1746 = {_T_1735,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10190.4]
  assign _T_1748 = {_T_1736,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@10192.4]
  assign _T_1750 = {_T_1737,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@10194.4]
  assign _T_1752 = {_T_1738,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@10196.4]
  assign _T_1754 = {_T_1739,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@10198.4]
  assign _T_1756 = {_T_1740,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@10200.4]
  assign _T_1757 = _T_1739 ? _T_1754 : _T_1756; // @[Mux.scala 31:69:@10201.4]
  assign _T_1758 = _T_1738 ? _T_1752 : _T_1757; // @[Mux.scala 31:69:@10202.4]
  assign _T_1759 = _T_1737 ? _T_1750 : _T_1758; // @[Mux.scala 31:69:@10203.4]
  assign _T_1760 = _T_1736 ? _T_1748 : _T_1759; // @[Mux.scala 31:69:@10204.4]
  assign _T_1761 = _T_1735 ? _T_1746 : _T_1760; // @[Mux.scala 31:69:@10205.4]
  assign _T_1762 = _T_1734 ? _T_1744 : _T_1761; // @[Mux.scala 31:69:@10206.4]
  assign _T_1763 = _T_1733 ? _T_1742 : _T_1762; // @[Mux.scala 31:69:@10207.4]
  assign _T_1768 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10214.4]
  assign _T_1773 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10217.4]
  assign _T_1778 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10220.4]
  assign _T_1783 = io_rPort_20_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10223.4]
  assign _T_1787 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@10233.4]
  assign _T_1788 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@10234.4]
  assign _T_1789 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@10235.4]
  assign _T_1790 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 123:41:@10236.4]
  assign _T_1792 = {_T_1787,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10238.4]
  assign _T_1794 = {_T_1788,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10240.4]
  assign _T_1796 = {_T_1789,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10242.4]
  assign _T_1798 = {_T_1790,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@10244.4]
  assign _T_1799 = _T_1789 ? _T_1796 : _T_1798; // @[Mux.scala 31:69:@10245.4]
  assign _T_1800 = _T_1788 ? _T_1794 : _T_1799; // @[Mux.scala 31:69:@10246.4]
  assign _T_1801 = _T_1787 ? _T_1792 : _T_1800; // @[Mux.scala 31:69:@10247.4]
  assign _T_1806 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10254.4]
  assign _T_1811 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10257.4]
  assign _T_1816 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10260.4]
  assign _T_1821 = io_rPort_21_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10263.4]
  assign _T_1825 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@10273.4]
  assign _T_1826 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@10274.4]
  assign _T_1827 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@10275.4]
  assign _T_1828 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 123:41:@10276.4]
  assign _T_1830 = {_T_1825,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10278.4]
  assign _T_1832 = {_T_1826,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10280.4]
  assign _T_1834 = {_T_1827,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10282.4]
  assign _T_1836 = {_T_1828,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@10284.4]
  assign _T_1837 = _T_1827 ? _T_1834 : _T_1836; // @[Mux.scala 31:69:@10285.4]
  assign _T_1838 = _T_1826 ? _T_1832 : _T_1837; // @[Mux.scala 31:69:@10286.4]
  assign _T_1839 = _T_1825 ? _T_1830 : _T_1838; // @[Mux.scala 31:69:@10287.4]
  assign _T_1844 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10294.4]
  assign _T_1849 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10297.4]
  assign _T_1854 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10300.4]
  assign _T_1859 = io_rPort_13_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10303.4]
  assign _T_1864 = io_rPort_15_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10306.4]
  assign _T_1869 = io_rPort_17_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10309.4]
  assign _T_1874 = io_rPort_22_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10312.4]
  assign _T_1879 = io_rPort_23_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10315.4]
  assign _T_1883 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@10329.4]
  assign _T_1884 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@10330.4]
  assign _T_1885 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@10331.4]
  assign _T_1886 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 123:41:@10332.4]
  assign _T_1887 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 123:41:@10333.4]
  assign _T_1888 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 123:41:@10334.4]
  assign _T_1889 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 123:41:@10335.4]
  assign _T_1890 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 123:41:@10336.4]
  assign _T_1892 = {_T_1883,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10338.4]
  assign _T_1894 = {_T_1884,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10340.4]
  assign _T_1896 = {_T_1885,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10342.4]
  assign _T_1898 = {_T_1886,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@10344.4]
  assign _T_1900 = {_T_1887,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@10346.4]
  assign _T_1902 = {_T_1888,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@10348.4]
  assign _T_1904 = {_T_1889,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@10350.4]
  assign _T_1906 = {_T_1890,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@10352.4]
  assign _T_1907 = _T_1889 ? _T_1904 : _T_1906; // @[Mux.scala 31:69:@10353.4]
  assign _T_1908 = _T_1888 ? _T_1902 : _T_1907; // @[Mux.scala 31:69:@10354.4]
  assign _T_1909 = _T_1887 ? _T_1900 : _T_1908; // @[Mux.scala 31:69:@10355.4]
  assign _T_1910 = _T_1886 ? _T_1898 : _T_1909; // @[Mux.scala 31:69:@10356.4]
  assign _T_1911 = _T_1885 ? _T_1896 : _T_1910; // @[Mux.scala 31:69:@10357.4]
  assign _T_1912 = _T_1884 ? _T_1894 : _T_1911; // @[Mux.scala 31:69:@10358.4]
  assign _T_1913 = _T_1883 ? _T_1892 : _T_1912; // @[Mux.scala 31:69:@10359.4]
  assign _T_1918 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10366.4]
  assign _T_1923 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10369.4]
  assign _T_1928 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10372.4]
  assign _T_1933 = io_rPort_12_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10375.4]
  assign _T_1938 = io_rPort_14_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10378.4]
  assign _T_1943 = io_rPort_16_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10381.4]
  assign _T_1948 = io_rPort_18_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10384.4]
  assign _T_1953 = io_rPort_19_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10387.4]
  assign _T_1957 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@10401.4]
  assign _T_1958 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@10402.4]
  assign _T_1959 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@10403.4]
  assign _T_1960 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@10404.4]
  assign _T_1961 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@10405.4]
  assign _T_1962 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@10406.4]
  assign _T_1963 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 123:41:@10407.4]
  assign _T_1964 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 123:41:@10408.4]
  assign _T_1966 = {_T_1957,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10410.4]
  assign _T_1968 = {_T_1958,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10412.4]
  assign _T_1970 = {_T_1959,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10414.4]
  assign _T_1972 = {_T_1960,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@10416.4]
  assign _T_1974 = {_T_1961,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@10418.4]
  assign _T_1976 = {_T_1962,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@10420.4]
  assign _T_1978 = {_T_1963,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@10422.4]
  assign _T_1980 = {_T_1964,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@10424.4]
  assign _T_1981 = _T_1963 ? _T_1978 : _T_1980; // @[Mux.scala 31:69:@10425.4]
  assign _T_1982 = _T_1962 ? _T_1976 : _T_1981; // @[Mux.scala 31:69:@10426.4]
  assign _T_1983 = _T_1961 ? _T_1974 : _T_1982; // @[Mux.scala 31:69:@10427.4]
  assign _T_1984 = _T_1960 ? _T_1972 : _T_1983; // @[Mux.scala 31:69:@10428.4]
  assign _T_1985 = _T_1959 ? _T_1970 : _T_1984; // @[Mux.scala 31:69:@10429.4]
  assign _T_1986 = _T_1958 ? _T_1968 : _T_1985; // @[Mux.scala 31:69:@10430.4]
  assign _T_1987 = _T_1957 ? _T_1966 : _T_1986; // @[Mux.scala 31:69:@10431.4]
  assign _T_1992 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10438.4]
  assign _T_1997 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10441.4]
  assign _T_2002 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10444.4]
  assign _T_2007 = io_rPort_20_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10447.4]
  assign _T_2011 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@10457.4]
  assign _T_2012 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@10458.4]
  assign _T_2013 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 123:41:@10459.4]
  assign _T_2014 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 123:41:@10460.4]
  assign _T_2016 = {_T_2011,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10462.4]
  assign _T_2018 = {_T_2012,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10464.4]
  assign _T_2020 = {_T_2013,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10466.4]
  assign _T_2022 = {_T_2014,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@10468.4]
  assign _T_2023 = _T_2013 ? _T_2020 : _T_2022; // @[Mux.scala 31:69:@10469.4]
  assign _T_2024 = _T_2012 ? _T_2018 : _T_2023; // @[Mux.scala 31:69:@10470.4]
  assign _T_2025 = _T_2011 ? _T_2016 : _T_2024; // @[Mux.scala 31:69:@10471.4]
  assign _T_2030 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10478.4]
  assign _T_2035 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10481.4]
  assign _T_2040 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10484.4]
  assign _T_2045 = io_rPort_21_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10487.4]
  assign _T_2049 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@10497.4]
  assign _T_2050 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@10498.4]
  assign _T_2051 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 123:41:@10499.4]
  assign _T_2052 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 123:41:@10500.4]
  assign _T_2054 = {_T_2049,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10502.4]
  assign _T_2056 = {_T_2050,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10504.4]
  assign _T_2058 = {_T_2051,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10506.4]
  assign _T_2060 = {_T_2052,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@10508.4]
  assign _T_2061 = _T_2051 ? _T_2058 : _T_2060; // @[Mux.scala 31:69:@10509.4]
  assign _T_2062 = _T_2050 ? _T_2056 : _T_2061; // @[Mux.scala 31:69:@10510.4]
  assign _T_2063 = _T_2049 ? _T_2054 : _T_2062; // @[Mux.scala 31:69:@10511.4]
  assign _T_2068 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10518.4]
  assign _T_2073 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10521.4]
  assign _T_2078 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10524.4]
  assign _T_2083 = io_rPort_13_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10527.4]
  assign _T_2088 = io_rPort_15_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10530.4]
  assign _T_2093 = io_rPort_17_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10533.4]
  assign _T_2098 = io_rPort_22_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10536.4]
  assign _T_2103 = io_rPort_23_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10539.4]
  assign _T_2107 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@10553.4]
  assign _T_2108 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@10554.4]
  assign _T_2109 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 123:41:@10555.4]
  assign _T_2110 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 123:41:@10556.4]
  assign _T_2111 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 123:41:@10557.4]
  assign _T_2112 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 123:41:@10558.4]
  assign _T_2113 = StickySelects_14_io_outs_6; // @[MemPrimitives.scala 123:41:@10559.4]
  assign _T_2114 = StickySelects_14_io_outs_7; // @[MemPrimitives.scala 123:41:@10560.4]
  assign _T_2116 = {_T_2107,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10562.4]
  assign _T_2118 = {_T_2108,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10564.4]
  assign _T_2120 = {_T_2109,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10566.4]
  assign _T_2122 = {_T_2110,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@10568.4]
  assign _T_2124 = {_T_2111,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@10570.4]
  assign _T_2126 = {_T_2112,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@10572.4]
  assign _T_2128 = {_T_2113,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@10574.4]
  assign _T_2130 = {_T_2114,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@10576.4]
  assign _T_2131 = _T_2113 ? _T_2128 : _T_2130; // @[Mux.scala 31:69:@10577.4]
  assign _T_2132 = _T_2112 ? _T_2126 : _T_2131; // @[Mux.scala 31:69:@10578.4]
  assign _T_2133 = _T_2111 ? _T_2124 : _T_2132; // @[Mux.scala 31:69:@10579.4]
  assign _T_2134 = _T_2110 ? _T_2122 : _T_2133; // @[Mux.scala 31:69:@10580.4]
  assign _T_2135 = _T_2109 ? _T_2120 : _T_2134; // @[Mux.scala 31:69:@10581.4]
  assign _T_2136 = _T_2108 ? _T_2118 : _T_2135; // @[Mux.scala 31:69:@10582.4]
  assign _T_2137 = _T_2107 ? _T_2116 : _T_2136; // @[Mux.scala 31:69:@10583.4]
  assign _T_2142 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10590.4]
  assign _T_2147 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10593.4]
  assign _T_2152 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10596.4]
  assign _T_2157 = io_rPort_12_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10599.4]
  assign _T_2162 = io_rPort_14_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10602.4]
  assign _T_2167 = io_rPort_16_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10605.4]
  assign _T_2172 = io_rPort_18_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10608.4]
  assign _T_2177 = io_rPort_19_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10611.4]
  assign _T_2181 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@10625.4]
  assign _T_2182 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@10626.4]
  assign _T_2183 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@10627.4]
  assign _T_2184 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@10628.4]
  assign _T_2185 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 123:41:@10629.4]
  assign _T_2186 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 123:41:@10630.4]
  assign _T_2187 = StickySelects_15_io_outs_6; // @[MemPrimitives.scala 123:41:@10631.4]
  assign _T_2188 = StickySelects_15_io_outs_7; // @[MemPrimitives.scala 123:41:@10632.4]
  assign _T_2190 = {_T_2181,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10634.4]
  assign _T_2192 = {_T_2182,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10636.4]
  assign _T_2194 = {_T_2183,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10638.4]
  assign _T_2196 = {_T_2184,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@10640.4]
  assign _T_2198 = {_T_2185,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@10642.4]
  assign _T_2200 = {_T_2186,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@10644.4]
  assign _T_2202 = {_T_2187,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@10646.4]
  assign _T_2204 = {_T_2188,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@10648.4]
  assign _T_2205 = _T_2187 ? _T_2202 : _T_2204; // @[Mux.scala 31:69:@10649.4]
  assign _T_2206 = _T_2186 ? _T_2200 : _T_2205; // @[Mux.scala 31:69:@10650.4]
  assign _T_2207 = _T_2185 ? _T_2198 : _T_2206; // @[Mux.scala 31:69:@10651.4]
  assign _T_2208 = _T_2184 ? _T_2196 : _T_2207; // @[Mux.scala 31:69:@10652.4]
  assign _T_2209 = _T_2183 ? _T_2194 : _T_2208; // @[Mux.scala 31:69:@10653.4]
  assign _T_2210 = _T_2182 ? _T_2192 : _T_2209; // @[Mux.scala 31:69:@10654.4]
  assign _T_2211 = _T_2181 ? _T_2190 : _T_2210; // @[Mux.scala 31:69:@10655.4]
  assign _T_2243 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@10696.4 package.scala 96:25:@10697.4]
  assign _T_2247 = _T_2243 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@10706.4]
  assign _T_2240 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@10688.4 package.scala 96:25:@10689.4]
  assign _T_2248 = _T_2240 ? Mem1D_5_io_output : _T_2247; // @[Mux.scala 31:69:@10707.4]
  assign _T_2237 = RetimeWrapper_io_out; // @[package.scala 96:25:@10680.4 package.scala 96:25:@10681.4]
  assign _T_2278 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@10744.4 package.scala 96:25:@10745.4]
  assign _T_2282 = _T_2278 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@10754.4]
  assign _T_2275 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@10736.4 package.scala 96:25:@10737.4]
  assign _T_2283 = _T_2275 ? Mem1D_7_io_output : _T_2282; // @[Mux.scala 31:69:@10755.4]
  assign _T_2272 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@10728.4 package.scala 96:25:@10729.4]
  assign _T_2313 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@10792.4 package.scala 96:25:@10793.4]
  assign _T_2317 = _T_2313 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@10802.4]
  assign _T_2310 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@10784.4 package.scala 96:25:@10785.4]
  assign _T_2318 = _T_2310 ? Mem1D_6_io_output : _T_2317; // @[Mux.scala 31:69:@10803.4]
  assign _T_2307 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@10776.4 package.scala 96:25:@10777.4]
  assign _T_2348 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@10840.4 package.scala 96:25:@10841.4]
  assign _T_2352 = _T_2348 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@10850.4]
  assign _T_2345 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@10832.4 package.scala 96:25:@10833.4]
  assign _T_2353 = _T_2345 ? Mem1D_5_io_output : _T_2352; // @[Mux.scala 31:69:@10851.4]
  assign _T_2342 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@10824.4 package.scala 96:25:@10825.4]
  assign _T_2383 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@10888.4 package.scala 96:25:@10889.4]
  assign _T_2387 = _T_2383 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@10898.4]
  assign _T_2380 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@10880.4 package.scala 96:25:@10881.4]
  assign _T_2388 = _T_2380 ? Mem1D_6_io_output : _T_2387; // @[Mux.scala 31:69:@10899.4]
  assign _T_2377 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@10872.4 package.scala 96:25:@10873.4]
  assign _T_2418 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@10936.4 package.scala 96:25:@10937.4]
  assign _T_2422 = _T_2418 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@10946.4]
  assign _T_2415 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@10928.4 package.scala 96:25:@10929.4]
  assign _T_2423 = _T_2415 ? Mem1D_4_io_output : _T_2422; // @[Mux.scala 31:69:@10947.4]
  assign _T_2412 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@10920.4 package.scala 96:25:@10921.4]
  assign _T_2453 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@10984.4 package.scala 96:25:@10985.4]
  assign _T_2457 = _T_2453 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@10994.4]
  assign _T_2450 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@10976.4 package.scala 96:25:@10977.4]
  assign _T_2458 = _T_2450 ? Mem1D_5_io_output : _T_2457; // @[Mux.scala 31:69:@10995.4]
  assign _T_2447 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@10968.4 package.scala 96:25:@10969.4]
  assign _T_2488 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@11032.4 package.scala 96:25:@11033.4]
  assign _T_2492 = _T_2488 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@11042.4]
  assign _T_2485 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@11024.4 package.scala 96:25:@11025.4]
  assign _T_2493 = _T_2485 ? Mem1D_4_io_output : _T_2492; // @[Mux.scala 31:69:@11043.4]
  assign _T_2482 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@11016.4 package.scala 96:25:@11017.4]
  assign _T_2523 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@11080.4 package.scala 96:25:@11081.4]
  assign _T_2527 = _T_2523 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11090.4]
  assign _T_2520 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@11072.4 package.scala 96:25:@11073.4]
  assign _T_2528 = _T_2520 ? Mem1D_7_io_output : _T_2527; // @[Mux.scala 31:69:@11091.4]
  assign _T_2517 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@11064.4 package.scala 96:25:@11065.4]
  assign _T_2558 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@11128.4 package.scala 96:25:@11129.4]
  assign _T_2562 = _T_2558 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11138.4]
  assign _T_2555 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@11120.4 package.scala 96:25:@11121.4]
  assign _T_2563 = _T_2555 ? Mem1D_7_io_output : _T_2562; // @[Mux.scala 31:69:@11139.4]
  assign _T_2552 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@11112.4 package.scala 96:25:@11113.4]
  assign _T_2593 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@11176.4 package.scala 96:25:@11177.4]
  assign _T_2597 = _T_2593 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@11186.4]
  assign _T_2590 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@11168.4 package.scala 96:25:@11169.4]
  assign _T_2598 = _T_2590 ? Mem1D_4_io_output : _T_2597; // @[Mux.scala 31:69:@11187.4]
  assign _T_2587 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@11160.4 package.scala 96:25:@11161.4]
  assign _T_2628 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@11224.4 package.scala 96:25:@11225.4]
  assign _T_2632 = _T_2628 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11234.4]
  assign _T_2625 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@11216.4 package.scala 96:25:@11217.4]
  assign _T_2633 = _T_2625 ? Mem1D_6_io_output : _T_2632; // @[Mux.scala 31:69:@11235.4]
  assign _T_2622 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@11208.4 package.scala 96:25:@11209.4]
  assign _T_2663 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@11272.4 package.scala 96:25:@11273.4]
  assign _T_2667 = _T_2663 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11282.4]
  assign _T_2660 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@11264.4 package.scala 96:25:@11265.4]
  assign _T_2668 = _T_2660 ? Mem1D_7_io_output : _T_2667; // @[Mux.scala 31:69:@11283.4]
  assign _T_2657 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@11256.4 package.scala 96:25:@11257.4]
  assign _T_2698 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@11320.4 package.scala 96:25:@11321.4]
  assign _T_2702 = _T_2698 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11330.4]
  assign _T_2695 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@11312.4 package.scala 96:25:@11313.4]
  assign _T_2703 = _T_2695 ? Mem1D_6_io_output : _T_2702; // @[Mux.scala 31:69:@11331.4]
  assign _T_2692 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@11304.4 package.scala 96:25:@11305.4]
  assign _T_2733 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@11368.4 package.scala 96:25:@11369.4]
  assign _T_2737 = _T_2733 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11378.4]
  assign _T_2730 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@11360.4 package.scala 96:25:@11361.4]
  assign _T_2738 = _T_2730 ? Mem1D_7_io_output : _T_2737; // @[Mux.scala 31:69:@11379.4]
  assign _T_2727 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@11352.4 package.scala 96:25:@11353.4]
  assign _T_2768 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@11416.4 package.scala 96:25:@11417.4]
  assign _T_2772 = _T_2768 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11426.4]
  assign _T_2765 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@11408.4 package.scala 96:25:@11409.4]
  assign _T_2773 = _T_2765 ? Mem1D_6_io_output : _T_2772; // @[Mux.scala 31:69:@11427.4]
  assign _T_2762 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@11400.4 package.scala 96:25:@11401.4]
  assign _T_2803 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@11464.4 package.scala 96:25:@11465.4]
  assign _T_2807 = _T_2803 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11474.4]
  assign _T_2800 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@11456.4 package.scala 96:25:@11457.4]
  assign _T_2808 = _T_2800 ? Mem1D_7_io_output : _T_2807; // @[Mux.scala 31:69:@11475.4]
  assign _T_2797 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@11448.4 package.scala 96:25:@11449.4]
  assign _T_2838 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@11512.4 package.scala 96:25:@11513.4]
  assign _T_2842 = _T_2838 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11522.4]
  assign _T_2835 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@11504.4 package.scala 96:25:@11505.4]
  assign _T_2843 = _T_2835 ? Mem1D_6_io_output : _T_2842; // @[Mux.scala 31:69:@11523.4]
  assign _T_2832 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@11496.4 package.scala 96:25:@11497.4]
  assign _T_2873 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@11560.4 package.scala 96:25:@11561.4]
  assign _T_2877 = _T_2873 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11570.4]
  assign _T_2870 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@11552.4 package.scala 96:25:@11553.4]
  assign _T_2878 = _T_2870 ? Mem1D_7_io_output : _T_2877; // @[Mux.scala 31:69:@11571.4]
  assign _T_2867 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@11544.4 package.scala 96:25:@11545.4]
  assign _T_2908 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@11608.4 package.scala 96:25:@11609.4]
  assign _T_2912 = _T_2908 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11618.4]
  assign _T_2905 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@11600.4 package.scala 96:25:@11601.4]
  assign _T_2913 = _T_2905 ? Mem1D_7_io_output : _T_2912; // @[Mux.scala 31:69:@11619.4]
  assign _T_2902 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@11592.4 package.scala 96:25:@11593.4]
  assign _T_2943 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@11656.4 package.scala 96:25:@11657.4]
  assign _T_2947 = _T_2943 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@11666.4]
  assign _T_2940 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@11648.4 package.scala 96:25:@11649.4]
  assign _T_2948 = _T_2940 ? Mem1D_4_io_output : _T_2947; // @[Mux.scala 31:69:@11667.4]
  assign _T_2937 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@11640.4 package.scala 96:25:@11641.4]
  assign _T_2978 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@11704.4 package.scala 96:25:@11705.4]
  assign _T_2982 = _T_2978 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@11714.4]
  assign _T_2975 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@11696.4 package.scala 96:25:@11697.4]
  assign _T_2983 = _T_2975 ? Mem1D_5_io_output : _T_2982; // @[Mux.scala 31:69:@11715.4]
  assign _T_2972 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@11688.4 package.scala 96:25:@11689.4]
  assign _T_3013 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@11752.4 package.scala 96:25:@11753.4]
  assign _T_3017 = _T_3013 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11762.4]
  assign _T_3010 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@11744.4 package.scala 96:25:@11745.4]
  assign _T_3018 = _T_3010 ? Mem1D_6_io_output : _T_3017; // @[Mux.scala 31:69:@11763.4]
  assign _T_3007 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@11736.4 package.scala 96:25:@11737.4]
  assign _T_3048 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@11800.4 package.scala 96:25:@11801.4]
  assign _T_3052 = _T_3048 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11810.4]
  assign _T_3045 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@11792.4 package.scala 96:25:@11793.4]
  assign _T_3053 = _T_3045 ? Mem1D_6_io_output : _T_3052; // @[Mux.scala 31:69:@11811.4]
  assign _T_3042 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@11784.4 package.scala 96:25:@11785.4]
  assign io_rPort_23_output_0 = _T_3042 ? Mem1D_2_io_output : _T_3053; // @[MemPrimitives.scala 148:13:@11813.4]
  assign io_rPort_22_output_0 = _T_3007 ? Mem1D_2_io_output : _T_3018; // @[MemPrimitives.scala 148:13:@11765.4]
  assign io_rPort_21_output_0 = _T_2972 ? Mem1D_1_io_output : _T_2983; // @[MemPrimitives.scala 148:13:@11717.4]
  assign io_rPort_20_output_0 = _T_2937 ? Mem1D_io_output : _T_2948; // @[MemPrimitives.scala 148:13:@11669.4]
  assign io_rPort_19_output_0 = _T_2902 ? Mem1D_3_io_output : _T_2913; // @[MemPrimitives.scala 148:13:@11621.4]
  assign io_rPort_18_output_0 = _T_2867 ? Mem1D_3_io_output : _T_2878; // @[MemPrimitives.scala 148:13:@11573.4]
  assign io_rPort_17_output_0 = _T_2832 ? Mem1D_2_io_output : _T_2843; // @[MemPrimitives.scala 148:13:@11525.4]
  assign io_rPort_16_output_0 = _T_2797 ? Mem1D_3_io_output : _T_2808; // @[MemPrimitives.scala 148:13:@11477.4]
  assign io_rPort_15_output_0 = _T_2762 ? Mem1D_2_io_output : _T_2773; // @[MemPrimitives.scala 148:13:@11429.4]
  assign io_rPort_14_output_0 = _T_2727 ? Mem1D_3_io_output : _T_2738; // @[MemPrimitives.scala 148:13:@11381.4]
  assign io_rPort_13_output_0 = _T_2692 ? Mem1D_2_io_output : _T_2703; // @[MemPrimitives.scala 148:13:@11333.4]
  assign io_rPort_12_output_0 = _T_2657 ? Mem1D_3_io_output : _T_2668; // @[MemPrimitives.scala 148:13:@11285.4]
  assign io_rPort_11_output_0 = _T_2622 ? Mem1D_2_io_output : _T_2633; // @[MemPrimitives.scala 148:13:@11237.4]
  assign io_rPort_10_output_0 = _T_2587 ? Mem1D_io_output : _T_2598; // @[MemPrimitives.scala 148:13:@11189.4]
  assign io_rPort_9_output_0 = _T_2552 ? Mem1D_3_io_output : _T_2563; // @[MemPrimitives.scala 148:13:@11141.4]
  assign io_rPort_8_output_0 = _T_2517 ? Mem1D_3_io_output : _T_2528; // @[MemPrimitives.scala 148:13:@11093.4]
  assign io_rPort_7_output_0 = _T_2482 ? Mem1D_io_output : _T_2493; // @[MemPrimitives.scala 148:13:@11045.4]
  assign io_rPort_6_output_0 = _T_2447 ? Mem1D_1_io_output : _T_2458; // @[MemPrimitives.scala 148:13:@10997.4]
  assign io_rPort_5_output_0 = _T_2412 ? Mem1D_io_output : _T_2423; // @[MemPrimitives.scala 148:13:@10949.4]
  assign io_rPort_4_output_0 = _T_2377 ? Mem1D_2_io_output : _T_2388; // @[MemPrimitives.scala 148:13:@10901.4]
  assign io_rPort_3_output_0 = _T_2342 ? Mem1D_1_io_output : _T_2353; // @[MemPrimitives.scala 148:13:@10853.4]
  assign io_rPort_2_output_0 = _T_2307 ? Mem1D_2_io_output : _T_2318; // @[MemPrimitives.scala 148:13:@10805.4]
  assign io_rPort_1_output_0 = _T_2272 ? Mem1D_3_io_output : _T_2283; // @[MemPrimitives.scala 148:13:@10757.4]
  assign io_rPort_0_output_0 = _T_2237 ? Mem1D_1_io_output : _T_2248; // @[MemPrimitives.scala 148:13:@10709.4]
  assign Mem1D_clock = clock; // @[:@9239.4]
  assign Mem1D_reset = reset; // @[:@9240.4]
  assign Mem1D_io_r_ofs_0 = _T_1353[0]; // @[MemPrimitives.scala 127:28:@9803.4]
  assign Mem1D_io_r_backpressure = _T_1353[1]; // @[MemPrimitives.scala 128:32:@9804.4]
  assign Mem1D_io_w_ofs_0 = _T_1045[0]; // @[MemPrimitives.scala 94:28:@9508.4]
  assign Mem1D_io_w_data_0 = _T_1045[8:1]; // @[MemPrimitives.scala 95:29:@9509.4]
  assign Mem1D_io_w_en_0 = _T_1045[9]; // @[MemPrimitives.scala 96:27:@9510.4]
  assign Mem1D_1_clock = clock; // @[:@9255.4]
  assign Mem1D_1_reset = reset; // @[:@9256.4]
  assign Mem1D_1_io_r_ofs_0 = _T_1391[0]; // @[MemPrimitives.scala 127:28:@9843.4]
  assign Mem1D_1_io_r_backpressure = _T_1391[1]; // @[MemPrimitives.scala 128:32:@9844.4]
  assign Mem1D_1_io_w_ofs_0 = _T_1063[0]; // @[MemPrimitives.scala 94:28:@9525.4]
  assign Mem1D_1_io_w_data_0 = _T_1063[8:1]; // @[MemPrimitives.scala 95:29:@9526.4]
  assign Mem1D_1_io_w_en_0 = _T_1063[9]; // @[MemPrimitives.scala 96:27:@9527.4]
  assign Mem1D_2_clock = clock; // @[:@9271.4]
  assign Mem1D_2_reset = reset; // @[:@9272.4]
  assign Mem1D_2_io_r_ofs_0 = _T_1465[0]; // @[MemPrimitives.scala 127:28:@9915.4]
  assign Mem1D_2_io_r_backpressure = _T_1465[1]; // @[MemPrimitives.scala 128:32:@9916.4]
  assign Mem1D_2_io_w_ofs_0 = _T_1081[0]; // @[MemPrimitives.scala 94:28:@9542.4]
  assign Mem1D_2_io_w_data_0 = _T_1081[8:1]; // @[MemPrimitives.scala 95:29:@9543.4]
  assign Mem1D_2_io_w_en_0 = _T_1081[9]; // @[MemPrimitives.scala 96:27:@9544.4]
  assign Mem1D_3_clock = clock; // @[:@9287.4]
  assign Mem1D_3_reset = reset; // @[:@9288.4]
  assign Mem1D_3_io_r_ofs_0 = _T_1539[0]; // @[MemPrimitives.scala 127:28:@9987.4]
  assign Mem1D_3_io_r_backpressure = _T_1539[1]; // @[MemPrimitives.scala 128:32:@9988.4]
  assign Mem1D_3_io_w_ofs_0 = _T_1099[0]; // @[MemPrimitives.scala 94:28:@9559.4]
  assign Mem1D_3_io_w_data_0 = _T_1099[8:1]; // @[MemPrimitives.scala 95:29:@9560.4]
  assign Mem1D_3_io_w_en_0 = _T_1099[9]; // @[MemPrimitives.scala 96:27:@9561.4]
  assign Mem1D_4_clock = clock; // @[:@9303.4]
  assign Mem1D_4_reset = reset; // @[:@9304.4]
  assign Mem1D_4_io_r_ofs_0 = _T_1577[0]; // @[MemPrimitives.scala 127:28:@10027.4]
  assign Mem1D_4_io_r_backpressure = _T_1577[1]; // @[MemPrimitives.scala 128:32:@10028.4]
  assign Mem1D_4_io_w_ofs_0 = _T_1117[0]; // @[MemPrimitives.scala 94:28:@9576.4]
  assign Mem1D_4_io_w_data_0 = _T_1117[8:1]; // @[MemPrimitives.scala 95:29:@9577.4]
  assign Mem1D_4_io_w_en_0 = _T_1117[9]; // @[MemPrimitives.scala 96:27:@9578.4]
  assign Mem1D_5_clock = clock; // @[:@9319.4]
  assign Mem1D_5_reset = reset; // @[:@9320.4]
  assign Mem1D_5_io_r_ofs_0 = _T_1615[0]; // @[MemPrimitives.scala 127:28:@10067.4]
  assign Mem1D_5_io_r_backpressure = _T_1615[1]; // @[MemPrimitives.scala 128:32:@10068.4]
  assign Mem1D_5_io_w_ofs_0 = _T_1135[0]; // @[MemPrimitives.scala 94:28:@9593.4]
  assign Mem1D_5_io_w_data_0 = _T_1135[8:1]; // @[MemPrimitives.scala 95:29:@9594.4]
  assign Mem1D_5_io_w_en_0 = _T_1135[9]; // @[MemPrimitives.scala 96:27:@9595.4]
  assign Mem1D_6_clock = clock; // @[:@9335.4]
  assign Mem1D_6_reset = reset; // @[:@9336.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1689[0]; // @[MemPrimitives.scala 127:28:@10139.4]
  assign Mem1D_6_io_r_backpressure = _T_1689[1]; // @[MemPrimitives.scala 128:32:@10140.4]
  assign Mem1D_6_io_w_ofs_0 = _T_1153[0]; // @[MemPrimitives.scala 94:28:@9610.4]
  assign Mem1D_6_io_w_data_0 = _T_1153[8:1]; // @[MemPrimitives.scala 95:29:@9611.4]
  assign Mem1D_6_io_w_en_0 = _T_1153[9]; // @[MemPrimitives.scala 96:27:@9612.4]
  assign Mem1D_7_clock = clock; // @[:@9351.4]
  assign Mem1D_7_reset = reset; // @[:@9352.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1763[0]; // @[MemPrimitives.scala 127:28:@10211.4]
  assign Mem1D_7_io_r_backpressure = _T_1763[1]; // @[MemPrimitives.scala 128:32:@10212.4]
  assign Mem1D_7_io_w_ofs_0 = _T_1171[0]; // @[MemPrimitives.scala 94:28:@9627.4]
  assign Mem1D_7_io_w_data_0 = _T_1171[8:1]; // @[MemPrimitives.scala 95:29:@9628.4]
  assign Mem1D_7_io_w_en_0 = _T_1171[9]; // @[MemPrimitives.scala 96:27:@9629.4]
  assign Mem1D_8_clock = clock; // @[:@9367.4]
  assign Mem1D_8_reset = reset; // @[:@9368.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1801[0]; // @[MemPrimitives.scala 127:28:@10251.4]
  assign Mem1D_8_io_r_backpressure = _T_1801[1]; // @[MemPrimitives.scala 128:32:@10252.4]
  assign Mem1D_8_io_w_ofs_0 = _T_1189[0]; // @[MemPrimitives.scala 94:28:@9644.4]
  assign Mem1D_8_io_w_data_0 = _T_1189[8:1]; // @[MemPrimitives.scala 95:29:@9645.4]
  assign Mem1D_8_io_w_en_0 = _T_1189[9]; // @[MemPrimitives.scala 96:27:@9646.4]
  assign Mem1D_9_clock = clock; // @[:@9383.4]
  assign Mem1D_9_reset = reset; // @[:@9384.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1839[0]; // @[MemPrimitives.scala 127:28:@10291.4]
  assign Mem1D_9_io_r_backpressure = _T_1839[1]; // @[MemPrimitives.scala 128:32:@10292.4]
  assign Mem1D_9_io_w_ofs_0 = _T_1207[0]; // @[MemPrimitives.scala 94:28:@9661.4]
  assign Mem1D_9_io_w_data_0 = _T_1207[8:1]; // @[MemPrimitives.scala 95:29:@9662.4]
  assign Mem1D_9_io_w_en_0 = _T_1207[9]; // @[MemPrimitives.scala 96:27:@9663.4]
  assign Mem1D_10_clock = clock; // @[:@9399.4]
  assign Mem1D_10_reset = reset; // @[:@9400.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1913[0]; // @[MemPrimitives.scala 127:28:@10363.4]
  assign Mem1D_10_io_r_backpressure = _T_1913[1]; // @[MemPrimitives.scala 128:32:@10364.4]
  assign Mem1D_10_io_w_ofs_0 = _T_1225[0]; // @[MemPrimitives.scala 94:28:@9678.4]
  assign Mem1D_10_io_w_data_0 = _T_1225[8:1]; // @[MemPrimitives.scala 95:29:@9679.4]
  assign Mem1D_10_io_w_en_0 = _T_1225[9]; // @[MemPrimitives.scala 96:27:@9680.4]
  assign Mem1D_11_clock = clock; // @[:@9415.4]
  assign Mem1D_11_reset = reset; // @[:@9416.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1987[0]; // @[MemPrimitives.scala 127:28:@10435.4]
  assign Mem1D_11_io_r_backpressure = _T_1987[1]; // @[MemPrimitives.scala 128:32:@10436.4]
  assign Mem1D_11_io_w_ofs_0 = _T_1243[0]; // @[MemPrimitives.scala 94:28:@9695.4]
  assign Mem1D_11_io_w_data_0 = _T_1243[8:1]; // @[MemPrimitives.scala 95:29:@9696.4]
  assign Mem1D_11_io_w_en_0 = _T_1243[9]; // @[MemPrimitives.scala 96:27:@9697.4]
  assign Mem1D_12_clock = clock; // @[:@9431.4]
  assign Mem1D_12_reset = reset; // @[:@9432.4]
  assign Mem1D_12_io_r_ofs_0 = _T_2025[0]; // @[MemPrimitives.scala 127:28:@10475.4]
  assign Mem1D_12_io_r_backpressure = _T_2025[1]; // @[MemPrimitives.scala 128:32:@10476.4]
  assign Mem1D_12_io_w_ofs_0 = _T_1261[0]; // @[MemPrimitives.scala 94:28:@9712.4]
  assign Mem1D_12_io_w_data_0 = _T_1261[8:1]; // @[MemPrimitives.scala 95:29:@9713.4]
  assign Mem1D_12_io_w_en_0 = _T_1261[9]; // @[MemPrimitives.scala 96:27:@9714.4]
  assign Mem1D_13_clock = clock; // @[:@9447.4]
  assign Mem1D_13_reset = reset; // @[:@9448.4]
  assign Mem1D_13_io_r_ofs_0 = _T_2063[0]; // @[MemPrimitives.scala 127:28:@10515.4]
  assign Mem1D_13_io_r_backpressure = _T_2063[1]; // @[MemPrimitives.scala 128:32:@10516.4]
  assign Mem1D_13_io_w_ofs_0 = _T_1279[0]; // @[MemPrimitives.scala 94:28:@9729.4]
  assign Mem1D_13_io_w_data_0 = _T_1279[8:1]; // @[MemPrimitives.scala 95:29:@9730.4]
  assign Mem1D_13_io_w_en_0 = _T_1279[9]; // @[MemPrimitives.scala 96:27:@9731.4]
  assign Mem1D_14_clock = clock; // @[:@9463.4]
  assign Mem1D_14_reset = reset; // @[:@9464.4]
  assign Mem1D_14_io_r_ofs_0 = _T_2137[0]; // @[MemPrimitives.scala 127:28:@10587.4]
  assign Mem1D_14_io_r_backpressure = _T_2137[1]; // @[MemPrimitives.scala 128:32:@10588.4]
  assign Mem1D_14_io_w_ofs_0 = _T_1297[0]; // @[MemPrimitives.scala 94:28:@9746.4]
  assign Mem1D_14_io_w_data_0 = _T_1297[8:1]; // @[MemPrimitives.scala 95:29:@9747.4]
  assign Mem1D_14_io_w_en_0 = _T_1297[9]; // @[MemPrimitives.scala 96:27:@9748.4]
  assign Mem1D_15_clock = clock; // @[:@9479.4]
  assign Mem1D_15_reset = reset; // @[:@9480.4]
  assign Mem1D_15_io_r_ofs_0 = _T_2211[0]; // @[MemPrimitives.scala 127:28:@10659.4]
  assign Mem1D_15_io_r_backpressure = _T_2211[1]; // @[MemPrimitives.scala 128:32:@10660.4]
  assign Mem1D_15_io_w_ofs_0 = _T_1315[0]; // @[MemPrimitives.scala 94:28:@9763.4]
  assign Mem1D_15_io_w_data_0 = _T_1315[8:1]; // @[MemPrimitives.scala 95:29:@9764.4]
  assign Mem1D_15_io_w_en_0 = _T_1315[9]; // @[MemPrimitives.scala 96:27:@9765.4]
  assign StickySelects_clock = clock; // @[:@9779.4]
  assign StickySelects_reset = reset; // @[:@9780.4]
  assign StickySelects_io_ins_0 = io_rPort_5_en_0 & _T_1320; // @[MemPrimitives.scala 122:60:@9781.4]
  assign StickySelects_io_ins_1 = io_rPort_7_en_0 & _T_1325; // @[MemPrimitives.scala 122:60:@9782.4]
  assign StickySelects_io_ins_2 = io_rPort_10_en_0 & _T_1330; // @[MemPrimitives.scala 122:60:@9783.4]
  assign StickySelects_io_ins_3 = io_rPort_20_en_0 & _T_1335; // @[MemPrimitives.scala 122:60:@9784.4]
  assign StickySelects_1_clock = clock; // @[:@9819.4]
  assign StickySelects_1_reset = reset; // @[:@9820.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_1358; // @[MemPrimitives.scala 122:60:@9821.4]
  assign StickySelects_1_io_ins_1 = io_rPort_3_en_0 & _T_1363; // @[MemPrimitives.scala 122:60:@9822.4]
  assign StickySelects_1_io_ins_2 = io_rPort_6_en_0 & _T_1368; // @[MemPrimitives.scala 122:60:@9823.4]
  assign StickySelects_1_io_ins_3 = io_rPort_21_en_0 & _T_1373; // @[MemPrimitives.scala 122:60:@9824.4]
  assign StickySelects_2_clock = clock; // @[:@9871.4]
  assign StickySelects_2_reset = reset; // @[:@9872.4]
  assign StickySelects_2_io_ins_0 = io_rPort_2_en_0 & _T_1396; // @[MemPrimitives.scala 122:60:@9873.4]
  assign StickySelects_2_io_ins_1 = io_rPort_4_en_0 & _T_1401; // @[MemPrimitives.scala 122:60:@9874.4]
  assign StickySelects_2_io_ins_2 = io_rPort_11_en_0 & _T_1406; // @[MemPrimitives.scala 122:60:@9875.4]
  assign StickySelects_2_io_ins_3 = io_rPort_13_en_0 & _T_1411; // @[MemPrimitives.scala 122:60:@9876.4]
  assign StickySelects_2_io_ins_4 = io_rPort_15_en_0 & _T_1416; // @[MemPrimitives.scala 122:60:@9877.4]
  assign StickySelects_2_io_ins_5 = io_rPort_17_en_0 & _T_1421; // @[MemPrimitives.scala 122:60:@9878.4]
  assign StickySelects_2_io_ins_6 = io_rPort_22_en_0 & _T_1426; // @[MemPrimitives.scala 122:60:@9879.4]
  assign StickySelects_2_io_ins_7 = io_rPort_23_en_0 & _T_1431; // @[MemPrimitives.scala 122:60:@9880.4]
  assign StickySelects_3_clock = clock; // @[:@9943.4]
  assign StickySelects_3_reset = reset; // @[:@9944.4]
  assign StickySelects_3_io_ins_0 = io_rPort_1_en_0 & _T_1470; // @[MemPrimitives.scala 122:60:@9945.4]
  assign StickySelects_3_io_ins_1 = io_rPort_8_en_0 & _T_1475; // @[MemPrimitives.scala 122:60:@9946.4]
  assign StickySelects_3_io_ins_2 = io_rPort_9_en_0 & _T_1480; // @[MemPrimitives.scala 122:60:@9947.4]
  assign StickySelects_3_io_ins_3 = io_rPort_12_en_0 & _T_1485; // @[MemPrimitives.scala 122:60:@9948.4]
  assign StickySelects_3_io_ins_4 = io_rPort_14_en_0 & _T_1490; // @[MemPrimitives.scala 122:60:@9949.4]
  assign StickySelects_3_io_ins_5 = io_rPort_16_en_0 & _T_1495; // @[MemPrimitives.scala 122:60:@9950.4]
  assign StickySelects_3_io_ins_6 = io_rPort_18_en_0 & _T_1500; // @[MemPrimitives.scala 122:60:@9951.4]
  assign StickySelects_3_io_ins_7 = io_rPort_19_en_0 & _T_1505; // @[MemPrimitives.scala 122:60:@9952.4]
  assign StickySelects_4_clock = clock; // @[:@10003.4]
  assign StickySelects_4_reset = reset; // @[:@10004.4]
  assign StickySelects_4_io_ins_0 = io_rPort_5_en_0 & _T_1544; // @[MemPrimitives.scala 122:60:@10005.4]
  assign StickySelects_4_io_ins_1 = io_rPort_7_en_0 & _T_1549; // @[MemPrimitives.scala 122:60:@10006.4]
  assign StickySelects_4_io_ins_2 = io_rPort_10_en_0 & _T_1554; // @[MemPrimitives.scala 122:60:@10007.4]
  assign StickySelects_4_io_ins_3 = io_rPort_20_en_0 & _T_1559; // @[MemPrimitives.scala 122:60:@10008.4]
  assign StickySelects_5_clock = clock; // @[:@10043.4]
  assign StickySelects_5_reset = reset; // @[:@10044.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_1582; // @[MemPrimitives.scala 122:60:@10045.4]
  assign StickySelects_5_io_ins_1 = io_rPort_3_en_0 & _T_1587; // @[MemPrimitives.scala 122:60:@10046.4]
  assign StickySelects_5_io_ins_2 = io_rPort_6_en_0 & _T_1592; // @[MemPrimitives.scala 122:60:@10047.4]
  assign StickySelects_5_io_ins_3 = io_rPort_21_en_0 & _T_1597; // @[MemPrimitives.scala 122:60:@10048.4]
  assign StickySelects_6_clock = clock; // @[:@10095.4]
  assign StickySelects_6_reset = reset; // @[:@10096.4]
  assign StickySelects_6_io_ins_0 = io_rPort_2_en_0 & _T_1620; // @[MemPrimitives.scala 122:60:@10097.4]
  assign StickySelects_6_io_ins_1 = io_rPort_4_en_0 & _T_1625; // @[MemPrimitives.scala 122:60:@10098.4]
  assign StickySelects_6_io_ins_2 = io_rPort_11_en_0 & _T_1630; // @[MemPrimitives.scala 122:60:@10099.4]
  assign StickySelects_6_io_ins_3 = io_rPort_13_en_0 & _T_1635; // @[MemPrimitives.scala 122:60:@10100.4]
  assign StickySelects_6_io_ins_4 = io_rPort_15_en_0 & _T_1640; // @[MemPrimitives.scala 122:60:@10101.4]
  assign StickySelects_6_io_ins_5 = io_rPort_17_en_0 & _T_1645; // @[MemPrimitives.scala 122:60:@10102.4]
  assign StickySelects_6_io_ins_6 = io_rPort_22_en_0 & _T_1650; // @[MemPrimitives.scala 122:60:@10103.4]
  assign StickySelects_6_io_ins_7 = io_rPort_23_en_0 & _T_1655; // @[MemPrimitives.scala 122:60:@10104.4]
  assign StickySelects_7_clock = clock; // @[:@10167.4]
  assign StickySelects_7_reset = reset; // @[:@10168.4]
  assign StickySelects_7_io_ins_0 = io_rPort_1_en_0 & _T_1694; // @[MemPrimitives.scala 122:60:@10169.4]
  assign StickySelects_7_io_ins_1 = io_rPort_8_en_0 & _T_1699; // @[MemPrimitives.scala 122:60:@10170.4]
  assign StickySelects_7_io_ins_2 = io_rPort_9_en_0 & _T_1704; // @[MemPrimitives.scala 122:60:@10171.4]
  assign StickySelects_7_io_ins_3 = io_rPort_12_en_0 & _T_1709; // @[MemPrimitives.scala 122:60:@10172.4]
  assign StickySelects_7_io_ins_4 = io_rPort_14_en_0 & _T_1714; // @[MemPrimitives.scala 122:60:@10173.4]
  assign StickySelects_7_io_ins_5 = io_rPort_16_en_0 & _T_1719; // @[MemPrimitives.scala 122:60:@10174.4]
  assign StickySelects_7_io_ins_6 = io_rPort_18_en_0 & _T_1724; // @[MemPrimitives.scala 122:60:@10175.4]
  assign StickySelects_7_io_ins_7 = io_rPort_19_en_0 & _T_1729; // @[MemPrimitives.scala 122:60:@10176.4]
  assign StickySelects_8_clock = clock; // @[:@10227.4]
  assign StickySelects_8_reset = reset; // @[:@10228.4]
  assign StickySelects_8_io_ins_0 = io_rPort_5_en_0 & _T_1768; // @[MemPrimitives.scala 122:60:@10229.4]
  assign StickySelects_8_io_ins_1 = io_rPort_7_en_0 & _T_1773; // @[MemPrimitives.scala 122:60:@10230.4]
  assign StickySelects_8_io_ins_2 = io_rPort_10_en_0 & _T_1778; // @[MemPrimitives.scala 122:60:@10231.4]
  assign StickySelects_8_io_ins_3 = io_rPort_20_en_0 & _T_1783; // @[MemPrimitives.scala 122:60:@10232.4]
  assign StickySelects_9_clock = clock; // @[:@10267.4]
  assign StickySelects_9_reset = reset; // @[:@10268.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_1806; // @[MemPrimitives.scala 122:60:@10269.4]
  assign StickySelects_9_io_ins_1 = io_rPort_3_en_0 & _T_1811; // @[MemPrimitives.scala 122:60:@10270.4]
  assign StickySelects_9_io_ins_2 = io_rPort_6_en_0 & _T_1816; // @[MemPrimitives.scala 122:60:@10271.4]
  assign StickySelects_9_io_ins_3 = io_rPort_21_en_0 & _T_1821; // @[MemPrimitives.scala 122:60:@10272.4]
  assign StickySelects_10_clock = clock; // @[:@10319.4]
  assign StickySelects_10_reset = reset; // @[:@10320.4]
  assign StickySelects_10_io_ins_0 = io_rPort_2_en_0 & _T_1844; // @[MemPrimitives.scala 122:60:@10321.4]
  assign StickySelects_10_io_ins_1 = io_rPort_4_en_0 & _T_1849; // @[MemPrimitives.scala 122:60:@10322.4]
  assign StickySelects_10_io_ins_2 = io_rPort_11_en_0 & _T_1854; // @[MemPrimitives.scala 122:60:@10323.4]
  assign StickySelects_10_io_ins_3 = io_rPort_13_en_0 & _T_1859; // @[MemPrimitives.scala 122:60:@10324.4]
  assign StickySelects_10_io_ins_4 = io_rPort_15_en_0 & _T_1864; // @[MemPrimitives.scala 122:60:@10325.4]
  assign StickySelects_10_io_ins_5 = io_rPort_17_en_0 & _T_1869; // @[MemPrimitives.scala 122:60:@10326.4]
  assign StickySelects_10_io_ins_6 = io_rPort_22_en_0 & _T_1874; // @[MemPrimitives.scala 122:60:@10327.4]
  assign StickySelects_10_io_ins_7 = io_rPort_23_en_0 & _T_1879; // @[MemPrimitives.scala 122:60:@10328.4]
  assign StickySelects_11_clock = clock; // @[:@10391.4]
  assign StickySelects_11_reset = reset; // @[:@10392.4]
  assign StickySelects_11_io_ins_0 = io_rPort_1_en_0 & _T_1918; // @[MemPrimitives.scala 122:60:@10393.4]
  assign StickySelects_11_io_ins_1 = io_rPort_8_en_0 & _T_1923; // @[MemPrimitives.scala 122:60:@10394.4]
  assign StickySelects_11_io_ins_2 = io_rPort_9_en_0 & _T_1928; // @[MemPrimitives.scala 122:60:@10395.4]
  assign StickySelects_11_io_ins_3 = io_rPort_12_en_0 & _T_1933; // @[MemPrimitives.scala 122:60:@10396.4]
  assign StickySelects_11_io_ins_4 = io_rPort_14_en_0 & _T_1938; // @[MemPrimitives.scala 122:60:@10397.4]
  assign StickySelects_11_io_ins_5 = io_rPort_16_en_0 & _T_1943; // @[MemPrimitives.scala 122:60:@10398.4]
  assign StickySelects_11_io_ins_6 = io_rPort_18_en_0 & _T_1948; // @[MemPrimitives.scala 122:60:@10399.4]
  assign StickySelects_11_io_ins_7 = io_rPort_19_en_0 & _T_1953; // @[MemPrimitives.scala 122:60:@10400.4]
  assign StickySelects_12_clock = clock; // @[:@10451.4]
  assign StickySelects_12_reset = reset; // @[:@10452.4]
  assign StickySelects_12_io_ins_0 = io_rPort_5_en_0 & _T_1992; // @[MemPrimitives.scala 122:60:@10453.4]
  assign StickySelects_12_io_ins_1 = io_rPort_7_en_0 & _T_1997; // @[MemPrimitives.scala 122:60:@10454.4]
  assign StickySelects_12_io_ins_2 = io_rPort_10_en_0 & _T_2002; // @[MemPrimitives.scala 122:60:@10455.4]
  assign StickySelects_12_io_ins_3 = io_rPort_20_en_0 & _T_2007; // @[MemPrimitives.scala 122:60:@10456.4]
  assign StickySelects_13_clock = clock; // @[:@10491.4]
  assign StickySelects_13_reset = reset; // @[:@10492.4]
  assign StickySelects_13_io_ins_0 = io_rPort_0_en_0 & _T_2030; // @[MemPrimitives.scala 122:60:@10493.4]
  assign StickySelects_13_io_ins_1 = io_rPort_3_en_0 & _T_2035; // @[MemPrimitives.scala 122:60:@10494.4]
  assign StickySelects_13_io_ins_2 = io_rPort_6_en_0 & _T_2040; // @[MemPrimitives.scala 122:60:@10495.4]
  assign StickySelects_13_io_ins_3 = io_rPort_21_en_0 & _T_2045; // @[MemPrimitives.scala 122:60:@10496.4]
  assign StickySelects_14_clock = clock; // @[:@10543.4]
  assign StickySelects_14_reset = reset; // @[:@10544.4]
  assign StickySelects_14_io_ins_0 = io_rPort_2_en_0 & _T_2068; // @[MemPrimitives.scala 122:60:@10545.4]
  assign StickySelects_14_io_ins_1 = io_rPort_4_en_0 & _T_2073; // @[MemPrimitives.scala 122:60:@10546.4]
  assign StickySelects_14_io_ins_2 = io_rPort_11_en_0 & _T_2078; // @[MemPrimitives.scala 122:60:@10547.4]
  assign StickySelects_14_io_ins_3 = io_rPort_13_en_0 & _T_2083; // @[MemPrimitives.scala 122:60:@10548.4]
  assign StickySelects_14_io_ins_4 = io_rPort_15_en_0 & _T_2088; // @[MemPrimitives.scala 122:60:@10549.4]
  assign StickySelects_14_io_ins_5 = io_rPort_17_en_0 & _T_2093; // @[MemPrimitives.scala 122:60:@10550.4]
  assign StickySelects_14_io_ins_6 = io_rPort_22_en_0 & _T_2098; // @[MemPrimitives.scala 122:60:@10551.4]
  assign StickySelects_14_io_ins_7 = io_rPort_23_en_0 & _T_2103; // @[MemPrimitives.scala 122:60:@10552.4]
  assign StickySelects_15_clock = clock; // @[:@10615.4]
  assign StickySelects_15_reset = reset; // @[:@10616.4]
  assign StickySelects_15_io_ins_0 = io_rPort_1_en_0 & _T_2142; // @[MemPrimitives.scala 122:60:@10617.4]
  assign StickySelects_15_io_ins_1 = io_rPort_8_en_0 & _T_2147; // @[MemPrimitives.scala 122:60:@10618.4]
  assign StickySelects_15_io_ins_2 = io_rPort_9_en_0 & _T_2152; // @[MemPrimitives.scala 122:60:@10619.4]
  assign StickySelects_15_io_ins_3 = io_rPort_12_en_0 & _T_2157; // @[MemPrimitives.scala 122:60:@10620.4]
  assign StickySelects_15_io_ins_4 = io_rPort_14_en_0 & _T_2162; // @[MemPrimitives.scala 122:60:@10621.4]
  assign StickySelects_15_io_ins_5 = io_rPort_16_en_0 & _T_2167; // @[MemPrimitives.scala 122:60:@10622.4]
  assign StickySelects_15_io_ins_6 = io_rPort_18_en_0 & _T_2172; // @[MemPrimitives.scala 122:60:@10623.4]
  assign StickySelects_15_io_ins_7 = io_rPort_19_en_0 & _T_2177; // @[MemPrimitives.scala 122:60:@10624.4]
  assign RetimeWrapper_clock = clock; // @[:@10676.4]
  assign RetimeWrapper_reset = reset; // @[:@10677.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10679.4]
  assign RetimeWrapper_io_in = _T_1358 & io_rPort_0_en_0; // @[package.scala 94:16:@10678.4]
  assign RetimeWrapper_1_clock = clock; // @[:@10684.4]
  assign RetimeWrapper_1_reset = reset; // @[:@10685.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10687.4]
  assign RetimeWrapper_1_io_in = _T_1582 & io_rPort_0_en_0; // @[package.scala 94:16:@10686.4]
  assign RetimeWrapper_2_clock = clock; // @[:@10692.4]
  assign RetimeWrapper_2_reset = reset; // @[:@10693.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10695.4]
  assign RetimeWrapper_2_io_in = _T_1806 & io_rPort_0_en_0; // @[package.scala 94:16:@10694.4]
  assign RetimeWrapper_3_clock = clock; // @[:@10700.4]
  assign RetimeWrapper_3_reset = reset; // @[:@10701.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10703.4]
  assign RetimeWrapper_3_io_in = _T_2030 & io_rPort_0_en_0; // @[package.scala 94:16:@10702.4]
  assign RetimeWrapper_4_clock = clock; // @[:@10724.4]
  assign RetimeWrapper_4_reset = reset; // @[:@10725.4]
  assign RetimeWrapper_4_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10727.4]
  assign RetimeWrapper_4_io_in = _T_1470 & io_rPort_1_en_0; // @[package.scala 94:16:@10726.4]
  assign RetimeWrapper_5_clock = clock; // @[:@10732.4]
  assign RetimeWrapper_5_reset = reset; // @[:@10733.4]
  assign RetimeWrapper_5_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10735.4]
  assign RetimeWrapper_5_io_in = _T_1694 & io_rPort_1_en_0; // @[package.scala 94:16:@10734.4]
  assign RetimeWrapper_6_clock = clock; // @[:@10740.4]
  assign RetimeWrapper_6_reset = reset; // @[:@10741.4]
  assign RetimeWrapper_6_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10743.4]
  assign RetimeWrapper_6_io_in = _T_1918 & io_rPort_1_en_0; // @[package.scala 94:16:@10742.4]
  assign RetimeWrapper_7_clock = clock; // @[:@10748.4]
  assign RetimeWrapper_7_reset = reset; // @[:@10749.4]
  assign RetimeWrapper_7_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10751.4]
  assign RetimeWrapper_7_io_in = _T_2142 & io_rPort_1_en_0; // @[package.scala 94:16:@10750.4]
  assign RetimeWrapper_8_clock = clock; // @[:@10772.4]
  assign RetimeWrapper_8_reset = reset; // @[:@10773.4]
  assign RetimeWrapper_8_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10775.4]
  assign RetimeWrapper_8_io_in = _T_1396 & io_rPort_2_en_0; // @[package.scala 94:16:@10774.4]
  assign RetimeWrapper_9_clock = clock; // @[:@10780.4]
  assign RetimeWrapper_9_reset = reset; // @[:@10781.4]
  assign RetimeWrapper_9_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10783.4]
  assign RetimeWrapper_9_io_in = _T_1620 & io_rPort_2_en_0; // @[package.scala 94:16:@10782.4]
  assign RetimeWrapper_10_clock = clock; // @[:@10788.4]
  assign RetimeWrapper_10_reset = reset; // @[:@10789.4]
  assign RetimeWrapper_10_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10791.4]
  assign RetimeWrapper_10_io_in = _T_1844 & io_rPort_2_en_0; // @[package.scala 94:16:@10790.4]
  assign RetimeWrapper_11_clock = clock; // @[:@10796.4]
  assign RetimeWrapper_11_reset = reset; // @[:@10797.4]
  assign RetimeWrapper_11_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10799.4]
  assign RetimeWrapper_11_io_in = _T_2068 & io_rPort_2_en_0; // @[package.scala 94:16:@10798.4]
  assign RetimeWrapper_12_clock = clock; // @[:@10820.4]
  assign RetimeWrapper_12_reset = reset; // @[:@10821.4]
  assign RetimeWrapper_12_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10823.4]
  assign RetimeWrapper_12_io_in = _T_1363 & io_rPort_3_en_0; // @[package.scala 94:16:@10822.4]
  assign RetimeWrapper_13_clock = clock; // @[:@10828.4]
  assign RetimeWrapper_13_reset = reset; // @[:@10829.4]
  assign RetimeWrapper_13_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10831.4]
  assign RetimeWrapper_13_io_in = _T_1587 & io_rPort_3_en_0; // @[package.scala 94:16:@10830.4]
  assign RetimeWrapper_14_clock = clock; // @[:@10836.4]
  assign RetimeWrapper_14_reset = reset; // @[:@10837.4]
  assign RetimeWrapper_14_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10839.4]
  assign RetimeWrapper_14_io_in = _T_1811 & io_rPort_3_en_0; // @[package.scala 94:16:@10838.4]
  assign RetimeWrapper_15_clock = clock; // @[:@10844.4]
  assign RetimeWrapper_15_reset = reset; // @[:@10845.4]
  assign RetimeWrapper_15_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10847.4]
  assign RetimeWrapper_15_io_in = _T_2035 & io_rPort_3_en_0; // @[package.scala 94:16:@10846.4]
  assign RetimeWrapper_16_clock = clock; // @[:@10868.4]
  assign RetimeWrapper_16_reset = reset; // @[:@10869.4]
  assign RetimeWrapper_16_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10871.4]
  assign RetimeWrapper_16_io_in = _T_1401 & io_rPort_4_en_0; // @[package.scala 94:16:@10870.4]
  assign RetimeWrapper_17_clock = clock; // @[:@10876.4]
  assign RetimeWrapper_17_reset = reset; // @[:@10877.4]
  assign RetimeWrapper_17_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10879.4]
  assign RetimeWrapper_17_io_in = _T_1625 & io_rPort_4_en_0; // @[package.scala 94:16:@10878.4]
  assign RetimeWrapper_18_clock = clock; // @[:@10884.4]
  assign RetimeWrapper_18_reset = reset; // @[:@10885.4]
  assign RetimeWrapper_18_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10887.4]
  assign RetimeWrapper_18_io_in = _T_1849 & io_rPort_4_en_0; // @[package.scala 94:16:@10886.4]
  assign RetimeWrapper_19_clock = clock; // @[:@10892.4]
  assign RetimeWrapper_19_reset = reset; // @[:@10893.4]
  assign RetimeWrapper_19_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10895.4]
  assign RetimeWrapper_19_io_in = _T_2073 & io_rPort_4_en_0; // @[package.scala 94:16:@10894.4]
  assign RetimeWrapper_20_clock = clock; // @[:@10916.4]
  assign RetimeWrapper_20_reset = reset; // @[:@10917.4]
  assign RetimeWrapper_20_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@10919.4]
  assign RetimeWrapper_20_io_in = _T_1320 & io_rPort_5_en_0; // @[package.scala 94:16:@10918.4]
  assign RetimeWrapper_21_clock = clock; // @[:@10924.4]
  assign RetimeWrapper_21_reset = reset; // @[:@10925.4]
  assign RetimeWrapper_21_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@10927.4]
  assign RetimeWrapper_21_io_in = _T_1544 & io_rPort_5_en_0; // @[package.scala 94:16:@10926.4]
  assign RetimeWrapper_22_clock = clock; // @[:@10932.4]
  assign RetimeWrapper_22_reset = reset; // @[:@10933.4]
  assign RetimeWrapper_22_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@10935.4]
  assign RetimeWrapper_22_io_in = _T_1768 & io_rPort_5_en_0; // @[package.scala 94:16:@10934.4]
  assign RetimeWrapper_23_clock = clock; // @[:@10940.4]
  assign RetimeWrapper_23_reset = reset; // @[:@10941.4]
  assign RetimeWrapper_23_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@10943.4]
  assign RetimeWrapper_23_io_in = _T_1992 & io_rPort_5_en_0; // @[package.scala 94:16:@10942.4]
  assign RetimeWrapper_24_clock = clock; // @[:@10964.4]
  assign RetimeWrapper_24_reset = reset; // @[:@10965.4]
  assign RetimeWrapper_24_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@10967.4]
  assign RetimeWrapper_24_io_in = _T_1368 & io_rPort_6_en_0; // @[package.scala 94:16:@10966.4]
  assign RetimeWrapper_25_clock = clock; // @[:@10972.4]
  assign RetimeWrapper_25_reset = reset; // @[:@10973.4]
  assign RetimeWrapper_25_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@10975.4]
  assign RetimeWrapper_25_io_in = _T_1592 & io_rPort_6_en_0; // @[package.scala 94:16:@10974.4]
  assign RetimeWrapper_26_clock = clock; // @[:@10980.4]
  assign RetimeWrapper_26_reset = reset; // @[:@10981.4]
  assign RetimeWrapper_26_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@10983.4]
  assign RetimeWrapper_26_io_in = _T_1816 & io_rPort_6_en_0; // @[package.scala 94:16:@10982.4]
  assign RetimeWrapper_27_clock = clock; // @[:@10988.4]
  assign RetimeWrapper_27_reset = reset; // @[:@10989.4]
  assign RetimeWrapper_27_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@10991.4]
  assign RetimeWrapper_27_io_in = _T_2040 & io_rPort_6_en_0; // @[package.scala 94:16:@10990.4]
  assign RetimeWrapper_28_clock = clock; // @[:@11012.4]
  assign RetimeWrapper_28_reset = reset; // @[:@11013.4]
  assign RetimeWrapper_28_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11015.4]
  assign RetimeWrapper_28_io_in = _T_1325 & io_rPort_7_en_0; // @[package.scala 94:16:@11014.4]
  assign RetimeWrapper_29_clock = clock; // @[:@11020.4]
  assign RetimeWrapper_29_reset = reset; // @[:@11021.4]
  assign RetimeWrapper_29_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11023.4]
  assign RetimeWrapper_29_io_in = _T_1549 & io_rPort_7_en_0; // @[package.scala 94:16:@11022.4]
  assign RetimeWrapper_30_clock = clock; // @[:@11028.4]
  assign RetimeWrapper_30_reset = reset; // @[:@11029.4]
  assign RetimeWrapper_30_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11031.4]
  assign RetimeWrapper_30_io_in = _T_1773 & io_rPort_7_en_0; // @[package.scala 94:16:@11030.4]
  assign RetimeWrapper_31_clock = clock; // @[:@11036.4]
  assign RetimeWrapper_31_reset = reset; // @[:@11037.4]
  assign RetimeWrapper_31_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11039.4]
  assign RetimeWrapper_31_io_in = _T_1997 & io_rPort_7_en_0; // @[package.scala 94:16:@11038.4]
  assign RetimeWrapper_32_clock = clock; // @[:@11060.4]
  assign RetimeWrapper_32_reset = reset; // @[:@11061.4]
  assign RetimeWrapper_32_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11063.4]
  assign RetimeWrapper_32_io_in = _T_1475 & io_rPort_8_en_0; // @[package.scala 94:16:@11062.4]
  assign RetimeWrapper_33_clock = clock; // @[:@11068.4]
  assign RetimeWrapper_33_reset = reset; // @[:@11069.4]
  assign RetimeWrapper_33_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11071.4]
  assign RetimeWrapper_33_io_in = _T_1699 & io_rPort_8_en_0; // @[package.scala 94:16:@11070.4]
  assign RetimeWrapper_34_clock = clock; // @[:@11076.4]
  assign RetimeWrapper_34_reset = reset; // @[:@11077.4]
  assign RetimeWrapper_34_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11079.4]
  assign RetimeWrapper_34_io_in = _T_1923 & io_rPort_8_en_0; // @[package.scala 94:16:@11078.4]
  assign RetimeWrapper_35_clock = clock; // @[:@11084.4]
  assign RetimeWrapper_35_reset = reset; // @[:@11085.4]
  assign RetimeWrapper_35_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11087.4]
  assign RetimeWrapper_35_io_in = _T_2147 & io_rPort_8_en_0; // @[package.scala 94:16:@11086.4]
  assign RetimeWrapper_36_clock = clock; // @[:@11108.4]
  assign RetimeWrapper_36_reset = reset; // @[:@11109.4]
  assign RetimeWrapper_36_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11111.4]
  assign RetimeWrapper_36_io_in = _T_1480 & io_rPort_9_en_0; // @[package.scala 94:16:@11110.4]
  assign RetimeWrapper_37_clock = clock; // @[:@11116.4]
  assign RetimeWrapper_37_reset = reset; // @[:@11117.4]
  assign RetimeWrapper_37_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11119.4]
  assign RetimeWrapper_37_io_in = _T_1704 & io_rPort_9_en_0; // @[package.scala 94:16:@11118.4]
  assign RetimeWrapper_38_clock = clock; // @[:@11124.4]
  assign RetimeWrapper_38_reset = reset; // @[:@11125.4]
  assign RetimeWrapper_38_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11127.4]
  assign RetimeWrapper_38_io_in = _T_1928 & io_rPort_9_en_0; // @[package.scala 94:16:@11126.4]
  assign RetimeWrapper_39_clock = clock; // @[:@11132.4]
  assign RetimeWrapper_39_reset = reset; // @[:@11133.4]
  assign RetimeWrapper_39_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11135.4]
  assign RetimeWrapper_39_io_in = _T_2152 & io_rPort_9_en_0; // @[package.scala 94:16:@11134.4]
  assign RetimeWrapper_40_clock = clock; // @[:@11156.4]
  assign RetimeWrapper_40_reset = reset; // @[:@11157.4]
  assign RetimeWrapper_40_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11159.4]
  assign RetimeWrapper_40_io_in = _T_1330 & io_rPort_10_en_0; // @[package.scala 94:16:@11158.4]
  assign RetimeWrapper_41_clock = clock; // @[:@11164.4]
  assign RetimeWrapper_41_reset = reset; // @[:@11165.4]
  assign RetimeWrapper_41_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11167.4]
  assign RetimeWrapper_41_io_in = _T_1554 & io_rPort_10_en_0; // @[package.scala 94:16:@11166.4]
  assign RetimeWrapper_42_clock = clock; // @[:@11172.4]
  assign RetimeWrapper_42_reset = reset; // @[:@11173.4]
  assign RetimeWrapper_42_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11175.4]
  assign RetimeWrapper_42_io_in = _T_1778 & io_rPort_10_en_0; // @[package.scala 94:16:@11174.4]
  assign RetimeWrapper_43_clock = clock; // @[:@11180.4]
  assign RetimeWrapper_43_reset = reset; // @[:@11181.4]
  assign RetimeWrapper_43_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11183.4]
  assign RetimeWrapper_43_io_in = _T_2002 & io_rPort_10_en_0; // @[package.scala 94:16:@11182.4]
  assign RetimeWrapper_44_clock = clock; // @[:@11204.4]
  assign RetimeWrapper_44_reset = reset; // @[:@11205.4]
  assign RetimeWrapper_44_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11207.4]
  assign RetimeWrapper_44_io_in = _T_1406 & io_rPort_11_en_0; // @[package.scala 94:16:@11206.4]
  assign RetimeWrapper_45_clock = clock; // @[:@11212.4]
  assign RetimeWrapper_45_reset = reset; // @[:@11213.4]
  assign RetimeWrapper_45_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11215.4]
  assign RetimeWrapper_45_io_in = _T_1630 & io_rPort_11_en_0; // @[package.scala 94:16:@11214.4]
  assign RetimeWrapper_46_clock = clock; // @[:@11220.4]
  assign RetimeWrapper_46_reset = reset; // @[:@11221.4]
  assign RetimeWrapper_46_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11223.4]
  assign RetimeWrapper_46_io_in = _T_1854 & io_rPort_11_en_0; // @[package.scala 94:16:@11222.4]
  assign RetimeWrapper_47_clock = clock; // @[:@11228.4]
  assign RetimeWrapper_47_reset = reset; // @[:@11229.4]
  assign RetimeWrapper_47_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11231.4]
  assign RetimeWrapper_47_io_in = _T_2078 & io_rPort_11_en_0; // @[package.scala 94:16:@11230.4]
  assign RetimeWrapper_48_clock = clock; // @[:@11252.4]
  assign RetimeWrapper_48_reset = reset; // @[:@11253.4]
  assign RetimeWrapper_48_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@11255.4]
  assign RetimeWrapper_48_io_in = _T_1485 & io_rPort_12_en_0; // @[package.scala 94:16:@11254.4]
  assign RetimeWrapper_49_clock = clock; // @[:@11260.4]
  assign RetimeWrapper_49_reset = reset; // @[:@11261.4]
  assign RetimeWrapper_49_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@11263.4]
  assign RetimeWrapper_49_io_in = _T_1709 & io_rPort_12_en_0; // @[package.scala 94:16:@11262.4]
  assign RetimeWrapper_50_clock = clock; // @[:@11268.4]
  assign RetimeWrapper_50_reset = reset; // @[:@11269.4]
  assign RetimeWrapper_50_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@11271.4]
  assign RetimeWrapper_50_io_in = _T_1933 & io_rPort_12_en_0; // @[package.scala 94:16:@11270.4]
  assign RetimeWrapper_51_clock = clock; // @[:@11276.4]
  assign RetimeWrapper_51_reset = reset; // @[:@11277.4]
  assign RetimeWrapper_51_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@11279.4]
  assign RetimeWrapper_51_io_in = _T_2157 & io_rPort_12_en_0; // @[package.scala 94:16:@11278.4]
  assign RetimeWrapper_52_clock = clock; // @[:@11300.4]
  assign RetimeWrapper_52_reset = reset; // @[:@11301.4]
  assign RetimeWrapper_52_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@11303.4]
  assign RetimeWrapper_52_io_in = _T_1411 & io_rPort_13_en_0; // @[package.scala 94:16:@11302.4]
  assign RetimeWrapper_53_clock = clock; // @[:@11308.4]
  assign RetimeWrapper_53_reset = reset; // @[:@11309.4]
  assign RetimeWrapper_53_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@11311.4]
  assign RetimeWrapper_53_io_in = _T_1635 & io_rPort_13_en_0; // @[package.scala 94:16:@11310.4]
  assign RetimeWrapper_54_clock = clock; // @[:@11316.4]
  assign RetimeWrapper_54_reset = reset; // @[:@11317.4]
  assign RetimeWrapper_54_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@11319.4]
  assign RetimeWrapper_54_io_in = _T_1859 & io_rPort_13_en_0; // @[package.scala 94:16:@11318.4]
  assign RetimeWrapper_55_clock = clock; // @[:@11324.4]
  assign RetimeWrapper_55_reset = reset; // @[:@11325.4]
  assign RetimeWrapper_55_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@11327.4]
  assign RetimeWrapper_55_io_in = _T_2083 & io_rPort_13_en_0; // @[package.scala 94:16:@11326.4]
  assign RetimeWrapper_56_clock = clock; // @[:@11348.4]
  assign RetimeWrapper_56_reset = reset; // @[:@11349.4]
  assign RetimeWrapper_56_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@11351.4]
  assign RetimeWrapper_56_io_in = _T_1490 & io_rPort_14_en_0; // @[package.scala 94:16:@11350.4]
  assign RetimeWrapper_57_clock = clock; // @[:@11356.4]
  assign RetimeWrapper_57_reset = reset; // @[:@11357.4]
  assign RetimeWrapper_57_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@11359.4]
  assign RetimeWrapper_57_io_in = _T_1714 & io_rPort_14_en_0; // @[package.scala 94:16:@11358.4]
  assign RetimeWrapper_58_clock = clock; // @[:@11364.4]
  assign RetimeWrapper_58_reset = reset; // @[:@11365.4]
  assign RetimeWrapper_58_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@11367.4]
  assign RetimeWrapper_58_io_in = _T_1938 & io_rPort_14_en_0; // @[package.scala 94:16:@11366.4]
  assign RetimeWrapper_59_clock = clock; // @[:@11372.4]
  assign RetimeWrapper_59_reset = reset; // @[:@11373.4]
  assign RetimeWrapper_59_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@11375.4]
  assign RetimeWrapper_59_io_in = _T_2162 & io_rPort_14_en_0; // @[package.scala 94:16:@11374.4]
  assign RetimeWrapper_60_clock = clock; // @[:@11396.4]
  assign RetimeWrapper_60_reset = reset; // @[:@11397.4]
  assign RetimeWrapper_60_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@11399.4]
  assign RetimeWrapper_60_io_in = _T_1416 & io_rPort_15_en_0; // @[package.scala 94:16:@11398.4]
  assign RetimeWrapper_61_clock = clock; // @[:@11404.4]
  assign RetimeWrapper_61_reset = reset; // @[:@11405.4]
  assign RetimeWrapper_61_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@11407.4]
  assign RetimeWrapper_61_io_in = _T_1640 & io_rPort_15_en_0; // @[package.scala 94:16:@11406.4]
  assign RetimeWrapper_62_clock = clock; // @[:@11412.4]
  assign RetimeWrapper_62_reset = reset; // @[:@11413.4]
  assign RetimeWrapper_62_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@11415.4]
  assign RetimeWrapper_62_io_in = _T_1864 & io_rPort_15_en_0; // @[package.scala 94:16:@11414.4]
  assign RetimeWrapper_63_clock = clock; // @[:@11420.4]
  assign RetimeWrapper_63_reset = reset; // @[:@11421.4]
  assign RetimeWrapper_63_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@11423.4]
  assign RetimeWrapper_63_io_in = _T_2088 & io_rPort_15_en_0; // @[package.scala 94:16:@11422.4]
  assign RetimeWrapper_64_clock = clock; // @[:@11444.4]
  assign RetimeWrapper_64_reset = reset; // @[:@11445.4]
  assign RetimeWrapper_64_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@11447.4]
  assign RetimeWrapper_64_io_in = _T_1495 & io_rPort_16_en_0; // @[package.scala 94:16:@11446.4]
  assign RetimeWrapper_65_clock = clock; // @[:@11452.4]
  assign RetimeWrapper_65_reset = reset; // @[:@11453.4]
  assign RetimeWrapper_65_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@11455.4]
  assign RetimeWrapper_65_io_in = _T_1719 & io_rPort_16_en_0; // @[package.scala 94:16:@11454.4]
  assign RetimeWrapper_66_clock = clock; // @[:@11460.4]
  assign RetimeWrapper_66_reset = reset; // @[:@11461.4]
  assign RetimeWrapper_66_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@11463.4]
  assign RetimeWrapper_66_io_in = _T_1943 & io_rPort_16_en_0; // @[package.scala 94:16:@11462.4]
  assign RetimeWrapper_67_clock = clock; // @[:@11468.4]
  assign RetimeWrapper_67_reset = reset; // @[:@11469.4]
  assign RetimeWrapper_67_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@11471.4]
  assign RetimeWrapper_67_io_in = _T_2167 & io_rPort_16_en_0; // @[package.scala 94:16:@11470.4]
  assign RetimeWrapper_68_clock = clock; // @[:@11492.4]
  assign RetimeWrapper_68_reset = reset; // @[:@11493.4]
  assign RetimeWrapper_68_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@11495.4]
  assign RetimeWrapper_68_io_in = _T_1421 & io_rPort_17_en_0; // @[package.scala 94:16:@11494.4]
  assign RetimeWrapper_69_clock = clock; // @[:@11500.4]
  assign RetimeWrapper_69_reset = reset; // @[:@11501.4]
  assign RetimeWrapper_69_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@11503.4]
  assign RetimeWrapper_69_io_in = _T_1645 & io_rPort_17_en_0; // @[package.scala 94:16:@11502.4]
  assign RetimeWrapper_70_clock = clock; // @[:@11508.4]
  assign RetimeWrapper_70_reset = reset; // @[:@11509.4]
  assign RetimeWrapper_70_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@11511.4]
  assign RetimeWrapper_70_io_in = _T_1869 & io_rPort_17_en_0; // @[package.scala 94:16:@11510.4]
  assign RetimeWrapper_71_clock = clock; // @[:@11516.4]
  assign RetimeWrapper_71_reset = reset; // @[:@11517.4]
  assign RetimeWrapper_71_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@11519.4]
  assign RetimeWrapper_71_io_in = _T_2093 & io_rPort_17_en_0; // @[package.scala 94:16:@11518.4]
  assign RetimeWrapper_72_clock = clock; // @[:@11540.4]
  assign RetimeWrapper_72_reset = reset; // @[:@11541.4]
  assign RetimeWrapper_72_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@11543.4]
  assign RetimeWrapper_72_io_in = _T_1500 & io_rPort_18_en_0; // @[package.scala 94:16:@11542.4]
  assign RetimeWrapper_73_clock = clock; // @[:@11548.4]
  assign RetimeWrapper_73_reset = reset; // @[:@11549.4]
  assign RetimeWrapper_73_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@11551.4]
  assign RetimeWrapper_73_io_in = _T_1724 & io_rPort_18_en_0; // @[package.scala 94:16:@11550.4]
  assign RetimeWrapper_74_clock = clock; // @[:@11556.4]
  assign RetimeWrapper_74_reset = reset; // @[:@11557.4]
  assign RetimeWrapper_74_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@11559.4]
  assign RetimeWrapper_74_io_in = _T_1948 & io_rPort_18_en_0; // @[package.scala 94:16:@11558.4]
  assign RetimeWrapper_75_clock = clock; // @[:@11564.4]
  assign RetimeWrapper_75_reset = reset; // @[:@11565.4]
  assign RetimeWrapper_75_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@11567.4]
  assign RetimeWrapper_75_io_in = _T_2172 & io_rPort_18_en_0; // @[package.scala 94:16:@11566.4]
  assign RetimeWrapper_76_clock = clock; // @[:@11588.4]
  assign RetimeWrapper_76_reset = reset; // @[:@11589.4]
  assign RetimeWrapper_76_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@11591.4]
  assign RetimeWrapper_76_io_in = _T_1505 & io_rPort_19_en_0; // @[package.scala 94:16:@11590.4]
  assign RetimeWrapper_77_clock = clock; // @[:@11596.4]
  assign RetimeWrapper_77_reset = reset; // @[:@11597.4]
  assign RetimeWrapper_77_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@11599.4]
  assign RetimeWrapper_77_io_in = _T_1729 & io_rPort_19_en_0; // @[package.scala 94:16:@11598.4]
  assign RetimeWrapper_78_clock = clock; // @[:@11604.4]
  assign RetimeWrapper_78_reset = reset; // @[:@11605.4]
  assign RetimeWrapper_78_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@11607.4]
  assign RetimeWrapper_78_io_in = _T_1953 & io_rPort_19_en_0; // @[package.scala 94:16:@11606.4]
  assign RetimeWrapper_79_clock = clock; // @[:@11612.4]
  assign RetimeWrapper_79_reset = reset; // @[:@11613.4]
  assign RetimeWrapper_79_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@11615.4]
  assign RetimeWrapper_79_io_in = _T_2177 & io_rPort_19_en_0; // @[package.scala 94:16:@11614.4]
  assign RetimeWrapper_80_clock = clock; // @[:@11636.4]
  assign RetimeWrapper_80_reset = reset; // @[:@11637.4]
  assign RetimeWrapper_80_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@11639.4]
  assign RetimeWrapper_80_io_in = _T_1335 & io_rPort_20_en_0; // @[package.scala 94:16:@11638.4]
  assign RetimeWrapper_81_clock = clock; // @[:@11644.4]
  assign RetimeWrapper_81_reset = reset; // @[:@11645.4]
  assign RetimeWrapper_81_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@11647.4]
  assign RetimeWrapper_81_io_in = _T_1559 & io_rPort_20_en_0; // @[package.scala 94:16:@11646.4]
  assign RetimeWrapper_82_clock = clock; // @[:@11652.4]
  assign RetimeWrapper_82_reset = reset; // @[:@11653.4]
  assign RetimeWrapper_82_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@11655.4]
  assign RetimeWrapper_82_io_in = _T_1783 & io_rPort_20_en_0; // @[package.scala 94:16:@11654.4]
  assign RetimeWrapper_83_clock = clock; // @[:@11660.4]
  assign RetimeWrapper_83_reset = reset; // @[:@11661.4]
  assign RetimeWrapper_83_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@11663.4]
  assign RetimeWrapper_83_io_in = _T_2007 & io_rPort_20_en_0; // @[package.scala 94:16:@11662.4]
  assign RetimeWrapper_84_clock = clock; // @[:@11684.4]
  assign RetimeWrapper_84_reset = reset; // @[:@11685.4]
  assign RetimeWrapper_84_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@11687.4]
  assign RetimeWrapper_84_io_in = _T_1373 & io_rPort_21_en_0; // @[package.scala 94:16:@11686.4]
  assign RetimeWrapper_85_clock = clock; // @[:@11692.4]
  assign RetimeWrapper_85_reset = reset; // @[:@11693.4]
  assign RetimeWrapper_85_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@11695.4]
  assign RetimeWrapper_85_io_in = _T_1597 & io_rPort_21_en_0; // @[package.scala 94:16:@11694.4]
  assign RetimeWrapper_86_clock = clock; // @[:@11700.4]
  assign RetimeWrapper_86_reset = reset; // @[:@11701.4]
  assign RetimeWrapper_86_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@11703.4]
  assign RetimeWrapper_86_io_in = _T_1821 & io_rPort_21_en_0; // @[package.scala 94:16:@11702.4]
  assign RetimeWrapper_87_clock = clock; // @[:@11708.4]
  assign RetimeWrapper_87_reset = reset; // @[:@11709.4]
  assign RetimeWrapper_87_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@11711.4]
  assign RetimeWrapper_87_io_in = _T_2045 & io_rPort_21_en_0; // @[package.scala 94:16:@11710.4]
  assign RetimeWrapper_88_clock = clock; // @[:@11732.4]
  assign RetimeWrapper_88_reset = reset; // @[:@11733.4]
  assign RetimeWrapper_88_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@11735.4]
  assign RetimeWrapper_88_io_in = _T_1426 & io_rPort_22_en_0; // @[package.scala 94:16:@11734.4]
  assign RetimeWrapper_89_clock = clock; // @[:@11740.4]
  assign RetimeWrapper_89_reset = reset; // @[:@11741.4]
  assign RetimeWrapper_89_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@11743.4]
  assign RetimeWrapper_89_io_in = _T_1650 & io_rPort_22_en_0; // @[package.scala 94:16:@11742.4]
  assign RetimeWrapper_90_clock = clock; // @[:@11748.4]
  assign RetimeWrapper_90_reset = reset; // @[:@11749.4]
  assign RetimeWrapper_90_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@11751.4]
  assign RetimeWrapper_90_io_in = _T_1874 & io_rPort_22_en_0; // @[package.scala 94:16:@11750.4]
  assign RetimeWrapper_91_clock = clock; // @[:@11756.4]
  assign RetimeWrapper_91_reset = reset; // @[:@11757.4]
  assign RetimeWrapper_91_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@11759.4]
  assign RetimeWrapper_91_io_in = _T_2098 & io_rPort_22_en_0; // @[package.scala 94:16:@11758.4]
  assign RetimeWrapper_92_clock = clock; // @[:@11780.4]
  assign RetimeWrapper_92_reset = reset; // @[:@11781.4]
  assign RetimeWrapper_92_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@11783.4]
  assign RetimeWrapper_92_io_in = _T_1431 & io_rPort_23_en_0; // @[package.scala 94:16:@11782.4]
  assign RetimeWrapper_93_clock = clock; // @[:@11788.4]
  assign RetimeWrapper_93_reset = reset; // @[:@11789.4]
  assign RetimeWrapper_93_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@11791.4]
  assign RetimeWrapper_93_io_in = _T_1655 & io_rPort_23_en_0; // @[package.scala 94:16:@11790.4]
  assign RetimeWrapper_94_clock = clock; // @[:@11796.4]
  assign RetimeWrapper_94_reset = reset; // @[:@11797.4]
  assign RetimeWrapper_94_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@11799.4]
  assign RetimeWrapper_94_io_in = _T_1879 & io_rPort_23_en_0; // @[package.scala 94:16:@11798.4]
  assign RetimeWrapper_95_clock = clock; // @[:@11804.4]
  assign RetimeWrapper_95_reset = reset; // @[:@11805.4]
  assign RetimeWrapper_95_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@11807.4]
  assign RetimeWrapper_95_io_in = _T_2103 & io_rPort_23_en_0; // @[package.scala 94:16:@11806.4]
endmodule
module StickySelects_16( // @[:@13335.2]
  input   clock, // @[:@13336.4]
  input   reset, // @[:@13337.4]
  input   io_ins_0, // @[:@13338.4]
  input   io_ins_1, // @[:@13338.4]
  input   io_ins_2, // @[:@13338.4]
  output  io_outs_0, // @[:@13338.4]
  output  io_outs_1, // @[:@13338.4]
  output  io_outs_2 // @[:@13338.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@13340.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@13341.4]
  wire  _T_22; // @[StickySelects.scala 24:52:@13342.4]
  wire  _T_23; // @[StickySelects.scala 24:21:@13343.4]
  reg  _T_26; // @[StickySelects.scala 21:22:@13345.4]
  reg [31:0] _RAND_1;
  wire  _T_27; // @[StickySelects.scala 22:54:@13346.4]
  wire  _T_29; // @[StickySelects.scala 24:52:@13347.4]
  wire  _T_30; // @[StickySelects.scala 24:21:@13348.4]
  reg  _T_33; // @[StickySelects.scala 21:22:@13350.4]
  reg [31:0] _RAND_2;
  wire  _T_34; // @[StickySelects.scala 22:54:@13351.4]
  wire  _T_36; // @[StickySelects.scala 24:52:@13352.4]
  wire  _T_37; // @[StickySelects.scala 24:21:@13353.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@13341.4]
  assign _T_22 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@13342.4]
  assign _T_23 = _T_20 ? 1'h0 : _T_22; // @[StickySelects.scala 24:21:@13343.4]
  assign _T_27 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@13346.4]
  assign _T_29 = io_ins_1 | _T_26; // @[StickySelects.scala 24:52:@13347.4]
  assign _T_30 = _T_27 ? 1'h0 : _T_29; // @[StickySelects.scala 24:21:@13348.4]
  assign _T_34 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@13351.4]
  assign _T_36 = io_ins_2 | _T_33; // @[StickySelects.scala 24:52:@13352.4]
  assign _T_37 = _T_34 ? 1'h0 : _T_36; // @[StickySelects.scala 24:21:@13353.4]
  assign io_outs_0 = _T_20 ? 1'h0 : _T_22; // @[StickySelects.scala 28:52:@13355.4]
  assign io_outs_1 = _T_27 ? 1'h0 : _T_29; // @[StickySelects.scala 28:52:@13356.4]
  assign io_outs_2 = _T_34 ? 1'h0 : _T_36; // @[StickySelects.scala 28:52:@13357.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_33 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_20) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_22;
      end
    end
    if (reset) begin
      _T_26 <= 1'h0;
    end else begin
      if (_T_27) begin
        _T_26 <= 1'h0;
      end else begin
        _T_26 <= _T_29;
      end
    end
    if (reset) begin
      _T_33 <= 1'h0;
    end else begin
      if (_T_34) begin
        _T_33 <= 1'h0;
      end else begin
        _T_33 <= _T_36;
      end
    end
  end
endmodule
module StickySelects_19( // @[:@13407.2]
  input   clock, // @[:@13408.4]
  input   reset, // @[:@13409.4]
  input   io_ins_0, // @[:@13410.4]
  input   io_ins_1, // @[:@13410.4]
  input   io_ins_2, // @[:@13410.4]
  input   io_ins_3, // @[:@13410.4]
  input   io_ins_4, // @[:@13410.4]
  input   io_ins_5, // @[:@13410.4]
  output  io_outs_0, // @[:@13410.4]
  output  io_outs_1, // @[:@13410.4]
  output  io_outs_2, // @[:@13410.4]
  output  io_outs_3, // @[:@13410.4]
  output  io_outs_4, // @[:@13410.4]
  output  io_outs_5 // @[:@13410.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@13412.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@13413.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@13414.4]
  wire  _T_22; // @[StickySelects.scala 22:54:@13415.4]
  wire  _T_23; // @[StickySelects.scala 22:54:@13416.4]
  wire  _T_25; // @[StickySelects.scala 24:52:@13417.4]
  wire  _T_26; // @[StickySelects.scala 24:21:@13418.4]
  reg  _T_29; // @[StickySelects.scala 21:22:@13420.4]
  reg [31:0] _RAND_1;
  wire  _T_30; // @[StickySelects.scala 22:54:@13421.4]
  wire  _T_31; // @[StickySelects.scala 22:54:@13422.4]
  wire  _T_32; // @[StickySelects.scala 22:54:@13423.4]
  wire  _T_33; // @[StickySelects.scala 22:54:@13424.4]
  wire  _T_35; // @[StickySelects.scala 24:52:@13425.4]
  wire  _T_36; // @[StickySelects.scala 24:21:@13426.4]
  reg  _T_39; // @[StickySelects.scala 21:22:@13428.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[StickySelects.scala 22:54:@13429.4]
  wire  _T_41; // @[StickySelects.scala 22:54:@13430.4]
  wire  _T_42; // @[StickySelects.scala 22:54:@13431.4]
  wire  _T_43; // @[StickySelects.scala 22:54:@13432.4]
  wire  _T_45; // @[StickySelects.scala 24:52:@13433.4]
  wire  _T_46; // @[StickySelects.scala 24:21:@13434.4]
  reg  _T_49; // @[StickySelects.scala 21:22:@13436.4]
  reg [31:0] _RAND_3;
  wire  _T_51; // @[StickySelects.scala 22:54:@13438.4]
  wire  _T_52; // @[StickySelects.scala 22:54:@13439.4]
  wire  _T_53; // @[StickySelects.scala 22:54:@13440.4]
  wire  _T_55; // @[StickySelects.scala 24:52:@13441.4]
  wire  _T_56; // @[StickySelects.scala 24:21:@13442.4]
  reg  _T_59; // @[StickySelects.scala 21:22:@13444.4]
  reg [31:0] _RAND_4;
  wire  _T_62; // @[StickySelects.scala 22:54:@13447.4]
  wire  _T_63; // @[StickySelects.scala 22:54:@13448.4]
  wire  _T_65; // @[StickySelects.scala 24:52:@13449.4]
  wire  _T_66; // @[StickySelects.scala 24:21:@13450.4]
  reg  _T_69; // @[StickySelects.scala 21:22:@13452.4]
  reg [31:0] _RAND_5;
  wire  _T_73; // @[StickySelects.scala 22:54:@13456.4]
  wire  _T_75; // @[StickySelects.scala 24:52:@13457.4]
  wire  _T_76; // @[StickySelects.scala 24:21:@13458.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@13413.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@13414.4]
  assign _T_22 = _T_21 | io_ins_4; // @[StickySelects.scala 22:54:@13415.4]
  assign _T_23 = _T_22 | io_ins_5; // @[StickySelects.scala 22:54:@13416.4]
  assign _T_25 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@13417.4]
  assign _T_26 = _T_23 ? 1'h0 : _T_25; // @[StickySelects.scala 24:21:@13418.4]
  assign _T_30 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@13421.4]
  assign _T_31 = _T_30 | io_ins_3; // @[StickySelects.scala 22:54:@13422.4]
  assign _T_32 = _T_31 | io_ins_4; // @[StickySelects.scala 22:54:@13423.4]
  assign _T_33 = _T_32 | io_ins_5; // @[StickySelects.scala 22:54:@13424.4]
  assign _T_35 = io_ins_1 | _T_29; // @[StickySelects.scala 24:52:@13425.4]
  assign _T_36 = _T_33 ? 1'h0 : _T_35; // @[StickySelects.scala 24:21:@13426.4]
  assign _T_40 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@13429.4]
  assign _T_41 = _T_40 | io_ins_3; // @[StickySelects.scala 22:54:@13430.4]
  assign _T_42 = _T_41 | io_ins_4; // @[StickySelects.scala 22:54:@13431.4]
  assign _T_43 = _T_42 | io_ins_5; // @[StickySelects.scala 22:54:@13432.4]
  assign _T_45 = io_ins_2 | _T_39; // @[StickySelects.scala 24:52:@13433.4]
  assign _T_46 = _T_43 ? 1'h0 : _T_45; // @[StickySelects.scala 24:21:@13434.4]
  assign _T_51 = _T_40 | io_ins_2; // @[StickySelects.scala 22:54:@13438.4]
  assign _T_52 = _T_51 | io_ins_4; // @[StickySelects.scala 22:54:@13439.4]
  assign _T_53 = _T_52 | io_ins_5; // @[StickySelects.scala 22:54:@13440.4]
  assign _T_55 = io_ins_3 | _T_49; // @[StickySelects.scala 24:52:@13441.4]
  assign _T_56 = _T_53 ? 1'h0 : _T_55; // @[StickySelects.scala 24:21:@13442.4]
  assign _T_62 = _T_51 | io_ins_3; // @[StickySelects.scala 22:54:@13447.4]
  assign _T_63 = _T_62 | io_ins_5; // @[StickySelects.scala 22:54:@13448.4]
  assign _T_65 = io_ins_4 | _T_59; // @[StickySelects.scala 24:52:@13449.4]
  assign _T_66 = _T_63 ? 1'h0 : _T_65; // @[StickySelects.scala 24:21:@13450.4]
  assign _T_73 = _T_62 | io_ins_4; // @[StickySelects.scala 22:54:@13456.4]
  assign _T_75 = io_ins_5 | _T_69; // @[StickySelects.scala 24:52:@13457.4]
  assign _T_76 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 24:21:@13458.4]
  assign io_outs_0 = _T_23 ? 1'h0 : _T_25; // @[StickySelects.scala 28:52:@13460.4]
  assign io_outs_1 = _T_33 ? 1'h0 : _T_35; // @[StickySelects.scala 28:52:@13461.4]
  assign io_outs_2 = _T_43 ? 1'h0 : _T_45; // @[StickySelects.scala 28:52:@13462.4]
  assign io_outs_3 = _T_53 ? 1'h0 : _T_55; // @[StickySelects.scala 28:52:@13463.4]
  assign io_outs_4 = _T_63 ? 1'h0 : _T_65; // @[StickySelects.scala 28:52:@13464.4]
  assign io_outs_5 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 28:52:@13465.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_29 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_39 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_49 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_59 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_69 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_23) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_25;
      end
    end
    if (reset) begin
      _T_29 <= 1'h0;
    end else begin
      if (_T_33) begin
        _T_29 <= 1'h0;
      end else begin
        _T_29 <= _T_35;
      end
    end
    if (reset) begin
      _T_39 <= 1'h0;
    end else begin
      if (_T_43) begin
        _T_39 <= 1'h0;
      end else begin
        _T_39 <= _T_45;
      end
    end
    if (reset) begin
      _T_49 <= 1'h0;
    end else begin
      if (_T_53) begin
        _T_49 <= 1'h0;
      end else begin
        _T_49 <= _T_55;
      end
    end
    if (reset) begin
      _T_59 <= 1'h0;
    end else begin
      if (_T_63) begin
        _T_59 <= 1'h0;
      end else begin
        _T_59 <= _T_65;
      end
    end
    if (reset) begin
      _T_69 <= 1'h0;
    end else begin
      if (_T_73) begin
        _T_69 <= 1'h0;
      end else begin
        _T_69 <= _T_75;
      end
    end
  end
endmodule
module x525_lb2_0( // @[:@15783.2]
  input        clock, // @[:@15784.4]
  input        reset, // @[:@15785.4]
  input  [2:0] io_rPort_14_banks_0, // @[:@15786.4]
  input        io_rPort_14_ofs_0, // @[:@15786.4]
  input        io_rPort_14_en_0, // @[:@15786.4]
  input        io_rPort_14_backpressure, // @[:@15786.4]
  output [7:0] io_rPort_14_output_0, // @[:@15786.4]
  input  [2:0] io_rPort_13_banks_0, // @[:@15786.4]
  input        io_rPort_13_ofs_0, // @[:@15786.4]
  input        io_rPort_13_en_0, // @[:@15786.4]
  input        io_rPort_13_backpressure, // @[:@15786.4]
  output [7:0] io_rPort_13_output_0, // @[:@15786.4]
  input  [2:0] io_rPort_12_banks_0, // @[:@15786.4]
  input        io_rPort_12_ofs_0, // @[:@15786.4]
  input        io_rPort_12_en_0, // @[:@15786.4]
  input        io_rPort_12_backpressure, // @[:@15786.4]
  output [7:0] io_rPort_12_output_0, // @[:@15786.4]
  input  [2:0] io_rPort_11_banks_0, // @[:@15786.4]
  input        io_rPort_11_ofs_0, // @[:@15786.4]
  input        io_rPort_11_en_0, // @[:@15786.4]
  input        io_rPort_11_backpressure, // @[:@15786.4]
  output [7:0] io_rPort_11_output_0, // @[:@15786.4]
  input  [2:0] io_rPort_10_banks_0, // @[:@15786.4]
  input        io_rPort_10_ofs_0, // @[:@15786.4]
  input        io_rPort_10_en_0, // @[:@15786.4]
  input        io_rPort_10_backpressure, // @[:@15786.4]
  output [7:0] io_rPort_10_output_0, // @[:@15786.4]
  input  [2:0] io_rPort_9_banks_0, // @[:@15786.4]
  input        io_rPort_9_ofs_0, // @[:@15786.4]
  input        io_rPort_9_en_0, // @[:@15786.4]
  input        io_rPort_9_backpressure, // @[:@15786.4]
  output [7:0] io_rPort_9_output_0, // @[:@15786.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@15786.4]
  input        io_rPort_8_ofs_0, // @[:@15786.4]
  input        io_rPort_8_en_0, // @[:@15786.4]
  input        io_rPort_8_backpressure, // @[:@15786.4]
  output [7:0] io_rPort_8_output_0, // @[:@15786.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@15786.4]
  input        io_rPort_7_ofs_0, // @[:@15786.4]
  input        io_rPort_7_en_0, // @[:@15786.4]
  input        io_rPort_7_backpressure, // @[:@15786.4]
  output [7:0] io_rPort_7_output_0, // @[:@15786.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@15786.4]
  input        io_rPort_6_ofs_0, // @[:@15786.4]
  input        io_rPort_6_en_0, // @[:@15786.4]
  input        io_rPort_6_backpressure, // @[:@15786.4]
  output [7:0] io_rPort_6_output_0, // @[:@15786.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@15786.4]
  input        io_rPort_5_ofs_0, // @[:@15786.4]
  input        io_rPort_5_en_0, // @[:@15786.4]
  input        io_rPort_5_backpressure, // @[:@15786.4]
  output [7:0] io_rPort_5_output_0, // @[:@15786.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@15786.4]
  input        io_rPort_4_ofs_0, // @[:@15786.4]
  input        io_rPort_4_en_0, // @[:@15786.4]
  input        io_rPort_4_backpressure, // @[:@15786.4]
  output [7:0] io_rPort_4_output_0, // @[:@15786.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@15786.4]
  input        io_rPort_3_ofs_0, // @[:@15786.4]
  input        io_rPort_3_en_0, // @[:@15786.4]
  input        io_rPort_3_backpressure, // @[:@15786.4]
  output [7:0] io_rPort_3_output_0, // @[:@15786.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@15786.4]
  input        io_rPort_2_ofs_0, // @[:@15786.4]
  input        io_rPort_2_en_0, // @[:@15786.4]
  input        io_rPort_2_backpressure, // @[:@15786.4]
  output [7:0] io_rPort_2_output_0, // @[:@15786.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@15786.4]
  input        io_rPort_1_ofs_0, // @[:@15786.4]
  input        io_rPort_1_en_0, // @[:@15786.4]
  input        io_rPort_1_backpressure, // @[:@15786.4]
  output [7:0] io_rPort_1_output_0, // @[:@15786.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@15786.4]
  input        io_rPort_0_ofs_0, // @[:@15786.4]
  input        io_rPort_0_en_0, // @[:@15786.4]
  input        io_rPort_0_backpressure, // @[:@15786.4]
  output [7:0] io_rPort_0_output_0, // @[:@15786.4]
  input  [2:0] io_wPort_7_banks_0, // @[:@15786.4]
  input        io_wPort_7_ofs_0, // @[:@15786.4]
  input  [7:0] io_wPort_7_data_0, // @[:@15786.4]
  input        io_wPort_7_en_0, // @[:@15786.4]
  input  [2:0] io_wPort_6_banks_0, // @[:@15786.4]
  input        io_wPort_6_ofs_0, // @[:@15786.4]
  input  [7:0] io_wPort_6_data_0, // @[:@15786.4]
  input        io_wPort_6_en_0, // @[:@15786.4]
  input  [2:0] io_wPort_5_banks_0, // @[:@15786.4]
  input        io_wPort_5_ofs_0, // @[:@15786.4]
  input  [7:0] io_wPort_5_data_0, // @[:@15786.4]
  input        io_wPort_5_en_0, // @[:@15786.4]
  input  [2:0] io_wPort_4_banks_0, // @[:@15786.4]
  input        io_wPort_4_ofs_0, // @[:@15786.4]
  input  [7:0] io_wPort_4_data_0, // @[:@15786.4]
  input        io_wPort_4_en_0, // @[:@15786.4]
  input  [2:0] io_wPort_3_banks_0, // @[:@15786.4]
  input        io_wPort_3_ofs_0, // @[:@15786.4]
  input  [7:0] io_wPort_3_data_0, // @[:@15786.4]
  input        io_wPort_3_en_0, // @[:@15786.4]
  input  [2:0] io_wPort_2_banks_0, // @[:@15786.4]
  input        io_wPort_2_ofs_0, // @[:@15786.4]
  input  [7:0] io_wPort_2_data_0, // @[:@15786.4]
  input        io_wPort_2_en_0, // @[:@15786.4]
  input  [2:0] io_wPort_1_banks_0, // @[:@15786.4]
  input        io_wPort_1_ofs_0, // @[:@15786.4]
  input  [7:0] io_wPort_1_data_0, // @[:@15786.4]
  input        io_wPort_1_en_0, // @[:@15786.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@15786.4]
  input        io_wPort_0_ofs_0, // @[:@15786.4]
  input  [7:0] io_wPort_0_data_0, // @[:@15786.4]
  input        io_wPort_0_en_0 // @[:@15786.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@15943.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@15943.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15943.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15943.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15943.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@15943.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@15943.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@15943.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@15959.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@15959.4]
  wire  Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15959.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15959.4]
  wire  Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15959.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@15959.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@15959.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@15959.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@15975.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@15975.4]
  wire  Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15975.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15975.4]
  wire  Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15975.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@15975.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@15975.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@15975.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@15991.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@15991.4]
  wire  Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@15991.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@15991.4]
  wire  Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@15991.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@15991.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@15991.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@15991.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@16007.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@16007.4]
  wire  Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@16007.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@16007.4]
  wire  Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@16007.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@16007.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@16007.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@16007.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@16023.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@16023.4]
  wire  Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@16023.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@16023.4]
  wire  Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@16023.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@16023.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@16023.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@16023.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@16039.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@16039.4]
  wire  Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@16039.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@16039.4]
  wire  Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@16039.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@16039.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@16039.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@16039.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@16055.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@16055.4]
  wire  Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@16055.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@16055.4]
  wire  Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@16055.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@16055.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@16055.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@16055.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@16071.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@16071.4]
  wire  Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@16071.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@16071.4]
  wire  Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@16071.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@16071.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@16071.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@16071.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@16087.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@16087.4]
  wire  Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@16087.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@16087.4]
  wire  Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@16087.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@16087.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@16087.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@16087.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@16103.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@16103.4]
  wire  Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@16103.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@16103.4]
  wire  Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@16103.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@16103.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@16103.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@16103.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@16119.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@16119.4]
  wire  Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@16119.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@16119.4]
  wire  Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@16119.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@16119.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@16119.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@16119.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@16135.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@16135.4]
  wire  Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@16135.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@16135.4]
  wire  Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@16135.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@16135.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@16135.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@16135.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@16151.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@16151.4]
  wire  Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@16151.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@16151.4]
  wire  Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@16151.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@16151.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@16151.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@16151.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@16167.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@16167.4]
  wire  Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@16167.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@16167.4]
  wire  Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@16167.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@16167.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@16167.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@16167.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@16183.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@16183.4]
  wire  Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@16183.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@16183.4]
  wire  Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@16183.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@16183.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@16183.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@16183.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@16480.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@16480.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@16480.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@16480.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@16480.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@16480.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@16480.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@16480.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@16512.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@16512.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@16512.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@16512.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@16512.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@16512.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@16512.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@16512.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@16544.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@16544.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@16544.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@16544.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@16544.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@16544.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@16544.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@16544.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@16585.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@16585.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@16585.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@16585.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@16585.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@16585.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@16585.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@16585.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@16585.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@16585.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@16585.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@16585.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@16585.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@16585.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@16632.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@16632.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@16632.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@16632.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@16632.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@16632.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@16632.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@16632.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@16664.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@16664.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@16664.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@16664.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@16664.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@16664.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@16664.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@16664.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@16696.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@16696.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@16696.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@16696.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@16696.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@16696.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@16696.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@16696.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@16737.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@16737.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@16737.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@16737.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@16737.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@16737.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@16737.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@16737.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@16737.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@16737.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@16737.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@16737.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@16737.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@16737.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@16784.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@16784.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@16784.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@16784.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@16784.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@16784.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@16784.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@16784.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@16816.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@16816.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@16816.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@16816.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@16816.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@16816.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@16816.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@16816.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@16848.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@16848.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@16848.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@16848.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@16848.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@16848.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@16848.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@16848.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@16889.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@16889.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@16889.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@16889.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@16889.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@16889.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@16889.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@16889.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@16889.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@16889.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@16889.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@16889.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@16889.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@16889.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@16936.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@16936.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@16936.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@16936.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 121:29:@16936.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@16936.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@16936.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 121:29:@16936.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@16968.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@16968.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@16968.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@16968.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 121:29:@16968.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@16968.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@16968.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 121:29:@16968.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@17000.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@17000.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@17000.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@17000.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 121:29:@17000.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@17000.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@17000.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 121:29:@17000.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@17041.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@17041.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@17041.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@17041.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@17041.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@17041.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 121:29:@17041.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 121:29:@17041.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@17041.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@17041.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@17041.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@17041.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 121:29:@17041.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 121:29:@17041.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@17092.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@17092.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@17092.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@17092.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@17092.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@17100.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@17100.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@17100.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@17100.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@17100.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@17108.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@17108.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@17108.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@17108.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@17108.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@17116.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@17116.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@17116.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@17116.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@17116.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@17140.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@17140.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@17140.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@17140.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@17140.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@17148.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@17148.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@17148.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@17148.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@17148.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@17156.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@17156.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@17156.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@17156.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@17156.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@17164.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@17164.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@17164.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@17164.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@17164.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@17188.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@17188.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@17188.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@17188.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@17188.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@17196.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@17196.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@17196.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@17196.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@17196.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@17204.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@17204.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@17204.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@17204.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@17204.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@17212.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@17212.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@17212.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@17212.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@17212.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@17236.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@17236.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@17236.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@17236.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@17236.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@17244.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@17244.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@17244.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@17244.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@17244.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@17252.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@17252.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@17252.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@17252.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@17252.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@17260.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@17260.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@17260.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@17260.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@17260.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@17284.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@17284.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@17284.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@17284.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@17284.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@17292.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@17292.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@17292.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@17292.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@17292.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@17300.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@17300.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@17300.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@17300.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@17300.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@17308.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@17308.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@17308.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@17308.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@17308.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@17332.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@17332.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@17332.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@17332.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@17332.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@17340.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@17340.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@17340.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@17340.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@17340.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@17348.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@17348.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@17348.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@17348.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@17348.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@17356.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@17356.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@17356.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@17356.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@17356.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@17380.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@17380.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@17380.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@17380.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@17380.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@17388.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@17388.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@17388.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@17388.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@17388.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@17396.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@17396.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@17396.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@17396.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@17396.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@17404.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@17404.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@17404.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@17404.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@17404.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@17428.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@17428.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@17428.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@17428.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@17428.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@17436.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@17436.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@17436.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@17436.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@17436.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@17444.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@17444.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@17444.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@17444.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@17444.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@17452.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@17452.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@17452.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@17452.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@17452.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@17476.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@17476.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@17476.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@17476.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@17476.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@17484.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@17484.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@17484.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@17484.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@17484.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@17492.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@17492.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@17492.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@17492.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@17492.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@17500.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@17500.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@17500.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@17500.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@17500.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@17524.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@17524.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@17524.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@17524.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@17524.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@17532.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@17532.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@17532.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@17532.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@17532.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@17540.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@17540.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@17540.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@17540.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@17540.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@17548.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@17548.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@17548.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@17548.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@17548.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@17572.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@17572.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@17572.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@17572.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@17572.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@17580.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@17580.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@17580.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@17580.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@17580.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@17588.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@17588.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@17588.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@17588.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@17588.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@17596.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@17596.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@17596.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@17596.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@17596.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@17620.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@17620.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@17620.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@17620.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@17620.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@17628.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@17628.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@17628.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@17628.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@17628.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@17636.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@17636.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@17636.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@17636.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@17636.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@17644.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@17644.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@17644.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@17644.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@17644.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@17668.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@17668.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@17668.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@17668.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@17668.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@17676.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@17676.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@17676.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@17676.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@17676.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@17684.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@17684.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@17684.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@17684.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@17684.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@17692.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@17692.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@17692.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@17692.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@17692.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@17716.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@17716.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@17716.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@17716.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@17716.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@17724.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@17724.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@17724.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@17724.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@17724.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@17732.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@17732.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@17732.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@17732.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@17732.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@17740.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@17740.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@17740.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@17740.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@17740.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@17764.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@17764.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@17764.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@17764.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@17764.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@17772.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@17772.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@17772.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@17772.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@17772.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@17780.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@17780.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@17780.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@17780.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@17780.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@17788.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@17788.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@17788.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@17788.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@17788.4]
  wire  _T_762; // @[MemPrimitives.scala 82:210:@16199.4]
  wire  _T_765; // @[MemPrimitives.scala 83:102:@16201.4]
  wire  _T_767; // @[MemPrimitives.scala 82:210:@16202.4]
  wire  _T_770; // @[MemPrimitives.scala 83:102:@16204.4]
  wire [9:0] _T_772; // @[Cat.scala 30:58:@16206.4]
  wire [9:0] _T_774; // @[Cat.scala 30:58:@16208.4]
  wire [9:0] _T_775; // @[Mux.scala 31:69:@16209.4]
  wire  _T_780; // @[MemPrimitives.scala 82:210:@16216.4]
  wire  _T_783; // @[MemPrimitives.scala 83:102:@16218.4]
  wire  _T_785; // @[MemPrimitives.scala 82:210:@16219.4]
  wire  _T_788; // @[MemPrimitives.scala 83:102:@16221.4]
  wire [9:0] _T_790; // @[Cat.scala 30:58:@16223.4]
  wire [9:0] _T_792; // @[Cat.scala 30:58:@16225.4]
  wire [9:0] _T_793; // @[Mux.scala 31:69:@16226.4]
  wire  _T_798; // @[MemPrimitives.scala 82:210:@16233.4]
  wire  _T_801; // @[MemPrimitives.scala 83:102:@16235.4]
  wire  _T_803; // @[MemPrimitives.scala 82:210:@16236.4]
  wire  _T_806; // @[MemPrimitives.scala 83:102:@16238.4]
  wire [9:0] _T_808; // @[Cat.scala 30:58:@16240.4]
  wire [9:0] _T_810; // @[Cat.scala 30:58:@16242.4]
  wire [9:0] _T_811; // @[Mux.scala 31:69:@16243.4]
  wire  _T_816; // @[MemPrimitives.scala 82:210:@16250.4]
  wire  _T_819; // @[MemPrimitives.scala 83:102:@16252.4]
  wire  _T_821; // @[MemPrimitives.scala 82:210:@16253.4]
  wire  _T_824; // @[MemPrimitives.scala 83:102:@16255.4]
  wire [9:0] _T_826; // @[Cat.scala 30:58:@16257.4]
  wire [9:0] _T_828; // @[Cat.scala 30:58:@16259.4]
  wire [9:0] _T_829; // @[Mux.scala 31:69:@16260.4]
  wire  _T_834; // @[MemPrimitives.scala 82:210:@16267.4]
  wire  _T_837; // @[MemPrimitives.scala 83:102:@16269.4]
  wire  _T_839; // @[MemPrimitives.scala 82:210:@16270.4]
  wire  _T_842; // @[MemPrimitives.scala 83:102:@16272.4]
  wire [9:0] _T_844; // @[Cat.scala 30:58:@16274.4]
  wire [9:0] _T_846; // @[Cat.scala 30:58:@16276.4]
  wire [9:0] _T_847; // @[Mux.scala 31:69:@16277.4]
  wire  _T_852; // @[MemPrimitives.scala 82:210:@16284.4]
  wire  _T_855; // @[MemPrimitives.scala 83:102:@16286.4]
  wire  _T_857; // @[MemPrimitives.scala 82:210:@16287.4]
  wire  _T_860; // @[MemPrimitives.scala 83:102:@16289.4]
  wire [9:0] _T_862; // @[Cat.scala 30:58:@16291.4]
  wire [9:0] _T_864; // @[Cat.scala 30:58:@16293.4]
  wire [9:0] _T_865; // @[Mux.scala 31:69:@16294.4]
  wire  _T_870; // @[MemPrimitives.scala 82:210:@16301.4]
  wire  _T_873; // @[MemPrimitives.scala 83:102:@16303.4]
  wire  _T_875; // @[MemPrimitives.scala 82:210:@16304.4]
  wire  _T_878; // @[MemPrimitives.scala 83:102:@16306.4]
  wire [9:0] _T_880; // @[Cat.scala 30:58:@16308.4]
  wire [9:0] _T_882; // @[Cat.scala 30:58:@16310.4]
  wire [9:0] _T_883; // @[Mux.scala 31:69:@16311.4]
  wire  _T_888; // @[MemPrimitives.scala 82:210:@16318.4]
  wire  _T_891; // @[MemPrimitives.scala 83:102:@16320.4]
  wire  _T_893; // @[MemPrimitives.scala 82:210:@16321.4]
  wire  _T_896; // @[MemPrimitives.scala 83:102:@16323.4]
  wire [9:0] _T_898; // @[Cat.scala 30:58:@16325.4]
  wire [9:0] _T_900; // @[Cat.scala 30:58:@16327.4]
  wire [9:0] _T_901; // @[Mux.scala 31:69:@16328.4]
  wire  _T_906; // @[MemPrimitives.scala 82:210:@16335.4]
  wire  _T_909; // @[MemPrimitives.scala 83:102:@16337.4]
  wire  _T_911; // @[MemPrimitives.scala 82:210:@16338.4]
  wire  _T_914; // @[MemPrimitives.scala 83:102:@16340.4]
  wire [9:0] _T_916; // @[Cat.scala 30:58:@16342.4]
  wire [9:0] _T_918; // @[Cat.scala 30:58:@16344.4]
  wire [9:0] _T_919; // @[Mux.scala 31:69:@16345.4]
  wire  _T_924; // @[MemPrimitives.scala 82:210:@16352.4]
  wire  _T_927; // @[MemPrimitives.scala 83:102:@16354.4]
  wire  _T_929; // @[MemPrimitives.scala 82:210:@16355.4]
  wire  _T_932; // @[MemPrimitives.scala 83:102:@16357.4]
  wire [9:0] _T_934; // @[Cat.scala 30:58:@16359.4]
  wire [9:0] _T_936; // @[Cat.scala 30:58:@16361.4]
  wire [9:0] _T_937; // @[Mux.scala 31:69:@16362.4]
  wire  _T_942; // @[MemPrimitives.scala 82:210:@16369.4]
  wire  _T_945; // @[MemPrimitives.scala 83:102:@16371.4]
  wire  _T_947; // @[MemPrimitives.scala 82:210:@16372.4]
  wire  _T_950; // @[MemPrimitives.scala 83:102:@16374.4]
  wire [9:0] _T_952; // @[Cat.scala 30:58:@16376.4]
  wire [9:0] _T_954; // @[Cat.scala 30:58:@16378.4]
  wire [9:0] _T_955; // @[Mux.scala 31:69:@16379.4]
  wire  _T_960; // @[MemPrimitives.scala 82:210:@16386.4]
  wire  _T_963; // @[MemPrimitives.scala 83:102:@16388.4]
  wire  _T_965; // @[MemPrimitives.scala 82:210:@16389.4]
  wire  _T_968; // @[MemPrimitives.scala 83:102:@16391.4]
  wire [9:0] _T_970; // @[Cat.scala 30:58:@16393.4]
  wire [9:0] _T_972; // @[Cat.scala 30:58:@16395.4]
  wire [9:0] _T_973; // @[Mux.scala 31:69:@16396.4]
  wire  _T_978; // @[MemPrimitives.scala 82:210:@16403.4]
  wire  _T_981; // @[MemPrimitives.scala 83:102:@16405.4]
  wire  _T_983; // @[MemPrimitives.scala 82:210:@16406.4]
  wire  _T_986; // @[MemPrimitives.scala 83:102:@16408.4]
  wire [9:0] _T_988; // @[Cat.scala 30:58:@16410.4]
  wire [9:0] _T_990; // @[Cat.scala 30:58:@16412.4]
  wire [9:0] _T_991; // @[Mux.scala 31:69:@16413.4]
  wire  _T_996; // @[MemPrimitives.scala 82:210:@16420.4]
  wire  _T_999; // @[MemPrimitives.scala 83:102:@16422.4]
  wire  _T_1001; // @[MemPrimitives.scala 82:210:@16423.4]
  wire  _T_1004; // @[MemPrimitives.scala 83:102:@16425.4]
  wire [9:0] _T_1006; // @[Cat.scala 30:58:@16427.4]
  wire [9:0] _T_1008; // @[Cat.scala 30:58:@16429.4]
  wire [9:0] _T_1009; // @[Mux.scala 31:69:@16430.4]
  wire  _T_1014; // @[MemPrimitives.scala 82:210:@16437.4]
  wire  _T_1017; // @[MemPrimitives.scala 83:102:@16439.4]
  wire  _T_1019; // @[MemPrimitives.scala 82:210:@16440.4]
  wire  _T_1022; // @[MemPrimitives.scala 83:102:@16442.4]
  wire [9:0] _T_1024; // @[Cat.scala 30:58:@16444.4]
  wire [9:0] _T_1026; // @[Cat.scala 30:58:@16446.4]
  wire [9:0] _T_1027; // @[Mux.scala 31:69:@16447.4]
  wire  _T_1032; // @[MemPrimitives.scala 82:210:@16454.4]
  wire  _T_1035; // @[MemPrimitives.scala 83:102:@16456.4]
  wire  _T_1037; // @[MemPrimitives.scala 82:210:@16457.4]
  wire  _T_1040; // @[MemPrimitives.scala 83:102:@16459.4]
  wire [9:0] _T_1042; // @[Cat.scala 30:58:@16461.4]
  wire [9:0] _T_1044; // @[Cat.scala 30:58:@16463.4]
  wire [9:0] _T_1045; // @[Mux.scala 31:69:@16464.4]
  wire  _T_1050; // @[MemPrimitives.scala 110:210:@16471.4]
  wire  _T_1055; // @[MemPrimitives.scala 110:210:@16474.4]
  wire  _T_1060; // @[MemPrimitives.scala 110:210:@16477.4]
  wire  _T_1064; // @[MemPrimitives.scala 123:41:@16486.4]
  wire  _T_1065; // @[MemPrimitives.scala 123:41:@16487.4]
  wire  _T_1066; // @[MemPrimitives.scala 123:41:@16488.4]
  wire [2:0] _T_1068; // @[Cat.scala 30:58:@16490.4]
  wire [2:0] _T_1070; // @[Cat.scala 30:58:@16492.4]
  wire [2:0] _T_1072; // @[Cat.scala 30:58:@16494.4]
  wire [2:0] _T_1073; // @[Mux.scala 31:69:@16495.4]
  wire [2:0] _T_1074; // @[Mux.scala 31:69:@16496.4]
  wire  _T_1079; // @[MemPrimitives.scala 110:210:@16503.4]
  wire  _T_1084; // @[MemPrimitives.scala 110:210:@16506.4]
  wire  _T_1089; // @[MemPrimitives.scala 110:210:@16509.4]
  wire  _T_1093; // @[MemPrimitives.scala 123:41:@16518.4]
  wire  _T_1094; // @[MemPrimitives.scala 123:41:@16519.4]
  wire  _T_1095; // @[MemPrimitives.scala 123:41:@16520.4]
  wire [2:0] _T_1097; // @[Cat.scala 30:58:@16522.4]
  wire [2:0] _T_1099; // @[Cat.scala 30:58:@16524.4]
  wire [2:0] _T_1101; // @[Cat.scala 30:58:@16526.4]
  wire [2:0] _T_1102; // @[Mux.scala 31:69:@16527.4]
  wire [2:0] _T_1103; // @[Mux.scala 31:69:@16528.4]
  wire  _T_1108; // @[MemPrimitives.scala 110:210:@16535.4]
  wire  _T_1113; // @[MemPrimitives.scala 110:210:@16538.4]
  wire  _T_1118; // @[MemPrimitives.scala 110:210:@16541.4]
  wire  _T_1122; // @[MemPrimitives.scala 123:41:@16550.4]
  wire  _T_1123; // @[MemPrimitives.scala 123:41:@16551.4]
  wire  _T_1124; // @[MemPrimitives.scala 123:41:@16552.4]
  wire [2:0] _T_1126; // @[Cat.scala 30:58:@16554.4]
  wire [2:0] _T_1128; // @[Cat.scala 30:58:@16556.4]
  wire [2:0] _T_1130; // @[Cat.scala 30:58:@16558.4]
  wire [2:0] _T_1131; // @[Mux.scala 31:69:@16559.4]
  wire [2:0] _T_1132; // @[Mux.scala 31:69:@16560.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:210:@16567.4]
  wire  _T_1142; // @[MemPrimitives.scala 110:210:@16570.4]
  wire  _T_1147; // @[MemPrimitives.scala 110:210:@16573.4]
  wire  _T_1152; // @[MemPrimitives.scala 110:210:@16576.4]
  wire  _T_1157; // @[MemPrimitives.scala 110:210:@16579.4]
  wire  _T_1162; // @[MemPrimitives.scala 110:210:@16582.4]
  wire  _T_1166; // @[MemPrimitives.scala 123:41:@16594.4]
  wire  _T_1167; // @[MemPrimitives.scala 123:41:@16595.4]
  wire  _T_1168; // @[MemPrimitives.scala 123:41:@16596.4]
  wire  _T_1169; // @[MemPrimitives.scala 123:41:@16597.4]
  wire  _T_1170; // @[MemPrimitives.scala 123:41:@16598.4]
  wire  _T_1171; // @[MemPrimitives.scala 123:41:@16599.4]
  wire [2:0] _T_1173; // @[Cat.scala 30:58:@16601.4]
  wire [2:0] _T_1175; // @[Cat.scala 30:58:@16603.4]
  wire [2:0] _T_1177; // @[Cat.scala 30:58:@16605.4]
  wire [2:0] _T_1179; // @[Cat.scala 30:58:@16607.4]
  wire [2:0] _T_1181; // @[Cat.scala 30:58:@16609.4]
  wire [2:0] _T_1183; // @[Cat.scala 30:58:@16611.4]
  wire [2:0] _T_1184; // @[Mux.scala 31:69:@16612.4]
  wire [2:0] _T_1185; // @[Mux.scala 31:69:@16613.4]
  wire [2:0] _T_1186; // @[Mux.scala 31:69:@16614.4]
  wire [2:0] _T_1187; // @[Mux.scala 31:69:@16615.4]
  wire [2:0] _T_1188; // @[Mux.scala 31:69:@16616.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:210:@16623.4]
  wire  _T_1198; // @[MemPrimitives.scala 110:210:@16626.4]
  wire  _T_1203; // @[MemPrimitives.scala 110:210:@16629.4]
  wire  _T_1207; // @[MemPrimitives.scala 123:41:@16638.4]
  wire  _T_1208; // @[MemPrimitives.scala 123:41:@16639.4]
  wire  _T_1209; // @[MemPrimitives.scala 123:41:@16640.4]
  wire [2:0] _T_1211; // @[Cat.scala 30:58:@16642.4]
  wire [2:0] _T_1213; // @[Cat.scala 30:58:@16644.4]
  wire [2:0] _T_1215; // @[Cat.scala 30:58:@16646.4]
  wire [2:0] _T_1216; // @[Mux.scala 31:69:@16647.4]
  wire [2:0] _T_1217; // @[Mux.scala 31:69:@16648.4]
  wire  _T_1222; // @[MemPrimitives.scala 110:210:@16655.4]
  wire  _T_1227; // @[MemPrimitives.scala 110:210:@16658.4]
  wire  _T_1232; // @[MemPrimitives.scala 110:210:@16661.4]
  wire  _T_1236; // @[MemPrimitives.scala 123:41:@16670.4]
  wire  _T_1237; // @[MemPrimitives.scala 123:41:@16671.4]
  wire  _T_1238; // @[MemPrimitives.scala 123:41:@16672.4]
  wire [2:0] _T_1240; // @[Cat.scala 30:58:@16674.4]
  wire [2:0] _T_1242; // @[Cat.scala 30:58:@16676.4]
  wire [2:0] _T_1244; // @[Cat.scala 30:58:@16678.4]
  wire [2:0] _T_1245; // @[Mux.scala 31:69:@16679.4]
  wire [2:0] _T_1246; // @[Mux.scala 31:69:@16680.4]
  wire  _T_1251; // @[MemPrimitives.scala 110:210:@16687.4]
  wire  _T_1256; // @[MemPrimitives.scala 110:210:@16690.4]
  wire  _T_1261; // @[MemPrimitives.scala 110:210:@16693.4]
  wire  _T_1265; // @[MemPrimitives.scala 123:41:@16702.4]
  wire  _T_1266; // @[MemPrimitives.scala 123:41:@16703.4]
  wire  _T_1267; // @[MemPrimitives.scala 123:41:@16704.4]
  wire [2:0] _T_1269; // @[Cat.scala 30:58:@16706.4]
  wire [2:0] _T_1271; // @[Cat.scala 30:58:@16708.4]
  wire [2:0] _T_1273; // @[Cat.scala 30:58:@16710.4]
  wire [2:0] _T_1274; // @[Mux.scala 31:69:@16711.4]
  wire [2:0] _T_1275; // @[Mux.scala 31:69:@16712.4]
  wire  _T_1280; // @[MemPrimitives.scala 110:210:@16719.4]
  wire  _T_1285; // @[MemPrimitives.scala 110:210:@16722.4]
  wire  _T_1290; // @[MemPrimitives.scala 110:210:@16725.4]
  wire  _T_1295; // @[MemPrimitives.scala 110:210:@16728.4]
  wire  _T_1300; // @[MemPrimitives.scala 110:210:@16731.4]
  wire  _T_1305; // @[MemPrimitives.scala 110:210:@16734.4]
  wire  _T_1309; // @[MemPrimitives.scala 123:41:@16746.4]
  wire  _T_1310; // @[MemPrimitives.scala 123:41:@16747.4]
  wire  _T_1311; // @[MemPrimitives.scala 123:41:@16748.4]
  wire  _T_1312; // @[MemPrimitives.scala 123:41:@16749.4]
  wire  _T_1313; // @[MemPrimitives.scala 123:41:@16750.4]
  wire  _T_1314; // @[MemPrimitives.scala 123:41:@16751.4]
  wire [2:0] _T_1316; // @[Cat.scala 30:58:@16753.4]
  wire [2:0] _T_1318; // @[Cat.scala 30:58:@16755.4]
  wire [2:0] _T_1320; // @[Cat.scala 30:58:@16757.4]
  wire [2:0] _T_1322; // @[Cat.scala 30:58:@16759.4]
  wire [2:0] _T_1324; // @[Cat.scala 30:58:@16761.4]
  wire [2:0] _T_1326; // @[Cat.scala 30:58:@16763.4]
  wire [2:0] _T_1327; // @[Mux.scala 31:69:@16764.4]
  wire [2:0] _T_1328; // @[Mux.scala 31:69:@16765.4]
  wire [2:0] _T_1329; // @[Mux.scala 31:69:@16766.4]
  wire [2:0] _T_1330; // @[Mux.scala 31:69:@16767.4]
  wire [2:0] _T_1331; // @[Mux.scala 31:69:@16768.4]
  wire  _T_1336; // @[MemPrimitives.scala 110:210:@16775.4]
  wire  _T_1341; // @[MemPrimitives.scala 110:210:@16778.4]
  wire  _T_1346; // @[MemPrimitives.scala 110:210:@16781.4]
  wire  _T_1350; // @[MemPrimitives.scala 123:41:@16790.4]
  wire  _T_1351; // @[MemPrimitives.scala 123:41:@16791.4]
  wire  _T_1352; // @[MemPrimitives.scala 123:41:@16792.4]
  wire [2:0] _T_1354; // @[Cat.scala 30:58:@16794.4]
  wire [2:0] _T_1356; // @[Cat.scala 30:58:@16796.4]
  wire [2:0] _T_1358; // @[Cat.scala 30:58:@16798.4]
  wire [2:0] _T_1359; // @[Mux.scala 31:69:@16799.4]
  wire [2:0] _T_1360; // @[Mux.scala 31:69:@16800.4]
  wire  _T_1365; // @[MemPrimitives.scala 110:210:@16807.4]
  wire  _T_1370; // @[MemPrimitives.scala 110:210:@16810.4]
  wire  _T_1375; // @[MemPrimitives.scala 110:210:@16813.4]
  wire  _T_1379; // @[MemPrimitives.scala 123:41:@16822.4]
  wire  _T_1380; // @[MemPrimitives.scala 123:41:@16823.4]
  wire  _T_1381; // @[MemPrimitives.scala 123:41:@16824.4]
  wire [2:0] _T_1383; // @[Cat.scala 30:58:@16826.4]
  wire [2:0] _T_1385; // @[Cat.scala 30:58:@16828.4]
  wire [2:0] _T_1387; // @[Cat.scala 30:58:@16830.4]
  wire [2:0] _T_1388; // @[Mux.scala 31:69:@16831.4]
  wire [2:0] _T_1389; // @[Mux.scala 31:69:@16832.4]
  wire  _T_1394; // @[MemPrimitives.scala 110:210:@16839.4]
  wire  _T_1399; // @[MemPrimitives.scala 110:210:@16842.4]
  wire  _T_1404; // @[MemPrimitives.scala 110:210:@16845.4]
  wire  _T_1408; // @[MemPrimitives.scala 123:41:@16854.4]
  wire  _T_1409; // @[MemPrimitives.scala 123:41:@16855.4]
  wire  _T_1410; // @[MemPrimitives.scala 123:41:@16856.4]
  wire [2:0] _T_1412; // @[Cat.scala 30:58:@16858.4]
  wire [2:0] _T_1414; // @[Cat.scala 30:58:@16860.4]
  wire [2:0] _T_1416; // @[Cat.scala 30:58:@16862.4]
  wire [2:0] _T_1417; // @[Mux.scala 31:69:@16863.4]
  wire [2:0] _T_1418; // @[Mux.scala 31:69:@16864.4]
  wire  _T_1423; // @[MemPrimitives.scala 110:210:@16871.4]
  wire  _T_1428; // @[MemPrimitives.scala 110:210:@16874.4]
  wire  _T_1433; // @[MemPrimitives.scala 110:210:@16877.4]
  wire  _T_1438; // @[MemPrimitives.scala 110:210:@16880.4]
  wire  _T_1443; // @[MemPrimitives.scala 110:210:@16883.4]
  wire  _T_1448; // @[MemPrimitives.scala 110:210:@16886.4]
  wire  _T_1452; // @[MemPrimitives.scala 123:41:@16898.4]
  wire  _T_1453; // @[MemPrimitives.scala 123:41:@16899.4]
  wire  _T_1454; // @[MemPrimitives.scala 123:41:@16900.4]
  wire  _T_1455; // @[MemPrimitives.scala 123:41:@16901.4]
  wire  _T_1456; // @[MemPrimitives.scala 123:41:@16902.4]
  wire  _T_1457; // @[MemPrimitives.scala 123:41:@16903.4]
  wire [2:0] _T_1459; // @[Cat.scala 30:58:@16905.4]
  wire [2:0] _T_1461; // @[Cat.scala 30:58:@16907.4]
  wire [2:0] _T_1463; // @[Cat.scala 30:58:@16909.4]
  wire [2:0] _T_1465; // @[Cat.scala 30:58:@16911.4]
  wire [2:0] _T_1467; // @[Cat.scala 30:58:@16913.4]
  wire [2:0] _T_1469; // @[Cat.scala 30:58:@16915.4]
  wire [2:0] _T_1470; // @[Mux.scala 31:69:@16916.4]
  wire [2:0] _T_1471; // @[Mux.scala 31:69:@16917.4]
  wire [2:0] _T_1472; // @[Mux.scala 31:69:@16918.4]
  wire [2:0] _T_1473; // @[Mux.scala 31:69:@16919.4]
  wire [2:0] _T_1474; // @[Mux.scala 31:69:@16920.4]
  wire  _T_1479; // @[MemPrimitives.scala 110:210:@16927.4]
  wire  _T_1484; // @[MemPrimitives.scala 110:210:@16930.4]
  wire  _T_1489; // @[MemPrimitives.scala 110:210:@16933.4]
  wire  _T_1493; // @[MemPrimitives.scala 123:41:@16942.4]
  wire  _T_1494; // @[MemPrimitives.scala 123:41:@16943.4]
  wire  _T_1495; // @[MemPrimitives.scala 123:41:@16944.4]
  wire [2:0] _T_1497; // @[Cat.scala 30:58:@16946.4]
  wire [2:0] _T_1499; // @[Cat.scala 30:58:@16948.4]
  wire [2:0] _T_1501; // @[Cat.scala 30:58:@16950.4]
  wire [2:0] _T_1502; // @[Mux.scala 31:69:@16951.4]
  wire [2:0] _T_1503; // @[Mux.scala 31:69:@16952.4]
  wire  _T_1508; // @[MemPrimitives.scala 110:210:@16959.4]
  wire  _T_1513; // @[MemPrimitives.scala 110:210:@16962.4]
  wire  _T_1518; // @[MemPrimitives.scala 110:210:@16965.4]
  wire  _T_1522; // @[MemPrimitives.scala 123:41:@16974.4]
  wire  _T_1523; // @[MemPrimitives.scala 123:41:@16975.4]
  wire  _T_1524; // @[MemPrimitives.scala 123:41:@16976.4]
  wire [2:0] _T_1526; // @[Cat.scala 30:58:@16978.4]
  wire [2:0] _T_1528; // @[Cat.scala 30:58:@16980.4]
  wire [2:0] _T_1530; // @[Cat.scala 30:58:@16982.4]
  wire [2:0] _T_1531; // @[Mux.scala 31:69:@16983.4]
  wire [2:0] _T_1532; // @[Mux.scala 31:69:@16984.4]
  wire  _T_1537; // @[MemPrimitives.scala 110:210:@16991.4]
  wire  _T_1542; // @[MemPrimitives.scala 110:210:@16994.4]
  wire  _T_1547; // @[MemPrimitives.scala 110:210:@16997.4]
  wire  _T_1551; // @[MemPrimitives.scala 123:41:@17006.4]
  wire  _T_1552; // @[MemPrimitives.scala 123:41:@17007.4]
  wire  _T_1553; // @[MemPrimitives.scala 123:41:@17008.4]
  wire [2:0] _T_1555; // @[Cat.scala 30:58:@17010.4]
  wire [2:0] _T_1557; // @[Cat.scala 30:58:@17012.4]
  wire [2:0] _T_1559; // @[Cat.scala 30:58:@17014.4]
  wire [2:0] _T_1560; // @[Mux.scala 31:69:@17015.4]
  wire [2:0] _T_1561; // @[Mux.scala 31:69:@17016.4]
  wire  _T_1566; // @[MemPrimitives.scala 110:210:@17023.4]
  wire  _T_1571; // @[MemPrimitives.scala 110:210:@17026.4]
  wire  _T_1576; // @[MemPrimitives.scala 110:210:@17029.4]
  wire  _T_1581; // @[MemPrimitives.scala 110:210:@17032.4]
  wire  _T_1586; // @[MemPrimitives.scala 110:210:@17035.4]
  wire  _T_1591; // @[MemPrimitives.scala 110:210:@17038.4]
  wire  _T_1595; // @[MemPrimitives.scala 123:41:@17050.4]
  wire  _T_1596; // @[MemPrimitives.scala 123:41:@17051.4]
  wire  _T_1597; // @[MemPrimitives.scala 123:41:@17052.4]
  wire  _T_1598; // @[MemPrimitives.scala 123:41:@17053.4]
  wire  _T_1599; // @[MemPrimitives.scala 123:41:@17054.4]
  wire  _T_1600; // @[MemPrimitives.scala 123:41:@17055.4]
  wire [2:0] _T_1602; // @[Cat.scala 30:58:@17057.4]
  wire [2:0] _T_1604; // @[Cat.scala 30:58:@17059.4]
  wire [2:0] _T_1606; // @[Cat.scala 30:58:@17061.4]
  wire [2:0] _T_1608; // @[Cat.scala 30:58:@17063.4]
  wire [2:0] _T_1610; // @[Cat.scala 30:58:@17065.4]
  wire [2:0] _T_1612; // @[Cat.scala 30:58:@17067.4]
  wire [2:0] _T_1613; // @[Mux.scala 31:69:@17068.4]
  wire [2:0] _T_1614; // @[Mux.scala 31:69:@17069.4]
  wire [2:0] _T_1615; // @[Mux.scala 31:69:@17070.4]
  wire [2:0] _T_1616; // @[Mux.scala 31:69:@17071.4]
  wire [2:0] _T_1617; // @[Mux.scala 31:69:@17072.4]
  wire  _T_1649; // @[package.scala 96:25:@17113.4 package.scala 96:25:@17114.4]
  wire [7:0] _T_1653; // @[Mux.scala 31:69:@17123.4]
  wire  _T_1646; // @[package.scala 96:25:@17105.4 package.scala 96:25:@17106.4]
  wire [7:0] _T_1654; // @[Mux.scala 31:69:@17124.4]
  wire  _T_1643; // @[package.scala 96:25:@17097.4 package.scala 96:25:@17098.4]
  wire  _T_1684; // @[package.scala 96:25:@17161.4 package.scala 96:25:@17162.4]
  wire [7:0] _T_1688; // @[Mux.scala 31:69:@17171.4]
  wire  _T_1681; // @[package.scala 96:25:@17153.4 package.scala 96:25:@17154.4]
  wire [7:0] _T_1689; // @[Mux.scala 31:69:@17172.4]
  wire  _T_1678; // @[package.scala 96:25:@17145.4 package.scala 96:25:@17146.4]
  wire  _T_1719; // @[package.scala 96:25:@17209.4 package.scala 96:25:@17210.4]
  wire [7:0] _T_1723; // @[Mux.scala 31:69:@17219.4]
  wire  _T_1716; // @[package.scala 96:25:@17201.4 package.scala 96:25:@17202.4]
  wire [7:0] _T_1724; // @[Mux.scala 31:69:@17220.4]
  wire  _T_1713; // @[package.scala 96:25:@17193.4 package.scala 96:25:@17194.4]
  wire  _T_1754; // @[package.scala 96:25:@17257.4 package.scala 96:25:@17258.4]
  wire [7:0] _T_1758; // @[Mux.scala 31:69:@17267.4]
  wire  _T_1751; // @[package.scala 96:25:@17249.4 package.scala 96:25:@17250.4]
  wire [7:0] _T_1759; // @[Mux.scala 31:69:@17268.4]
  wire  _T_1748; // @[package.scala 96:25:@17241.4 package.scala 96:25:@17242.4]
  wire  _T_1789; // @[package.scala 96:25:@17305.4 package.scala 96:25:@17306.4]
  wire [7:0] _T_1793; // @[Mux.scala 31:69:@17315.4]
  wire  _T_1786; // @[package.scala 96:25:@17297.4 package.scala 96:25:@17298.4]
  wire [7:0] _T_1794; // @[Mux.scala 31:69:@17316.4]
  wire  _T_1783; // @[package.scala 96:25:@17289.4 package.scala 96:25:@17290.4]
  wire  _T_1824; // @[package.scala 96:25:@17353.4 package.scala 96:25:@17354.4]
  wire [7:0] _T_1828; // @[Mux.scala 31:69:@17363.4]
  wire  _T_1821; // @[package.scala 96:25:@17345.4 package.scala 96:25:@17346.4]
  wire [7:0] _T_1829; // @[Mux.scala 31:69:@17364.4]
  wire  _T_1818; // @[package.scala 96:25:@17337.4 package.scala 96:25:@17338.4]
  wire  _T_1859; // @[package.scala 96:25:@17401.4 package.scala 96:25:@17402.4]
  wire [7:0] _T_1863; // @[Mux.scala 31:69:@17411.4]
  wire  _T_1856; // @[package.scala 96:25:@17393.4 package.scala 96:25:@17394.4]
  wire [7:0] _T_1864; // @[Mux.scala 31:69:@17412.4]
  wire  _T_1853; // @[package.scala 96:25:@17385.4 package.scala 96:25:@17386.4]
  wire  _T_1894; // @[package.scala 96:25:@17449.4 package.scala 96:25:@17450.4]
  wire [7:0] _T_1898; // @[Mux.scala 31:69:@17459.4]
  wire  _T_1891; // @[package.scala 96:25:@17441.4 package.scala 96:25:@17442.4]
  wire [7:0] _T_1899; // @[Mux.scala 31:69:@17460.4]
  wire  _T_1888; // @[package.scala 96:25:@17433.4 package.scala 96:25:@17434.4]
  wire  _T_1929; // @[package.scala 96:25:@17497.4 package.scala 96:25:@17498.4]
  wire [7:0] _T_1933; // @[Mux.scala 31:69:@17507.4]
  wire  _T_1926; // @[package.scala 96:25:@17489.4 package.scala 96:25:@17490.4]
  wire [7:0] _T_1934; // @[Mux.scala 31:69:@17508.4]
  wire  _T_1923; // @[package.scala 96:25:@17481.4 package.scala 96:25:@17482.4]
  wire  _T_1964; // @[package.scala 96:25:@17545.4 package.scala 96:25:@17546.4]
  wire [7:0] _T_1968; // @[Mux.scala 31:69:@17555.4]
  wire  _T_1961; // @[package.scala 96:25:@17537.4 package.scala 96:25:@17538.4]
  wire [7:0] _T_1969; // @[Mux.scala 31:69:@17556.4]
  wire  _T_1958; // @[package.scala 96:25:@17529.4 package.scala 96:25:@17530.4]
  wire  _T_1999; // @[package.scala 96:25:@17593.4 package.scala 96:25:@17594.4]
  wire [7:0] _T_2003; // @[Mux.scala 31:69:@17603.4]
  wire  _T_1996; // @[package.scala 96:25:@17585.4 package.scala 96:25:@17586.4]
  wire [7:0] _T_2004; // @[Mux.scala 31:69:@17604.4]
  wire  _T_1993; // @[package.scala 96:25:@17577.4 package.scala 96:25:@17578.4]
  wire  _T_2034; // @[package.scala 96:25:@17641.4 package.scala 96:25:@17642.4]
  wire [7:0] _T_2038; // @[Mux.scala 31:69:@17651.4]
  wire  _T_2031; // @[package.scala 96:25:@17633.4 package.scala 96:25:@17634.4]
  wire [7:0] _T_2039; // @[Mux.scala 31:69:@17652.4]
  wire  _T_2028; // @[package.scala 96:25:@17625.4 package.scala 96:25:@17626.4]
  wire  _T_2069; // @[package.scala 96:25:@17689.4 package.scala 96:25:@17690.4]
  wire [7:0] _T_2073; // @[Mux.scala 31:69:@17699.4]
  wire  _T_2066; // @[package.scala 96:25:@17681.4 package.scala 96:25:@17682.4]
  wire [7:0] _T_2074; // @[Mux.scala 31:69:@17700.4]
  wire  _T_2063; // @[package.scala 96:25:@17673.4 package.scala 96:25:@17674.4]
  wire  _T_2104; // @[package.scala 96:25:@17737.4 package.scala 96:25:@17738.4]
  wire [7:0] _T_2108; // @[Mux.scala 31:69:@17747.4]
  wire  _T_2101; // @[package.scala 96:25:@17729.4 package.scala 96:25:@17730.4]
  wire [7:0] _T_2109; // @[Mux.scala 31:69:@17748.4]
  wire  _T_2098; // @[package.scala 96:25:@17721.4 package.scala 96:25:@17722.4]
  wire  _T_2139; // @[package.scala 96:25:@17785.4 package.scala 96:25:@17786.4]
  wire [7:0] _T_2143; // @[Mux.scala 31:69:@17795.4]
  wire  _T_2136; // @[package.scala 96:25:@17777.4 package.scala 96:25:@17778.4]
  wire [7:0] _T_2144; // @[Mux.scala 31:69:@17796.4]
  wire  _T_2133; // @[package.scala 96:25:@17769.4 package.scala 96:25:@17770.4]
  Mem1D_4 Mem1D ( // @[MemPrimitives.scala 64:21:@15943.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_4 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@15959.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_4 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@15975.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_4 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@15991.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_4 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@16007.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_4 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@16023.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_4 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@16039.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_4 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@16055.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_4 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@16071.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_4 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@16087.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_4 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@16103.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_4 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@16119.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_4 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@16135.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_4 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@16151.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_4 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@16167.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_4 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@16183.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects_16 StickySelects ( // @[MemPrimitives.scala 121:29:@16480.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2)
  );
  StickySelects_16 StickySelects_1 ( // @[MemPrimitives.scala 121:29:@16512.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2)
  );
  StickySelects_16 StickySelects_2 ( // @[MemPrimitives.scala 121:29:@16544.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2)
  );
  StickySelects_19 StickySelects_3 ( // @[MemPrimitives.scala 121:29:@16585.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5)
  );
  StickySelects_16 StickySelects_4 ( // @[MemPrimitives.scala 121:29:@16632.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2)
  );
  StickySelects_16 StickySelects_5 ( // @[MemPrimitives.scala 121:29:@16664.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2)
  );
  StickySelects_16 StickySelects_6 ( // @[MemPrimitives.scala 121:29:@16696.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2)
  );
  StickySelects_19 StickySelects_7 ( // @[MemPrimitives.scala 121:29:@16737.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5)
  );
  StickySelects_16 StickySelects_8 ( // @[MemPrimitives.scala 121:29:@16784.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2)
  );
  StickySelects_16 StickySelects_9 ( // @[MemPrimitives.scala 121:29:@16816.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2)
  );
  StickySelects_16 StickySelects_10 ( // @[MemPrimitives.scala 121:29:@16848.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2)
  );
  StickySelects_19 StickySelects_11 ( // @[MemPrimitives.scala 121:29:@16889.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5)
  );
  StickySelects_16 StickySelects_12 ( // @[MemPrimitives.scala 121:29:@16936.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2)
  );
  StickySelects_16 StickySelects_13 ( // @[MemPrimitives.scala 121:29:@16968.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2)
  );
  StickySelects_16 StickySelects_14 ( // @[MemPrimitives.scala 121:29:@17000.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2)
  );
  StickySelects_19 StickySelects_15 ( // @[MemPrimitives.scala 121:29:@17041.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@17092.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_1 ( // @[package.scala 93:22:@17100.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_2 ( // @[package.scala 93:22:@17108.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_3 ( // @[package.scala 93:22:@17116.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_4 ( // @[package.scala 93:22:@17140.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_5 ( // @[package.scala 93:22:@17148.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_6 ( // @[package.scala 93:22:@17156.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_7 ( // @[package.scala 93:22:@17164.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_8 ( // @[package.scala 93:22:@17188.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_9 ( // @[package.scala 93:22:@17196.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_10 ( // @[package.scala 93:22:@17204.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_11 ( // @[package.scala 93:22:@17212.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_12 ( // @[package.scala 93:22:@17236.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_13 ( // @[package.scala 93:22:@17244.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_14 ( // @[package.scala 93:22:@17252.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_15 ( // @[package.scala 93:22:@17260.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_16 ( // @[package.scala 93:22:@17284.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_17 ( // @[package.scala 93:22:@17292.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_18 ( // @[package.scala 93:22:@17300.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_19 ( // @[package.scala 93:22:@17308.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_20 ( // @[package.scala 93:22:@17332.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_21 ( // @[package.scala 93:22:@17340.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_22 ( // @[package.scala 93:22:@17348.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_23 ( // @[package.scala 93:22:@17356.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_24 ( // @[package.scala 93:22:@17380.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_25 ( // @[package.scala 93:22:@17388.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_26 ( // @[package.scala 93:22:@17396.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_27 ( // @[package.scala 93:22:@17404.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_28 ( // @[package.scala 93:22:@17428.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_29 ( // @[package.scala 93:22:@17436.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_30 ( // @[package.scala 93:22:@17444.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_31 ( // @[package.scala 93:22:@17452.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_32 ( // @[package.scala 93:22:@17476.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_33 ( // @[package.scala 93:22:@17484.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_34 ( // @[package.scala 93:22:@17492.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_35 ( // @[package.scala 93:22:@17500.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_36 ( // @[package.scala 93:22:@17524.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_37 ( // @[package.scala 93:22:@17532.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_38 ( // @[package.scala 93:22:@17540.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_39 ( // @[package.scala 93:22:@17548.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_40 ( // @[package.scala 93:22:@17572.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_41 ( // @[package.scala 93:22:@17580.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_42 ( // @[package.scala 93:22:@17588.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_43 ( // @[package.scala 93:22:@17596.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_44 ( // @[package.scala 93:22:@17620.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_45 ( // @[package.scala 93:22:@17628.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_46 ( // @[package.scala 93:22:@17636.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_47 ( // @[package.scala 93:22:@17644.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_48 ( // @[package.scala 93:22:@17668.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_49 ( // @[package.scala 93:22:@17676.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_50 ( // @[package.scala 93:22:@17684.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_51 ( // @[package.scala 93:22:@17692.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_52 ( // @[package.scala 93:22:@17716.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_53 ( // @[package.scala 93:22:@17724.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_54 ( // @[package.scala 93:22:@17732.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_55 ( // @[package.scala 93:22:@17740.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_56 ( // @[package.scala 93:22:@17764.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_57 ( // @[package.scala 93:22:@17772.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_58 ( // @[package.scala 93:22:@17780.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_59 ( // @[package.scala 93:22:@17788.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  assign _T_762 = io_wPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@16199.4]
  assign _T_765 = io_wPort_3_en_0 & _T_762; // @[MemPrimitives.scala 83:102:@16201.4]
  assign _T_767 = io_wPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@16202.4]
  assign _T_770 = io_wPort_5_en_0 & _T_767; // @[MemPrimitives.scala 83:102:@16204.4]
  assign _T_772 = {_T_765,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16206.4]
  assign _T_774 = {_T_770,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@16208.4]
  assign _T_775 = _T_765 ? _T_772 : _T_774; // @[Mux.scala 31:69:@16209.4]
  assign _T_780 = io_wPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@16216.4]
  assign _T_783 = io_wPort_4_en_0 & _T_780; // @[MemPrimitives.scala 83:102:@16218.4]
  assign _T_785 = io_wPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@16219.4]
  assign _T_788 = io_wPort_7_en_0 & _T_785; // @[MemPrimitives.scala 83:102:@16221.4]
  assign _T_790 = {_T_783,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@16223.4]
  assign _T_792 = {_T_788,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@16225.4]
  assign _T_793 = _T_783 ? _T_790 : _T_792; // @[Mux.scala 31:69:@16226.4]
  assign _T_798 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@16233.4]
  assign _T_801 = io_wPort_0_en_0 & _T_798; // @[MemPrimitives.scala 83:102:@16235.4]
  assign _T_803 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@16236.4]
  assign _T_806 = io_wPort_1_en_0 & _T_803; // @[MemPrimitives.scala 83:102:@16238.4]
  assign _T_808 = {_T_801,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16240.4]
  assign _T_810 = {_T_806,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16242.4]
  assign _T_811 = _T_801 ? _T_808 : _T_810; // @[Mux.scala 31:69:@16243.4]
  assign _T_816 = io_wPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@16250.4]
  assign _T_819 = io_wPort_2_en_0 & _T_816; // @[MemPrimitives.scala 83:102:@16252.4]
  assign _T_821 = io_wPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@16253.4]
  assign _T_824 = io_wPort_6_en_0 & _T_821; // @[MemPrimitives.scala 83:102:@16255.4]
  assign _T_826 = {_T_819,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16257.4]
  assign _T_828 = {_T_824,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@16259.4]
  assign _T_829 = _T_819 ? _T_826 : _T_828; // @[Mux.scala 31:69:@16260.4]
  assign _T_834 = io_wPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@16267.4]
  assign _T_837 = io_wPort_3_en_0 & _T_834; // @[MemPrimitives.scala 83:102:@16269.4]
  assign _T_839 = io_wPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@16270.4]
  assign _T_842 = io_wPort_5_en_0 & _T_839; // @[MemPrimitives.scala 83:102:@16272.4]
  assign _T_844 = {_T_837,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16274.4]
  assign _T_846 = {_T_842,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@16276.4]
  assign _T_847 = _T_837 ? _T_844 : _T_846; // @[Mux.scala 31:69:@16277.4]
  assign _T_852 = io_wPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@16284.4]
  assign _T_855 = io_wPort_4_en_0 & _T_852; // @[MemPrimitives.scala 83:102:@16286.4]
  assign _T_857 = io_wPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@16287.4]
  assign _T_860 = io_wPort_7_en_0 & _T_857; // @[MemPrimitives.scala 83:102:@16289.4]
  assign _T_862 = {_T_855,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@16291.4]
  assign _T_864 = {_T_860,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@16293.4]
  assign _T_865 = _T_855 ? _T_862 : _T_864; // @[Mux.scala 31:69:@16294.4]
  assign _T_870 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@16301.4]
  assign _T_873 = io_wPort_0_en_0 & _T_870; // @[MemPrimitives.scala 83:102:@16303.4]
  assign _T_875 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@16304.4]
  assign _T_878 = io_wPort_1_en_0 & _T_875; // @[MemPrimitives.scala 83:102:@16306.4]
  assign _T_880 = {_T_873,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16308.4]
  assign _T_882 = {_T_878,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16310.4]
  assign _T_883 = _T_873 ? _T_880 : _T_882; // @[Mux.scala 31:69:@16311.4]
  assign _T_888 = io_wPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@16318.4]
  assign _T_891 = io_wPort_2_en_0 & _T_888; // @[MemPrimitives.scala 83:102:@16320.4]
  assign _T_893 = io_wPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@16321.4]
  assign _T_896 = io_wPort_6_en_0 & _T_893; // @[MemPrimitives.scala 83:102:@16323.4]
  assign _T_898 = {_T_891,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16325.4]
  assign _T_900 = {_T_896,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@16327.4]
  assign _T_901 = _T_891 ? _T_898 : _T_900; // @[Mux.scala 31:69:@16328.4]
  assign _T_906 = io_wPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@16335.4]
  assign _T_909 = io_wPort_3_en_0 & _T_906; // @[MemPrimitives.scala 83:102:@16337.4]
  assign _T_911 = io_wPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@16338.4]
  assign _T_914 = io_wPort_5_en_0 & _T_911; // @[MemPrimitives.scala 83:102:@16340.4]
  assign _T_916 = {_T_909,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16342.4]
  assign _T_918 = {_T_914,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@16344.4]
  assign _T_919 = _T_909 ? _T_916 : _T_918; // @[Mux.scala 31:69:@16345.4]
  assign _T_924 = io_wPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@16352.4]
  assign _T_927 = io_wPort_4_en_0 & _T_924; // @[MemPrimitives.scala 83:102:@16354.4]
  assign _T_929 = io_wPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@16355.4]
  assign _T_932 = io_wPort_7_en_0 & _T_929; // @[MemPrimitives.scala 83:102:@16357.4]
  assign _T_934 = {_T_927,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@16359.4]
  assign _T_936 = {_T_932,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@16361.4]
  assign _T_937 = _T_927 ? _T_934 : _T_936; // @[Mux.scala 31:69:@16362.4]
  assign _T_942 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@16369.4]
  assign _T_945 = io_wPort_0_en_0 & _T_942; // @[MemPrimitives.scala 83:102:@16371.4]
  assign _T_947 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@16372.4]
  assign _T_950 = io_wPort_1_en_0 & _T_947; // @[MemPrimitives.scala 83:102:@16374.4]
  assign _T_952 = {_T_945,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16376.4]
  assign _T_954 = {_T_950,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16378.4]
  assign _T_955 = _T_945 ? _T_952 : _T_954; // @[Mux.scala 31:69:@16379.4]
  assign _T_960 = io_wPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@16386.4]
  assign _T_963 = io_wPort_2_en_0 & _T_960; // @[MemPrimitives.scala 83:102:@16388.4]
  assign _T_965 = io_wPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@16389.4]
  assign _T_968 = io_wPort_6_en_0 & _T_965; // @[MemPrimitives.scala 83:102:@16391.4]
  assign _T_970 = {_T_963,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16393.4]
  assign _T_972 = {_T_968,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@16395.4]
  assign _T_973 = _T_963 ? _T_970 : _T_972; // @[Mux.scala 31:69:@16396.4]
  assign _T_978 = io_wPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@16403.4]
  assign _T_981 = io_wPort_3_en_0 & _T_978; // @[MemPrimitives.scala 83:102:@16405.4]
  assign _T_983 = io_wPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@16406.4]
  assign _T_986 = io_wPort_5_en_0 & _T_983; // @[MemPrimitives.scala 83:102:@16408.4]
  assign _T_988 = {_T_981,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@16410.4]
  assign _T_990 = {_T_986,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@16412.4]
  assign _T_991 = _T_981 ? _T_988 : _T_990; // @[Mux.scala 31:69:@16413.4]
  assign _T_996 = io_wPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@16420.4]
  assign _T_999 = io_wPort_4_en_0 & _T_996; // @[MemPrimitives.scala 83:102:@16422.4]
  assign _T_1001 = io_wPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@16423.4]
  assign _T_1004 = io_wPort_7_en_0 & _T_1001; // @[MemPrimitives.scala 83:102:@16425.4]
  assign _T_1006 = {_T_999,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@16427.4]
  assign _T_1008 = {_T_1004,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@16429.4]
  assign _T_1009 = _T_999 ? _T_1006 : _T_1008; // @[Mux.scala 31:69:@16430.4]
  assign _T_1014 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@16437.4]
  assign _T_1017 = io_wPort_0_en_0 & _T_1014; // @[MemPrimitives.scala 83:102:@16439.4]
  assign _T_1019 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@16440.4]
  assign _T_1022 = io_wPort_1_en_0 & _T_1019; // @[MemPrimitives.scala 83:102:@16442.4]
  assign _T_1024 = {_T_1017,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@16444.4]
  assign _T_1026 = {_T_1022,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@16446.4]
  assign _T_1027 = _T_1017 ? _T_1024 : _T_1026; // @[Mux.scala 31:69:@16447.4]
  assign _T_1032 = io_wPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@16454.4]
  assign _T_1035 = io_wPort_2_en_0 & _T_1032; // @[MemPrimitives.scala 83:102:@16456.4]
  assign _T_1037 = io_wPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@16457.4]
  assign _T_1040 = io_wPort_6_en_0 & _T_1037; // @[MemPrimitives.scala 83:102:@16459.4]
  assign _T_1042 = {_T_1035,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@16461.4]
  assign _T_1044 = {_T_1040,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@16463.4]
  assign _T_1045 = _T_1035 ? _T_1042 : _T_1044; // @[Mux.scala 31:69:@16464.4]
  assign _T_1050 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16471.4]
  assign _T_1055 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16474.4]
  assign _T_1060 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16477.4]
  assign _T_1064 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@16486.4]
  assign _T_1065 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@16487.4]
  assign _T_1066 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@16488.4]
  assign _T_1068 = {_T_1064,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@16490.4]
  assign _T_1070 = {_T_1065,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@16492.4]
  assign _T_1072 = {_T_1066,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@16494.4]
  assign _T_1073 = _T_1065 ? _T_1070 : _T_1072; // @[Mux.scala 31:69:@16495.4]
  assign _T_1074 = _T_1064 ? _T_1068 : _T_1073; // @[Mux.scala 31:69:@16496.4]
  assign _T_1079 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16503.4]
  assign _T_1084 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16506.4]
  assign _T_1089 = io_rPort_14_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16509.4]
  assign _T_1093 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@16518.4]
  assign _T_1094 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@16519.4]
  assign _T_1095 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@16520.4]
  assign _T_1097 = {_T_1093,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@16522.4]
  assign _T_1099 = {_T_1094,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@16524.4]
  assign _T_1101 = {_T_1095,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@16526.4]
  assign _T_1102 = _T_1094 ? _T_1099 : _T_1101; // @[Mux.scala 31:69:@16527.4]
  assign _T_1103 = _T_1093 ? _T_1097 : _T_1102; // @[Mux.scala 31:69:@16528.4]
  assign _T_1108 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16535.4]
  assign _T_1113 = io_rPort_12_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16538.4]
  assign _T_1118 = io_rPort_13_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16541.4]
  assign _T_1122 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@16550.4]
  assign _T_1123 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@16551.4]
  assign _T_1124 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@16552.4]
  assign _T_1126 = {_T_1122,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@16554.4]
  assign _T_1128 = {_T_1123,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@16556.4]
  assign _T_1130 = {_T_1124,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@16558.4]
  assign _T_1131 = _T_1123 ? _T_1128 : _T_1130; // @[Mux.scala 31:69:@16559.4]
  assign _T_1132 = _T_1122 ? _T_1126 : _T_1131; // @[Mux.scala 31:69:@16560.4]
  assign _T_1137 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16567.4]
  assign _T_1142 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16570.4]
  assign _T_1147 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16573.4]
  assign _T_1152 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16576.4]
  assign _T_1157 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16579.4]
  assign _T_1162 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@16582.4]
  assign _T_1166 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@16594.4]
  assign _T_1167 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@16595.4]
  assign _T_1168 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@16596.4]
  assign _T_1169 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@16597.4]
  assign _T_1170 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@16598.4]
  assign _T_1171 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@16599.4]
  assign _T_1173 = {_T_1166,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@16601.4]
  assign _T_1175 = {_T_1167,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@16603.4]
  assign _T_1177 = {_T_1168,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@16605.4]
  assign _T_1179 = {_T_1169,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@16607.4]
  assign _T_1181 = {_T_1170,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@16609.4]
  assign _T_1183 = {_T_1171,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@16611.4]
  assign _T_1184 = _T_1170 ? _T_1181 : _T_1183; // @[Mux.scala 31:69:@16612.4]
  assign _T_1185 = _T_1169 ? _T_1179 : _T_1184; // @[Mux.scala 31:69:@16613.4]
  assign _T_1186 = _T_1168 ? _T_1177 : _T_1185; // @[Mux.scala 31:69:@16614.4]
  assign _T_1187 = _T_1167 ? _T_1175 : _T_1186; // @[Mux.scala 31:69:@16615.4]
  assign _T_1188 = _T_1166 ? _T_1173 : _T_1187; // @[Mux.scala 31:69:@16616.4]
  assign _T_1193 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16623.4]
  assign _T_1198 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16626.4]
  assign _T_1203 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16629.4]
  assign _T_1207 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@16638.4]
  assign _T_1208 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@16639.4]
  assign _T_1209 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@16640.4]
  assign _T_1211 = {_T_1207,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@16642.4]
  assign _T_1213 = {_T_1208,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@16644.4]
  assign _T_1215 = {_T_1209,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@16646.4]
  assign _T_1216 = _T_1208 ? _T_1213 : _T_1215; // @[Mux.scala 31:69:@16647.4]
  assign _T_1217 = _T_1207 ? _T_1211 : _T_1216; // @[Mux.scala 31:69:@16648.4]
  assign _T_1222 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16655.4]
  assign _T_1227 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16658.4]
  assign _T_1232 = io_rPort_14_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16661.4]
  assign _T_1236 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@16670.4]
  assign _T_1237 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@16671.4]
  assign _T_1238 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@16672.4]
  assign _T_1240 = {_T_1236,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@16674.4]
  assign _T_1242 = {_T_1237,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@16676.4]
  assign _T_1244 = {_T_1238,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@16678.4]
  assign _T_1245 = _T_1237 ? _T_1242 : _T_1244; // @[Mux.scala 31:69:@16679.4]
  assign _T_1246 = _T_1236 ? _T_1240 : _T_1245; // @[Mux.scala 31:69:@16680.4]
  assign _T_1251 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16687.4]
  assign _T_1256 = io_rPort_12_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16690.4]
  assign _T_1261 = io_rPort_13_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16693.4]
  assign _T_1265 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@16702.4]
  assign _T_1266 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@16703.4]
  assign _T_1267 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@16704.4]
  assign _T_1269 = {_T_1265,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@16706.4]
  assign _T_1271 = {_T_1266,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@16708.4]
  assign _T_1273 = {_T_1267,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@16710.4]
  assign _T_1274 = _T_1266 ? _T_1271 : _T_1273; // @[Mux.scala 31:69:@16711.4]
  assign _T_1275 = _T_1265 ? _T_1269 : _T_1274; // @[Mux.scala 31:69:@16712.4]
  assign _T_1280 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16719.4]
  assign _T_1285 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16722.4]
  assign _T_1290 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16725.4]
  assign _T_1295 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16728.4]
  assign _T_1300 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16731.4]
  assign _T_1305 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@16734.4]
  assign _T_1309 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@16746.4]
  assign _T_1310 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@16747.4]
  assign _T_1311 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@16748.4]
  assign _T_1312 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@16749.4]
  assign _T_1313 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@16750.4]
  assign _T_1314 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@16751.4]
  assign _T_1316 = {_T_1309,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@16753.4]
  assign _T_1318 = {_T_1310,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@16755.4]
  assign _T_1320 = {_T_1311,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@16757.4]
  assign _T_1322 = {_T_1312,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@16759.4]
  assign _T_1324 = {_T_1313,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@16761.4]
  assign _T_1326 = {_T_1314,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@16763.4]
  assign _T_1327 = _T_1313 ? _T_1324 : _T_1326; // @[Mux.scala 31:69:@16764.4]
  assign _T_1328 = _T_1312 ? _T_1322 : _T_1327; // @[Mux.scala 31:69:@16765.4]
  assign _T_1329 = _T_1311 ? _T_1320 : _T_1328; // @[Mux.scala 31:69:@16766.4]
  assign _T_1330 = _T_1310 ? _T_1318 : _T_1329; // @[Mux.scala 31:69:@16767.4]
  assign _T_1331 = _T_1309 ? _T_1316 : _T_1330; // @[Mux.scala 31:69:@16768.4]
  assign _T_1336 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@16775.4]
  assign _T_1341 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@16778.4]
  assign _T_1346 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@16781.4]
  assign _T_1350 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@16790.4]
  assign _T_1351 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@16791.4]
  assign _T_1352 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@16792.4]
  assign _T_1354 = {_T_1350,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@16794.4]
  assign _T_1356 = {_T_1351,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@16796.4]
  assign _T_1358 = {_T_1352,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@16798.4]
  assign _T_1359 = _T_1351 ? _T_1356 : _T_1358; // @[Mux.scala 31:69:@16799.4]
  assign _T_1360 = _T_1350 ? _T_1354 : _T_1359; // @[Mux.scala 31:69:@16800.4]
  assign _T_1365 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@16807.4]
  assign _T_1370 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@16810.4]
  assign _T_1375 = io_rPort_14_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@16813.4]
  assign _T_1379 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@16822.4]
  assign _T_1380 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@16823.4]
  assign _T_1381 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@16824.4]
  assign _T_1383 = {_T_1379,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@16826.4]
  assign _T_1385 = {_T_1380,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@16828.4]
  assign _T_1387 = {_T_1381,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@16830.4]
  assign _T_1388 = _T_1380 ? _T_1385 : _T_1387; // @[Mux.scala 31:69:@16831.4]
  assign _T_1389 = _T_1379 ? _T_1383 : _T_1388; // @[Mux.scala 31:69:@16832.4]
  assign _T_1394 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@16839.4]
  assign _T_1399 = io_rPort_12_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@16842.4]
  assign _T_1404 = io_rPort_13_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@16845.4]
  assign _T_1408 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@16854.4]
  assign _T_1409 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@16855.4]
  assign _T_1410 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@16856.4]
  assign _T_1412 = {_T_1408,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@16858.4]
  assign _T_1414 = {_T_1409,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@16860.4]
  assign _T_1416 = {_T_1410,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@16862.4]
  assign _T_1417 = _T_1409 ? _T_1414 : _T_1416; // @[Mux.scala 31:69:@16863.4]
  assign _T_1418 = _T_1408 ? _T_1412 : _T_1417; // @[Mux.scala 31:69:@16864.4]
  assign _T_1423 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@16871.4]
  assign _T_1428 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@16874.4]
  assign _T_1433 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@16877.4]
  assign _T_1438 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@16880.4]
  assign _T_1443 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@16883.4]
  assign _T_1448 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@16886.4]
  assign _T_1452 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@16898.4]
  assign _T_1453 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@16899.4]
  assign _T_1454 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@16900.4]
  assign _T_1455 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@16901.4]
  assign _T_1456 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@16902.4]
  assign _T_1457 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@16903.4]
  assign _T_1459 = {_T_1452,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@16905.4]
  assign _T_1461 = {_T_1453,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@16907.4]
  assign _T_1463 = {_T_1454,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@16909.4]
  assign _T_1465 = {_T_1455,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@16911.4]
  assign _T_1467 = {_T_1456,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@16913.4]
  assign _T_1469 = {_T_1457,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@16915.4]
  assign _T_1470 = _T_1456 ? _T_1467 : _T_1469; // @[Mux.scala 31:69:@16916.4]
  assign _T_1471 = _T_1455 ? _T_1465 : _T_1470; // @[Mux.scala 31:69:@16917.4]
  assign _T_1472 = _T_1454 ? _T_1463 : _T_1471; // @[Mux.scala 31:69:@16918.4]
  assign _T_1473 = _T_1453 ? _T_1461 : _T_1472; // @[Mux.scala 31:69:@16919.4]
  assign _T_1474 = _T_1452 ? _T_1459 : _T_1473; // @[Mux.scala 31:69:@16920.4]
  assign _T_1479 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@16927.4]
  assign _T_1484 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@16930.4]
  assign _T_1489 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@16933.4]
  assign _T_1493 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@16942.4]
  assign _T_1494 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@16943.4]
  assign _T_1495 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 123:41:@16944.4]
  assign _T_1497 = {_T_1493,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@16946.4]
  assign _T_1499 = {_T_1494,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@16948.4]
  assign _T_1501 = {_T_1495,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@16950.4]
  assign _T_1502 = _T_1494 ? _T_1499 : _T_1501; // @[Mux.scala 31:69:@16951.4]
  assign _T_1503 = _T_1493 ? _T_1497 : _T_1502; // @[Mux.scala 31:69:@16952.4]
  assign _T_1508 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@16959.4]
  assign _T_1513 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@16962.4]
  assign _T_1518 = io_rPort_14_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@16965.4]
  assign _T_1522 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@16974.4]
  assign _T_1523 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@16975.4]
  assign _T_1524 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 123:41:@16976.4]
  assign _T_1526 = {_T_1522,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@16978.4]
  assign _T_1528 = {_T_1523,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@16980.4]
  assign _T_1530 = {_T_1524,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@16982.4]
  assign _T_1531 = _T_1523 ? _T_1528 : _T_1530; // @[Mux.scala 31:69:@16983.4]
  assign _T_1532 = _T_1522 ? _T_1526 : _T_1531; // @[Mux.scala 31:69:@16984.4]
  assign _T_1537 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@16991.4]
  assign _T_1542 = io_rPort_12_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@16994.4]
  assign _T_1547 = io_rPort_13_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@16997.4]
  assign _T_1551 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@17006.4]
  assign _T_1552 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@17007.4]
  assign _T_1553 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 123:41:@17008.4]
  assign _T_1555 = {_T_1551,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@17010.4]
  assign _T_1557 = {_T_1552,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@17012.4]
  assign _T_1559 = {_T_1553,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@17014.4]
  assign _T_1560 = _T_1552 ? _T_1557 : _T_1559; // @[Mux.scala 31:69:@17015.4]
  assign _T_1561 = _T_1551 ? _T_1555 : _T_1560; // @[Mux.scala 31:69:@17016.4]
  assign _T_1566 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@17023.4]
  assign _T_1571 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@17026.4]
  assign _T_1576 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@17029.4]
  assign _T_1581 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@17032.4]
  assign _T_1586 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@17035.4]
  assign _T_1591 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@17038.4]
  assign _T_1595 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@17050.4]
  assign _T_1596 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@17051.4]
  assign _T_1597 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@17052.4]
  assign _T_1598 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@17053.4]
  assign _T_1599 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 123:41:@17054.4]
  assign _T_1600 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 123:41:@17055.4]
  assign _T_1602 = {_T_1595,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@17057.4]
  assign _T_1604 = {_T_1596,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@17059.4]
  assign _T_1606 = {_T_1597,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@17061.4]
  assign _T_1608 = {_T_1598,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@17063.4]
  assign _T_1610 = {_T_1599,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@17065.4]
  assign _T_1612 = {_T_1600,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@17067.4]
  assign _T_1613 = _T_1599 ? _T_1610 : _T_1612; // @[Mux.scala 31:69:@17068.4]
  assign _T_1614 = _T_1598 ? _T_1608 : _T_1613; // @[Mux.scala 31:69:@17069.4]
  assign _T_1615 = _T_1597 ? _T_1606 : _T_1614; // @[Mux.scala 31:69:@17070.4]
  assign _T_1616 = _T_1596 ? _T_1604 : _T_1615; // @[Mux.scala 31:69:@17071.4]
  assign _T_1617 = _T_1595 ? _T_1602 : _T_1616; // @[Mux.scala 31:69:@17072.4]
  assign _T_1649 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@17113.4 package.scala 96:25:@17114.4]
  assign _T_1653 = _T_1649 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@17123.4]
  assign _T_1646 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@17105.4 package.scala 96:25:@17106.4]
  assign _T_1654 = _T_1646 ? Mem1D_5_io_output : _T_1653; // @[Mux.scala 31:69:@17124.4]
  assign _T_1643 = RetimeWrapper_io_out; // @[package.scala 96:25:@17097.4 package.scala 96:25:@17098.4]
  assign _T_1684 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@17161.4 package.scala 96:25:@17162.4]
  assign _T_1688 = _T_1684 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@17171.4]
  assign _T_1681 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@17153.4 package.scala 96:25:@17154.4]
  assign _T_1689 = _T_1681 ? Mem1D_7_io_output : _T_1688; // @[Mux.scala 31:69:@17172.4]
  assign _T_1678 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@17145.4 package.scala 96:25:@17146.4]
  assign _T_1719 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@17209.4 package.scala 96:25:@17210.4]
  assign _T_1723 = _T_1719 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@17219.4]
  assign _T_1716 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@17201.4 package.scala 96:25:@17202.4]
  assign _T_1724 = _T_1716 ? Mem1D_7_io_output : _T_1723; // @[Mux.scala 31:69:@17220.4]
  assign _T_1713 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@17193.4 package.scala 96:25:@17194.4]
  assign _T_1754 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@17257.4 package.scala 96:25:@17258.4]
  assign _T_1758 = _T_1754 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@17267.4]
  assign _T_1751 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@17249.4 package.scala 96:25:@17250.4]
  assign _T_1759 = _T_1751 ? Mem1D_5_io_output : _T_1758; // @[Mux.scala 31:69:@17268.4]
  assign _T_1748 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@17241.4 package.scala 96:25:@17242.4]
  assign _T_1789 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@17305.4 package.scala 96:25:@17306.4]
  assign _T_1793 = _T_1789 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@17315.4]
  assign _T_1786 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@17297.4 package.scala 96:25:@17298.4]
  assign _T_1794 = _T_1786 ? Mem1D_4_io_output : _T_1793; // @[Mux.scala 31:69:@17316.4]
  assign _T_1783 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@17289.4 package.scala 96:25:@17290.4]
  assign _T_1824 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@17353.4 package.scala 96:25:@17354.4]
  assign _T_1828 = _T_1824 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@17363.4]
  assign _T_1821 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@17345.4 package.scala 96:25:@17346.4]
  assign _T_1829 = _T_1821 ? Mem1D_7_io_output : _T_1828; // @[Mux.scala 31:69:@17364.4]
  assign _T_1818 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@17337.4 package.scala 96:25:@17338.4]
  assign _T_1859 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@17401.4 package.scala 96:25:@17402.4]
  assign _T_1863 = _T_1859 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@17411.4]
  assign _T_1856 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@17393.4 package.scala 96:25:@17394.4]
  assign _T_1864 = _T_1856 ? Mem1D_6_io_output : _T_1863; // @[Mux.scala 31:69:@17412.4]
  assign _T_1853 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@17385.4 package.scala 96:25:@17386.4]
  assign _T_1894 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@17449.4 package.scala 96:25:@17450.4]
  assign _T_1898 = _T_1894 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@17459.4]
  assign _T_1891 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@17441.4 package.scala 96:25:@17442.4]
  assign _T_1899 = _T_1891 ? Mem1D_7_io_output : _T_1898; // @[Mux.scala 31:69:@17460.4]
  assign _T_1888 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@17433.4 package.scala 96:25:@17434.4]
  assign _T_1929 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@17497.4 package.scala 96:25:@17498.4]
  assign _T_1933 = _T_1929 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@17507.4]
  assign _T_1926 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@17489.4 package.scala 96:25:@17490.4]
  assign _T_1934 = _T_1926 ? Mem1D_7_io_output : _T_1933; // @[Mux.scala 31:69:@17508.4]
  assign _T_1923 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@17481.4 package.scala 96:25:@17482.4]
  assign _T_1964 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@17545.4 package.scala 96:25:@17546.4]
  assign _T_1968 = _T_1964 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@17555.4]
  assign _T_1961 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@17537.4 package.scala 96:25:@17538.4]
  assign _T_1969 = _T_1961 ? Mem1D_4_io_output : _T_1968; // @[Mux.scala 31:69:@17556.4]
  assign _T_1958 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@17529.4 package.scala 96:25:@17530.4]
  assign _T_1999 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@17593.4 package.scala 96:25:@17594.4]
  assign _T_2003 = _T_1999 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@17603.4]
  assign _T_1996 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@17585.4 package.scala 96:25:@17586.4]
  assign _T_2004 = _T_1996 ? Mem1D_4_io_output : _T_2003; // @[Mux.scala 31:69:@17604.4]
  assign _T_1993 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@17577.4 package.scala 96:25:@17578.4]
  assign _T_2034 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@17641.4 package.scala 96:25:@17642.4]
  assign _T_2038 = _T_2034 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@17651.4]
  assign _T_2031 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@17633.4 package.scala 96:25:@17634.4]
  assign _T_2039 = _T_2031 ? Mem1D_7_io_output : _T_2038; // @[Mux.scala 31:69:@17652.4]
  assign _T_2028 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@17625.4 package.scala 96:25:@17626.4]
  assign _T_2069 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@17689.4 package.scala 96:25:@17690.4]
  assign _T_2073 = _T_2069 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@17699.4]
  assign _T_2066 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@17681.4 package.scala 96:25:@17682.4]
  assign _T_2074 = _T_2066 ? Mem1D_6_io_output : _T_2073; // @[Mux.scala 31:69:@17700.4]
  assign _T_2063 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@17673.4 package.scala 96:25:@17674.4]
  assign _T_2104 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@17737.4 package.scala 96:25:@17738.4]
  assign _T_2108 = _T_2104 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@17747.4]
  assign _T_2101 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@17729.4 package.scala 96:25:@17730.4]
  assign _T_2109 = _T_2101 ? Mem1D_6_io_output : _T_2108; // @[Mux.scala 31:69:@17748.4]
  assign _T_2098 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@17721.4 package.scala 96:25:@17722.4]
  assign _T_2139 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@17785.4 package.scala 96:25:@17786.4]
  assign _T_2143 = _T_2139 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@17795.4]
  assign _T_2136 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@17777.4 package.scala 96:25:@17778.4]
  assign _T_2144 = _T_2136 ? Mem1D_5_io_output : _T_2143; // @[Mux.scala 31:69:@17796.4]
  assign _T_2133 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@17769.4 package.scala 96:25:@17770.4]
  assign io_rPort_14_output_0 = _T_2133 ? Mem1D_1_io_output : _T_2144; // @[MemPrimitives.scala 148:13:@17798.4]
  assign io_rPort_13_output_0 = _T_2098 ? Mem1D_2_io_output : _T_2109; // @[MemPrimitives.scala 148:13:@17750.4]
  assign io_rPort_12_output_0 = _T_2063 ? Mem1D_2_io_output : _T_2074; // @[MemPrimitives.scala 148:13:@17702.4]
  assign io_rPort_11_output_0 = _T_2028 ? Mem1D_3_io_output : _T_2039; // @[MemPrimitives.scala 148:13:@17654.4]
  assign io_rPort_10_output_0 = _T_1993 ? Mem1D_io_output : _T_2004; // @[MemPrimitives.scala 148:13:@17606.4]
  assign io_rPort_9_output_0 = _T_1958 ? Mem1D_io_output : _T_1969; // @[MemPrimitives.scala 148:13:@17558.4]
  assign io_rPort_8_output_0 = _T_1923 ? Mem1D_3_io_output : _T_1934; // @[MemPrimitives.scala 148:13:@17510.4]
  assign io_rPort_7_output_0 = _T_1888 ? Mem1D_3_io_output : _T_1899; // @[MemPrimitives.scala 148:13:@17462.4]
  assign io_rPort_6_output_0 = _T_1853 ? Mem1D_2_io_output : _T_1864; // @[MemPrimitives.scala 148:13:@17414.4]
  assign io_rPort_5_output_0 = _T_1818 ? Mem1D_3_io_output : _T_1829; // @[MemPrimitives.scala 148:13:@17366.4]
  assign io_rPort_4_output_0 = _T_1783 ? Mem1D_io_output : _T_1794; // @[MemPrimitives.scala 148:13:@17318.4]
  assign io_rPort_3_output_0 = _T_1748 ? Mem1D_1_io_output : _T_1759; // @[MemPrimitives.scala 148:13:@17270.4]
  assign io_rPort_2_output_0 = _T_1713 ? Mem1D_3_io_output : _T_1724; // @[MemPrimitives.scala 148:13:@17222.4]
  assign io_rPort_1_output_0 = _T_1678 ? Mem1D_3_io_output : _T_1689; // @[MemPrimitives.scala 148:13:@17174.4]
  assign io_rPort_0_output_0 = _T_1643 ? Mem1D_1_io_output : _T_1654; // @[MemPrimitives.scala 148:13:@17126.4]
  assign Mem1D_clock = clock; // @[:@15944.4]
  assign Mem1D_reset = reset; // @[:@15945.4]
  assign Mem1D_io_r_ofs_0 = _T_1074[0]; // @[MemPrimitives.scala 127:28:@16500.4]
  assign Mem1D_io_r_backpressure = _T_1074[1]; // @[MemPrimitives.scala 128:32:@16501.4]
  assign Mem1D_io_w_ofs_0 = _T_775[0]; // @[MemPrimitives.scala 94:28:@16213.4]
  assign Mem1D_io_w_data_0 = _T_775[8:1]; // @[MemPrimitives.scala 95:29:@16214.4]
  assign Mem1D_io_w_en_0 = _T_775[9]; // @[MemPrimitives.scala 96:27:@16215.4]
  assign Mem1D_1_clock = clock; // @[:@15960.4]
  assign Mem1D_1_reset = reset; // @[:@15961.4]
  assign Mem1D_1_io_r_ofs_0 = _T_1103[0]; // @[MemPrimitives.scala 127:28:@16532.4]
  assign Mem1D_1_io_r_backpressure = _T_1103[1]; // @[MemPrimitives.scala 128:32:@16533.4]
  assign Mem1D_1_io_w_ofs_0 = _T_793[0]; // @[MemPrimitives.scala 94:28:@16230.4]
  assign Mem1D_1_io_w_data_0 = _T_793[8:1]; // @[MemPrimitives.scala 95:29:@16231.4]
  assign Mem1D_1_io_w_en_0 = _T_793[9]; // @[MemPrimitives.scala 96:27:@16232.4]
  assign Mem1D_2_clock = clock; // @[:@15976.4]
  assign Mem1D_2_reset = reset; // @[:@15977.4]
  assign Mem1D_2_io_r_ofs_0 = _T_1132[0]; // @[MemPrimitives.scala 127:28:@16564.4]
  assign Mem1D_2_io_r_backpressure = _T_1132[1]; // @[MemPrimitives.scala 128:32:@16565.4]
  assign Mem1D_2_io_w_ofs_0 = _T_811[0]; // @[MemPrimitives.scala 94:28:@16247.4]
  assign Mem1D_2_io_w_data_0 = _T_811[8:1]; // @[MemPrimitives.scala 95:29:@16248.4]
  assign Mem1D_2_io_w_en_0 = _T_811[9]; // @[MemPrimitives.scala 96:27:@16249.4]
  assign Mem1D_3_clock = clock; // @[:@15992.4]
  assign Mem1D_3_reset = reset; // @[:@15993.4]
  assign Mem1D_3_io_r_ofs_0 = _T_1188[0]; // @[MemPrimitives.scala 127:28:@16620.4]
  assign Mem1D_3_io_r_backpressure = _T_1188[1]; // @[MemPrimitives.scala 128:32:@16621.4]
  assign Mem1D_3_io_w_ofs_0 = _T_829[0]; // @[MemPrimitives.scala 94:28:@16264.4]
  assign Mem1D_3_io_w_data_0 = _T_829[8:1]; // @[MemPrimitives.scala 95:29:@16265.4]
  assign Mem1D_3_io_w_en_0 = _T_829[9]; // @[MemPrimitives.scala 96:27:@16266.4]
  assign Mem1D_4_clock = clock; // @[:@16008.4]
  assign Mem1D_4_reset = reset; // @[:@16009.4]
  assign Mem1D_4_io_r_ofs_0 = _T_1217[0]; // @[MemPrimitives.scala 127:28:@16652.4]
  assign Mem1D_4_io_r_backpressure = _T_1217[1]; // @[MemPrimitives.scala 128:32:@16653.4]
  assign Mem1D_4_io_w_ofs_0 = _T_847[0]; // @[MemPrimitives.scala 94:28:@16281.4]
  assign Mem1D_4_io_w_data_0 = _T_847[8:1]; // @[MemPrimitives.scala 95:29:@16282.4]
  assign Mem1D_4_io_w_en_0 = _T_847[9]; // @[MemPrimitives.scala 96:27:@16283.4]
  assign Mem1D_5_clock = clock; // @[:@16024.4]
  assign Mem1D_5_reset = reset; // @[:@16025.4]
  assign Mem1D_5_io_r_ofs_0 = _T_1246[0]; // @[MemPrimitives.scala 127:28:@16684.4]
  assign Mem1D_5_io_r_backpressure = _T_1246[1]; // @[MemPrimitives.scala 128:32:@16685.4]
  assign Mem1D_5_io_w_ofs_0 = _T_865[0]; // @[MemPrimitives.scala 94:28:@16298.4]
  assign Mem1D_5_io_w_data_0 = _T_865[8:1]; // @[MemPrimitives.scala 95:29:@16299.4]
  assign Mem1D_5_io_w_en_0 = _T_865[9]; // @[MemPrimitives.scala 96:27:@16300.4]
  assign Mem1D_6_clock = clock; // @[:@16040.4]
  assign Mem1D_6_reset = reset; // @[:@16041.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1275[0]; // @[MemPrimitives.scala 127:28:@16716.4]
  assign Mem1D_6_io_r_backpressure = _T_1275[1]; // @[MemPrimitives.scala 128:32:@16717.4]
  assign Mem1D_6_io_w_ofs_0 = _T_883[0]; // @[MemPrimitives.scala 94:28:@16315.4]
  assign Mem1D_6_io_w_data_0 = _T_883[8:1]; // @[MemPrimitives.scala 95:29:@16316.4]
  assign Mem1D_6_io_w_en_0 = _T_883[9]; // @[MemPrimitives.scala 96:27:@16317.4]
  assign Mem1D_7_clock = clock; // @[:@16056.4]
  assign Mem1D_7_reset = reset; // @[:@16057.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1331[0]; // @[MemPrimitives.scala 127:28:@16772.4]
  assign Mem1D_7_io_r_backpressure = _T_1331[1]; // @[MemPrimitives.scala 128:32:@16773.4]
  assign Mem1D_7_io_w_ofs_0 = _T_901[0]; // @[MemPrimitives.scala 94:28:@16332.4]
  assign Mem1D_7_io_w_data_0 = _T_901[8:1]; // @[MemPrimitives.scala 95:29:@16333.4]
  assign Mem1D_7_io_w_en_0 = _T_901[9]; // @[MemPrimitives.scala 96:27:@16334.4]
  assign Mem1D_8_clock = clock; // @[:@16072.4]
  assign Mem1D_8_reset = reset; // @[:@16073.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1360[0]; // @[MemPrimitives.scala 127:28:@16804.4]
  assign Mem1D_8_io_r_backpressure = _T_1360[1]; // @[MemPrimitives.scala 128:32:@16805.4]
  assign Mem1D_8_io_w_ofs_0 = _T_919[0]; // @[MemPrimitives.scala 94:28:@16349.4]
  assign Mem1D_8_io_w_data_0 = _T_919[8:1]; // @[MemPrimitives.scala 95:29:@16350.4]
  assign Mem1D_8_io_w_en_0 = _T_919[9]; // @[MemPrimitives.scala 96:27:@16351.4]
  assign Mem1D_9_clock = clock; // @[:@16088.4]
  assign Mem1D_9_reset = reset; // @[:@16089.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1389[0]; // @[MemPrimitives.scala 127:28:@16836.4]
  assign Mem1D_9_io_r_backpressure = _T_1389[1]; // @[MemPrimitives.scala 128:32:@16837.4]
  assign Mem1D_9_io_w_ofs_0 = _T_937[0]; // @[MemPrimitives.scala 94:28:@16366.4]
  assign Mem1D_9_io_w_data_0 = _T_937[8:1]; // @[MemPrimitives.scala 95:29:@16367.4]
  assign Mem1D_9_io_w_en_0 = _T_937[9]; // @[MemPrimitives.scala 96:27:@16368.4]
  assign Mem1D_10_clock = clock; // @[:@16104.4]
  assign Mem1D_10_reset = reset; // @[:@16105.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1418[0]; // @[MemPrimitives.scala 127:28:@16868.4]
  assign Mem1D_10_io_r_backpressure = _T_1418[1]; // @[MemPrimitives.scala 128:32:@16869.4]
  assign Mem1D_10_io_w_ofs_0 = _T_955[0]; // @[MemPrimitives.scala 94:28:@16383.4]
  assign Mem1D_10_io_w_data_0 = _T_955[8:1]; // @[MemPrimitives.scala 95:29:@16384.4]
  assign Mem1D_10_io_w_en_0 = _T_955[9]; // @[MemPrimitives.scala 96:27:@16385.4]
  assign Mem1D_11_clock = clock; // @[:@16120.4]
  assign Mem1D_11_reset = reset; // @[:@16121.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1474[0]; // @[MemPrimitives.scala 127:28:@16924.4]
  assign Mem1D_11_io_r_backpressure = _T_1474[1]; // @[MemPrimitives.scala 128:32:@16925.4]
  assign Mem1D_11_io_w_ofs_0 = _T_973[0]; // @[MemPrimitives.scala 94:28:@16400.4]
  assign Mem1D_11_io_w_data_0 = _T_973[8:1]; // @[MemPrimitives.scala 95:29:@16401.4]
  assign Mem1D_11_io_w_en_0 = _T_973[9]; // @[MemPrimitives.scala 96:27:@16402.4]
  assign Mem1D_12_clock = clock; // @[:@16136.4]
  assign Mem1D_12_reset = reset; // @[:@16137.4]
  assign Mem1D_12_io_r_ofs_0 = _T_1503[0]; // @[MemPrimitives.scala 127:28:@16956.4]
  assign Mem1D_12_io_r_backpressure = _T_1503[1]; // @[MemPrimitives.scala 128:32:@16957.4]
  assign Mem1D_12_io_w_ofs_0 = _T_991[0]; // @[MemPrimitives.scala 94:28:@16417.4]
  assign Mem1D_12_io_w_data_0 = _T_991[8:1]; // @[MemPrimitives.scala 95:29:@16418.4]
  assign Mem1D_12_io_w_en_0 = _T_991[9]; // @[MemPrimitives.scala 96:27:@16419.4]
  assign Mem1D_13_clock = clock; // @[:@16152.4]
  assign Mem1D_13_reset = reset; // @[:@16153.4]
  assign Mem1D_13_io_r_ofs_0 = _T_1532[0]; // @[MemPrimitives.scala 127:28:@16988.4]
  assign Mem1D_13_io_r_backpressure = _T_1532[1]; // @[MemPrimitives.scala 128:32:@16989.4]
  assign Mem1D_13_io_w_ofs_0 = _T_1009[0]; // @[MemPrimitives.scala 94:28:@16434.4]
  assign Mem1D_13_io_w_data_0 = _T_1009[8:1]; // @[MemPrimitives.scala 95:29:@16435.4]
  assign Mem1D_13_io_w_en_0 = _T_1009[9]; // @[MemPrimitives.scala 96:27:@16436.4]
  assign Mem1D_14_clock = clock; // @[:@16168.4]
  assign Mem1D_14_reset = reset; // @[:@16169.4]
  assign Mem1D_14_io_r_ofs_0 = _T_1561[0]; // @[MemPrimitives.scala 127:28:@17020.4]
  assign Mem1D_14_io_r_backpressure = _T_1561[1]; // @[MemPrimitives.scala 128:32:@17021.4]
  assign Mem1D_14_io_w_ofs_0 = _T_1027[0]; // @[MemPrimitives.scala 94:28:@16451.4]
  assign Mem1D_14_io_w_data_0 = _T_1027[8:1]; // @[MemPrimitives.scala 95:29:@16452.4]
  assign Mem1D_14_io_w_en_0 = _T_1027[9]; // @[MemPrimitives.scala 96:27:@16453.4]
  assign Mem1D_15_clock = clock; // @[:@16184.4]
  assign Mem1D_15_reset = reset; // @[:@16185.4]
  assign Mem1D_15_io_r_ofs_0 = _T_1617[0]; // @[MemPrimitives.scala 127:28:@17076.4]
  assign Mem1D_15_io_r_backpressure = _T_1617[1]; // @[MemPrimitives.scala 128:32:@17077.4]
  assign Mem1D_15_io_w_ofs_0 = _T_1045[0]; // @[MemPrimitives.scala 94:28:@16468.4]
  assign Mem1D_15_io_w_data_0 = _T_1045[8:1]; // @[MemPrimitives.scala 95:29:@16469.4]
  assign Mem1D_15_io_w_en_0 = _T_1045[9]; // @[MemPrimitives.scala 96:27:@16470.4]
  assign StickySelects_clock = clock; // @[:@16481.4]
  assign StickySelects_reset = reset; // @[:@16482.4]
  assign StickySelects_io_ins_0 = io_rPort_4_en_0 & _T_1050; // @[MemPrimitives.scala 122:60:@16483.4]
  assign StickySelects_io_ins_1 = io_rPort_9_en_0 & _T_1055; // @[MemPrimitives.scala 122:60:@16484.4]
  assign StickySelects_io_ins_2 = io_rPort_10_en_0 & _T_1060; // @[MemPrimitives.scala 122:60:@16485.4]
  assign StickySelects_1_clock = clock; // @[:@16513.4]
  assign StickySelects_1_reset = reset; // @[:@16514.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_1079; // @[MemPrimitives.scala 122:60:@16515.4]
  assign StickySelects_1_io_ins_1 = io_rPort_3_en_0 & _T_1084; // @[MemPrimitives.scala 122:60:@16516.4]
  assign StickySelects_1_io_ins_2 = io_rPort_14_en_0 & _T_1089; // @[MemPrimitives.scala 122:60:@16517.4]
  assign StickySelects_2_clock = clock; // @[:@16545.4]
  assign StickySelects_2_reset = reset; // @[:@16546.4]
  assign StickySelects_2_io_ins_0 = io_rPort_6_en_0 & _T_1108; // @[MemPrimitives.scala 122:60:@16547.4]
  assign StickySelects_2_io_ins_1 = io_rPort_12_en_0 & _T_1113; // @[MemPrimitives.scala 122:60:@16548.4]
  assign StickySelects_2_io_ins_2 = io_rPort_13_en_0 & _T_1118; // @[MemPrimitives.scala 122:60:@16549.4]
  assign StickySelects_3_clock = clock; // @[:@16586.4]
  assign StickySelects_3_reset = reset; // @[:@16587.4]
  assign StickySelects_3_io_ins_0 = io_rPort_1_en_0 & _T_1137; // @[MemPrimitives.scala 122:60:@16588.4]
  assign StickySelects_3_io_ins_1 = io_rPort_2_en_0 & _T_1142; // @[MemPrimitives.scala 122:60:@16589.4]
  assign StickySelects_3_io_ins_2 = io_rPort_5_en_0 & _T_1147; // @[MemPrimitives.scala 122:60:@16590.4]
  assign StickySelects_3_io_ins_3 = io_rPort_7_en_0 & _T_1152; // @[MemPrimitives.scala 122:60:@16591.4]
  assign StickySelects_3_io_ins_4 = io_rPort_8_en_0 & _T_1157; // @[MemPrimitives.scala 122:60:@16592.4]
  assign StickySelects_3_io_ins_5 = io_rPort_11_en_0 & _T_1162; // @[MemPrimitives.scala 122:60:@16593.4]
  assign StickySelects_4_clock = clock; // @[:@16633.4]
  assign StickySelects_4_reset = reset; // @[:@16634.4]
  assign StickySelects_4_io_ins_0 = io_rPort_4_en_0 & _T_1193; // @[MemPrimitives.scala 122:60:@16635.4]
  assign StickySelects_4_io_ins_1 = io_rPort_9_en_0 & _T_1198; // @[MemPrimitives.scala 122:60:@16636.4]
  assign StickySelects_4_io_ins_2 = io_rPort_10_en_0 & _T_1203; // @[MemPrimitives.scala 122:60:@16637.4]
  assign StickySelects_5_clock = clock; // @[:@16665.4]
  assign StickySelects_5_reset = reset; // @[:@16666.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_1222; // @[MemPrimitives.scala 122:60:@16667.4]
  assign StickySelects_5_io_ins_1 = io_rPort_3_en_0 & _T_1227; // @[MemPrimitives.scala 122:60:@16668.4]
  assign StickySelects_5_io_ins_2 = io_rPort_14_en_0 & _T_1232; // @[MemPrimitives.scala 122:60:@16669.4]
  assign StickySelects_6_clock = clock; // @[:@16697.4]
  assign StickySelects_6_reset = reset; // @[:@16698.4]
  assign StickySelects_6_io_ins_0 = io_rPort_6_en_0 & _T_1251; // @[MemPrimitives.scala 122:60:@16699.4]
  assign StickySelects_6_io_ins_1 = io_rPort_12_en_0 & _T_1256; // @[MemPrimitives.scala 122:60:@16700.4]
  assign StickySelects_6_io_ins_2 = io_rPort_13_en_0 & _T_1261; // @[MemPrimitives.scala 122:60:@16701.4]
  assign StickySelects_7_clock = clock; // @[:@16738.4]
  assign StickySelects_7_reset = reset; // @[:@16739.4]
  assign StickySelects_7_io_ins_0 = io_rPort_1_en_0 & _T_1280; // @[MemPrimitives.scala 122:60:@16740.4]
  assign StickySelects_7_io_ins_1 = io_rPort_2_en_0 & _T_1285; // @[MemPrimitives.scala 122:60:@16741.4]
  assign StickySelects_7_io_ins_2 = io_rPort_5_en_0 & _T_1290; // @[MemPrimitives.scala 122:60:@16742.4]
  assign StickySelects_7_io_ins_3 = io_rPort_7_en_0 & _T_1295; // @[MemPrimitives.scala 122:60:@16743.4]
  assign StickySelects_7_io_ins_4 = io_rPort_8_en_0 & _T_1300; // @[MemPrimitives.scala 122:60:@16744.4]
  assign StickySelects_7_io_ins_5 = io_rPort_11_en_0 & _T_1305; // @[MemPrimitives.scala 122:60:@16745.4]
  assign StickySelects_8_clock = clock; // @[:@16785.4]
  assign StickySelects_8_reset = reset; // @[:@16786.4]
  assign StickySelects_8_io_ins_0 = io_rPort_4_en_0 & _T_1336; // @[MemPrimitives.scala 122:60:@16787.4]
  assign StickySelects_8_io_ins_1 = io_rPort_9_en_0 & _T_1341; // @[MemPrimitives.scala 122:60:@16788.4]
  assign StickySelects_8_io_ins_2 = io_rPort_10_en_0 & _T_1346; // @[MemPrimitives.scala 122:60:@16789.4]
  assign StickySelects_9_clock = clock; // @[:@16817.4]
  assign StickySelects_9_reset = reset; // @[:@16818.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_1365; // @[MemPrimitives.scala 122:60:@16819.4]
  assign StickySelects_9_io_ins_1 = io_rPort_3_en_0 & _T_1370; // @[MemPrimitives.scala 122:60:@16820.4]
  assign StickySelects_9_io_ins_2 = io_rPort_14_en_0 & _T_1375; // @[MemPrimitives.scala 122:60:@16821.4]
  assign StickySelects_10_clock = clock; // @[:@16849.4]
  assign StickySelects_10_reset = reset; // @[:@16850.4]
  assign StickySelects_10_io_ins_0 = io_rPort_6_en_0 & _T_1394; // @[MemPrimitives.scala 122:60:@16851.4]
  assign StickySelects_10_io_ins_1 = io_rPort_12_en_0 & _T_1399; // @[MemPrimitives.scala 122:60:@16852.4]
  assign StickySelects_10_io_ins_2 = io_rPort_13_en_0 & _T_1404; // @[MemPrimitives.scala 122:60:@16853.4]
  assign StickySelects_11_clock = clock; // @[:@16890.4]
  assign StickySelects_11_reset = reset; // @[:@16891.4]
  assign StickySelects_11_io_ins_0 = io_rPort_1_en_0 & _T_1423; // @[MemPrimitives.scala 122:60:@16892.4]
  assign StickySelects_11_io_ins_1 = io_rPort_2_en_0 & _T_1428; // @[MemPrimitives.scala 122:60:@16893.4]
  assign StickySelects_11_io_ins_2 = io_rPort_5_en_0 & _T_1433; // @[MemPrimitives.scala 122:60:@16894.4]
  assign StickySelects_11_io_ins_3 = io_rPort_7_en_0 & _T_1438; // @[MemPrimitives.scala 122:60:@16895.4]
  assign StickySelects_11_io_ins_4 = io_rPort_8_en_0 & _T_1443; // @[MemPrimitives.scala 122:60:@16896.4]
  assign StickySelects_11_io_ins_5 = io_rPort_11_en_0 & _T_1448; // @[MemPrimitives.scala 122:60:@16897.4]
  assign StickySelects_12_clock = clock; // @[:@16937.4]
  assign StickySelects_12_reset = reset; // @[:@16938.4]
  assign StickySelects_12_io_ins_0 = io_rPort_4_en_0 & _T_1479; // @[MemPrimitives.scala 122:60:@16939.4]
  assign StickySelects_12_io_ins_1 = io_rPort_9_en_0 & _T_1484; // @[MemPrimitives.scala 122:60:@16940.4]
  assign StickySelects_12_io_ins_2 = io_rPort_10_en_0 & _T_1489; // @[MemPrimitives.scala 122:60:@16941.4]
  assign StickySelects_13_clock = clock; // @[:@16969.4]
  assign StickySelects_13_reset = reset; // @[:@16970.4]
  assign StickySelects_13_io_ins_0 = io_rPort_0_en_0 & _T_1508; // @[MemPrimitives.scala 122:60:@16971.4]
  assign StickySelects_13_io_ins_1 = io_rPort_3_en_0 & _T_1513; // @[MemPrimitives.scala 122:60:@16972.4]
  assign StickySelects_13_io_ins_2 = io_rPort_14_en_0 & _T_1518; // @[MemPrimitives.scala 122:60:@16973.4]
  assign StickySelects_14_clock = clock; // @[:@17001.4]
  assign StickySelects_14_reset = reset; // @[:@17002.4]
  assign StickySelects_14_io_ins_0 = io_rPort_6_en_0 & _T_1537; // @[MemPrimitives.scala 122:60:@17003.4]
  assign StickySelects_14_io_ins_1 = io_rPort_12_en_0 & _T_1542; // @[MemPrimitives.scala 122:60:@17004.4]
  assign StickySelects_14_io_ins_2 = io_rPort_13_en_0 & _T_1547; // @[MemPrimitives.scala 122:60:@17005.4]
  assign StickySelects_15_clock = clock; // @[:@17042.4]
  assign StickySelects_15_reset = reset; // @[:@17043.4]
  assign StickySelects_15_io_ins_0 = io_rPort_1_en_0 & _T_1566; // @[MemPrimitives.scala 122:60:@17044.4]
  assign StickySelects_15_io_ins_1 = io_rPort_2_en_0 & _T_1571; // @[MemPrimitives.scala 122:60:@17045.4]
  assign StickySelects_15_io_ins_2 = io_rPort_5_en_0 & _T_1576; // @[MemPrimitives.scala 122:60:@17046.4]
  assign StickySelects_15_io_ins_3 = io_rPort_7_en_0 & _T_1581; // @[MemPrimitives.scala 122:60:@17047.4]
  assign StickySelects_15_io_ins_4 = io_rPort_8_en_0 & _T_1586; // @[MemPrimitives.scala 122:60:@17048.4]
  assign StickySelects_15_io_ins_5 = io_rPort_11_en_0 & _T_1591; // @[MemPrimitives.scala 122:60:@17049.4]
  assign RetimeWrapper_clock = clock; // @[:@17093.4]
  assign RetimeWrapper_reset = reset; // @[:@17094.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@17096.4]
  assign RetimeWrapper_io_in = _T_1079 & io_rPort_0_en_0; // @[package.scala 94:16:@17095.4]
  assign RetimeWrapper_1_clock = clock; // @[:@17101.4]
  assign RetimeWrapper_1_reset = reset; // @[:@17102.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@17104.4]
  assign RetimeWrapper_1_io_in = _T_1222 & io_rPort_0_en_0; // @[package.scala 94:16:@17103.4]
  assign RetimeWrapper_2_clock = clock; // @[:@17109.4]
  assign RetimeWrapper_2_reset = reset; // @[:@17110.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@17112.4]
  assign RetimeWrapper_2_io_in = _T_1365 & io_rPort_0_en_0; // @[package.scala 94:16:@17111.4]
  assign RetimeWrapper_3_clock = clock; // @[:@17117.4]
  assign RetimeWrapper_3_reset = reset; // @[:@17118.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@17120.4]
  assign RetimeWrapper_3_io_in = _T_1508 & io_rPort_0_en_0; // @[package.scala 94:16:@17119.4]
  assign RetimeWrapper_4_clock = clock; // @[:@17141.4]
  assign RetimeWrapper_4_reset = reset; // @[:@17142.4]
  assign RetimeWrapper_4_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@17144.4]
  assign RetimeWrapper_4_io_in = _T_1137 & io_rPort_1_en_0; // @[package.scala 94:16:@17143.4]
  assign RetimeWrapper_5_clock = clock; // @[:@17149.4]
  assign RetimeWrapper_5_reset = reset; // @[:@17150.4]
  assign RetimeWrapper_5_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@17152.4]
  assign RetimeWrapper_5_io_in = _T_1280 & io_rPort_1_en_0; // @[package.scala 94:16:@17151.4]
  assign RetimeWrapper_6_clock = clock; // @[:@17157.4]
  assign RetimeWrapper_6_reset = reset; // @[:@17158.4]
  assign RetimeWrapper_6_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@17160.4]
  assign RetimeWrapper_6_io_in = _T_1423 & io_rPort_1_en_0; // @[package.scala 94:16:@17159.4]
  assign RetimeWrapper_7_clock = clock; // @[:@17165.4]
  assign RetimeWrapper_7_reset = reset; // @[:@17166.4]
  assign RetimeWrapper_7_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@17168.4]
  assign RetimeWrapper_7_io_in = _T_1566 & io_rPort_1_en_0; // @[package.scala 94:16:@17167.4]
  assign RetimeWrapper_8_clock = clock; // @[:@17189.4]
  assign RetimeWrapper_8_reset = reset; // @[:@17190.4]
  assign RetimeWrapper_8_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@17192.4]
  assign RetimeWrapper_8_io_in = _T_1142 & io_rPort_2_en_0; // @[package.scala 94:16:@17191.4]
  assign RetimeWrapper_9_clock = clock; // @[:@17197.4]
  assign RetimeWrapper_9_reset = reset; // @[:@17198.4]
  assign RetimeWrapper_9_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@17200.4]
  assign RetimeWrapper_9_io_in = _T_1285 & io_rPort_2_en_0; // @[package.scala 94:16:@17199.4]
  assign RetimeWrapper_10_clock = clock; // @[:@17205.4]
  assign RetimeWrapper_10_reset = reset; // @[:@17206.4]
  assign RetimeWrapper_10_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@17208.4]
  assign RetimeWrapper_10_io_in = _T_1428 & io_rPort_2_en_0; // @[package.scala 94:16:@17207.4]
  assign RetimeWrapper_11_clock = clock; // @[:@17213.4]
  assign RetimeWrapper_11_reset = reset; // @[:@17214.4]
  assign RetimeWrapper_11_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@17216.4]
  assign RetimeWrapper_11_io_in = _T_1571 & io_rPort_2_en_0; // @[package.scala 94:16:@17215.4]
  assign RetimeWrapper_12_clock = clock; // @[:@17237.4]
  assign RetimeWrapper_12_reset = reset; // @[:@17238.4]
  assign RetimeWrapper_12_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@17240.4]
  assign RetimeWrapper_12_io_in = _T_1084 & io_rPort_3_en_0; // @[package.scala 94:16:@17239.4]
  assign RetimeWrapper_13_clock = clock; // @[:@17245.4]
  assign RetimeWrapper_13_reset = reset; // @[:@17246.4]
  assign RetimeWrapper_13_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@17248.4]
  assign RetimeWrapper_13_io_in = _T_1227 & io_rPort_3_en_0; // @[package.scala 94:16:@17247.4]
  assign RetimeWrapper_14_clock = clock; // @[:@17253.4]
  assign RetimeWrapper_14_reset = reset; // @[:@17254.4]
  assign RetimeWrapper_14_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@17256.4]
  assign RetimeWrapper_14_io_in = _T_1370 & io_rPort_3_en_0; // @[package.scala 94:16:@17255.4]
  assign RetimeWrapper_15_clock = clock; // @[:@17261.4]
  assign RetimeWrapper_15_reset = reset; // @[:@17262.4]
  assign RetimeWrapper_15_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@17264.4]
  assign RetimeWrapper_15_io_in = _T_1513 & io_rPort_3_en_0; // @[package.scala 94:16:@17263.4]
  assign RetimeWrapper_16_clock = clock; // @[:@17285.4]
  assign RetimeWrapper_16_reset = reset; // @[:@17286.4]
  assign RetimeWrapper_16_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@17288.4]
  assign RetimeWrapper_16_io_in = _T_1050 & io_rPort_4_en_0; // @[package.scala 94:16:@17287.4]
  assign RetimeWrapper_17_clock = clock; // @[:@17293.4]
  assign RetimeWrapper_17_reset = reset; // @[:@17294.4]
  assign RetimeWrapper_17_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@17296.4]
  assign RetimeWrapper_17_io_in = _T_1193 & io_rPort_4_en_0; // @[package.scala 94:16:@17295.4]
  assign RetimeWrapper_18_clock = clock; // @[:@17301.4]
  assign RetimeWrapper_18_reset = reset; // @[:@17302.4]
  assign RetimeWrapper_18_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@17304.4]
  assign RetimeWrapper_18_io_in = _T_1336 & io_rPort_4_en_0; // @[package.scala 94:16:@17303.4]
  assign RetimeWrapper_19_clock = clock; // @[:@17309.4]
  assign RetimeWrapper_19_reset = reset; // @[:@17310.4]
  assign RetimeWrapper_19_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@17312.4]
  assign RetimeWrapper_19_io_in = _T_1479 & io_rPort_4_en_0; // @[package.scala 94:16:@17311.4]
  assign RetimeWrapper_20_clock = clock; // @[:@17333.4]
  assign RetimeWrapper_20_reset = reset; // @[:@17334.4]
  assign RetimeWrapper_20_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@17336.4]
  assign RetimeWrapper_20_io_in = _T_1147 & io_rPort_5_en_0; // @[package.scala 94:16:@17335.4]
  assign RetimeWrapper_21_clock = clock; // @[:@17341.4]
  assign RetimeWrapper_21_reset = reset; // @[:@17342.4]
  assign RetimeWrapper_21_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@17344.4]
  assign RetimeWrapper_21_io_in = _T_1290 & io_rPort_5_en_0; // @[package.scala 94:16:@17343.4]
  assign RetimeWrapper_22_clock = clock; // @[:@17349.4]
  assign RetimeWrapper_22_reset = reset; // @[:@17350.4]
  assign RetimeWrapper_22_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@17352.4]
  assign RetimeWrapper_22_io_in = _T_1433 & io_rPort_5_en_0; // @[package.scala 94:16:@17351.4]
  assign RetimeWrapper_23_clock = clock; // @[:@17357.4]
  assign RetimeWrapper_23_reset = reset; // @[:@17358.4]
  assign RetimeWrapper_23_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@17360.4]
  assign RetimeWrapper_23_io_in = _T_1576 & io_rPort_5_en_0; // @[package.scala 94:16:@17359.4]
  assign RetimeWrapper_24_clock = clock; // @[:@17381.4]
  assign RetimeWrapper_24_reset = reset; // @[:@17382.4]
  assign RetimeWrapper_24_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@17384.4]
  assign RetimeWrapper_24_io_in = _T_1108 & io_rPort_6_en_0; // @[package.scala 94:16:@17383.4]
  assign RetimeWrapper_25_clock = clock; // @[:@17389.4]
  assign RetimeWrapper_25_reset = reset; // @[:@17390.4]
  assign RetimeWrapper_25_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@17392.4]
  assign RetimeWrapper_25_io_in = _T_1251 & io_rPort_6_en_0; // @[package.scala 94:16:@17391.4]
  assign RetimeWrapper_26_clock = clock; // @[:@17397.4]
  assign RetimeWrapper_26_reset = reset; // @[:@17398.4]
  assign RetimeWrapper_26_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@17400.4]
  assign RetimeWrapper_26_io_in = _T_1394 & io_rPort_6_en_0; // @[package.scala 94:16:@17399.4]
  assign RetimeWrapper_27_clock = clock; // @[:@17405.4]
  assign RetimeWrapper_27_reset = reset; // @[:@17406.4]
  assign RetimeWrapper_27_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@17408.4]
  assign RetimeWrapper_27_io_in = _T_1537 & io_rPort_6_en_0; // @[package.scala 94:16:@17407.4]
  assign RetimeWrapper_28_clock = clock; // @[:@17429.4]
  assign RetimeWrapper_28_reset = reset; // @[:@17430.4]
  assign RetimeWrapper_28_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@17432.4]
  assign RetimeWrapper_28_io_in = _T_1152 & io_rPort_7_en_0; // @[package.scala 94:16:@17431.4]
  assign RetimeWrapper_29_clock = clock; // @[:@17437.4]
  assign RetimeWrapper_29_reset = reset; // @[:@17438.4]
  assign RetimeWrapper_29_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@17440.4]
  assign RetimeWrapper_29_io_in = _T_1295 & io_rPort_7_en_0; // @[package.scala 94:16:@17439.4]
  assign RetimeWrapper_30_clock = clock; // @[:@17445.4]
  assign RetimeWrapper_30_reset = reset; // @[:@17446.4]
  assign RetimeWrapper_30_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@17448.4]
  assign RetimeWrapper_30_io_in = _T_1438 & io_rPort_7_en_0; // @[package.scala 94:16:@17447.4]
  assign RetimeWrapper_31_clock = clock; // @[:@17453.4]
  assign RetimeWrapper_31_reset = reset; // @[:@17454.4]
  assign RetimeWrapper_31_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@17456.4]
  assign RetimeWrapper_31_io_in = _T_1581 & io_rPort_7_en_0; // @[package.scala 94:16:@17455.4]
  assign RetimeWrapper_32_clock = clock; // @[:@17477.4]
  assign RetimeWrapper_32_reset = reset; // @[:@17478.4]
  assign RetimeWrapper_32_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@17480.4]
  assign RetimeWrapper_32_io_in = _T_1157 & io_rPort_8_en_0; // @[package.scala 94:16:@17479.4]
  assign RetimeWrapper_33_clock = clock; // @[:@17485.4]
  assign RetimeWrapper_33_reset = reset; // @[:@17486.4]
  assign RetimeWrapper_33_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@17488.4]
  assign RetimeWrapper_33_io_in = _T_1300 & io_rPort_8_en_0; // @[package.scala 94:16:@17487.4]
  assign RetimeWrapper_34_clock = clock; // @[:@17493.4]
  assign RetimeWrapper_34_reset = reset; // @[:@17494.4]
  assign RetimeWrapper_34_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@17496.4]
  assign RetimeWrapper_34_io_in = _T_1443 & io_rPort_8_en_0; // @[package.scala 94:16:@17495.4]
  assign RetimeWrapper_35_clock = clock; // @[:@17501.4]
  assign RetimeWrapper_35_reset = reset; // @[:@17502.4]
  assign RetimeWrapper_35_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@17504.4]
  assign RetimeWrapper_35_io_in = _T_1586 & io_rPort_8_en_0; // @[package.scala 94:16:@17503.4]
  assign RetimeWrapper_36_clock = clock; // @[:@17525.4]
  assign RetimeWrapper_36_reset = reset; // @[:@17526.4]
  assign RetimeWrapper_36_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@17528.4]
  assign RetimeWrapper_36_io_in = _T_1055 & io_rPort_9_en_0; // @[package.scala 94:16:@17527.4]
  assign RetimeWrapper_37_clock = clock; // @[:@17533.4]
  assign RetimeWrapper_37_reset = reset; // @[:@17534.4]
  assign RetimeWrapper_37_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@17536.4]
  assign RetimeWrapper_37_io_in = _T_1198 & io_rPort_9_en_0; // @[package.scala 94:16:@17535.4]
  assign RetimeWrapper_38_clock = clock; // @[:@17541.4]
  assign RetimeWrapper_38_reset = reset; // @[:@17542.4]
  assign RetimeWrapper_38_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@17544.4]
  assign RetimeWrapper_38_io_in = _T_1341 & io_rPort_9_en_0; // @[package.scala 94:16:@17543.4]
  assign RetimeWrapper_39_clock = clock; // @[:@17549.4]
  assign RetimeWrapper_39_reset = reset; // @[:@17550.4]
  assign RetimeWrapper_39_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@17552.4]
  assign RetimeWrapper_39_io_in = _T_1484 & io_rPort_9_en_0; // @[package.scala 94:16:@17551.4]
  assign RetimeWrapper_40_clock = clock; // @[:@17573.4]
  assign RetimeWrapper_40_reset = reset; // @[:@17574.4]
  assign RetimeWrapper_40_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@17576.4]
  assign RetimeWrapper_40_io_in = _T_1060 & io_rPort_10_en_0; // @[package.scala 94:16:@17575.4]
  assign RetimeWrapper_41_clock = clock; // @[:@17581.4]
  assign RetimeWrapper_41_reset = reset; // @[:@17582.4]
  assign RetimeWrapper_41_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@17584.4]
  assign RetimeWrapper_41_io_in = _T_1203 & io_rPort_10_en_0; // @[package.scala 94:16:@17583.4]
  assign RetimeWrapper_42_clock = clock; // @[:@17589.4]
  assign RetimeWrapper_42_reset = reset; // @[:@17590.4]
  assign RetimeWrapper_42_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@17592.4]
  assign RetimeWrapper_42_io_in = _T_1346 & io_rPort_10_en_0; // @[package.scala 94:16:@17591.4]
  assign RetimeWrapper_43_clock = clock; // @[:@17597.4]
  assign RetimeWrapper_43_reset = reset; // @[:@17598.4]
  assign RetimeWrapper_43_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@17600.4]
  assign RetimeWrapper_43_io_in = _T_1489 & io_rPort_10_en_0; // @[package.scala 94:16:@17599.4]
  assign RetimeWrapper_44_clock = clock; // @[:@17621.4]
  assign RetimeWrapper_44_reset = reset; // @[:@17622.4]
  assign RetimeWrapper_44_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@17624.4]
  assign RetimeWrapper_44_io_in = _T_1162 & io_rPort_11_en_0; // @[package.scala 94:16:@17623.4]
  assign RetimeWrapper_45_clock = clock; // @[:@17629.4]
  assign RetimeWrapper_45_reset = reset; // @[:@17630.4]
  assign RetimeWrapper_45_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@17632.4]
  assign RetimeWrapper_45_io_in = _T_1305 & io_rPort_11_en_0; // @[package.scala 94:16:@17631.4]
  assign RetimeWrapper_46_clock = clock; // @[:@17637.4]
  assign RetimeWrapper_46_reset = reset; // @[:@17638.4]
  assign RetimeWrapper_46_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@17640.4]
  assign RetimeWrapper_46_io_in = _T_1448 & io_rPort_11_en_0; // @[package.scala 94:16:@17639.4]
  assign RetimeWrapper_47_clock = clock; // @[:@17645.4]
  assign RetimeWrapper_47_reset = reset; // @[:@17646.4]
  assign RetimeWrapper_47_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@17648.4]
  assign RetimeWrapper_47_io_in = _T_1591 & io_rPort_11_en_0; // @[package.scala 94:16:@17647.4]
  assign RetimeWrapper_48_clock = clock; // @[:@17669.4]
  assign RetimeWrapper_48_reset = reset; // @[:@17670.4]
  assign RetimeWrapper_48_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@17672.4]
  assign RetimeWrapper_48_io_in = _T_1113 & io_rPort_12_en_0; // @[package.scala 94:16:@17671.4]
  assign RetimeWrapper_49_clock = clock; // @[:@17677.4]
  assign RetimeWrapper_49_reset = reset; // @[:@17678.4]
  assign RetimeWrapper_49_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@17680.4]
  assign RetimeWrapper_49_io_in = _T_1256 & io_rPort_12_en_0; // @[package.scala 94:16:@17679.4]
  assign RetimeWrapper_50_clock = clock; // @[:@17685.4]
  assign RetimeWrapper_50_reset = reset; // @[:@17686.4]
  assign RetimeWrapper_50_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@17688.4]
  assign RetimeWrapper_50_io_in = _T_1399 & io_rPort_12_en_0; // @[package.scala 94:16:@17687.4]
  assign RetimeWrapper_51_clock = clock; // @[:@17693.4]
  assign RetimeWrapper_51_reset = reset; // @[:@17694.4]
  assign RetimeWrapper_51_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@17696.4]
  assign RetimeWrapper_51_io_in = _T_1542 & io_rPort_12_en_0; // @[package.scala 94:16:@17695.4]
  assign RetimeWrapper_52_clock = clock; // @[:@17717.4]
  assign RetimeWrapper_52_reset = reset; // @[:@17718.4]
  assign RetimeWrapper_52_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@17720.4]
  assign RetimeWrapper_52_io_in = _T_1118 & io_rPort_13_en_0; // @[package.scala 94:16:@17719.4]
  assign RetimeWrapper_53_clock = clock; // @[:@17725.4]
  assign RetimeWrapper_53_reset = reset; // @[:@17726.4]
  assign RetimeWrapper_53_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@17728.4]
  assign RetimeWrapper_53_io_in = _T_1261 & io_rPort_13_en_0; // @[package.scala 94:16:@17727.4]
  assign RetimeWrapper_54_clock = clock; // @[:@17733.4]
  assign RetimeWrapper_54_reset = reset; // @[:@17734.4]
  assign RetimeWrapper_54_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@17736.4]
  assign RetimeWrapper_54_io_in = _T_1404 & io_rPort_13_en_0; // @[package.scala 94:16:@17735.4]
  assign RetimeWrapper_55_clock = clock; // @[:@17741.4]
  assign RetimeWrapper_55_reset = reset; // @[:@17742.4]
  assign RetimeWrapper_55_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@17744.4]
  assign RetimeWrapper_55_io_in = _T_1547 & io_rPort_13_en_0; // @[package.scala 94:16:@17743.4]
  assign RetimeWrapper_56_clock = clock; // @[:@17765.4]
  assign RetimeWrapper_56_reset = reset; // @[:@17766.4]
  assign RetimeWrapper_56_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@17768.4]
  assign RetimeWrapper_56_io_in = _T_1089 & io_rPort_14_en_0; // @[package.scala 94:16:@17767.4]
  assign RetimeWrapper_57_clock = clock; // @[:@17773.4]
  assign RetimeWrapper_57_reset = reset; // @[:@17774.4]
  assign RetimeWrapper_57_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@17776.4]
  assign RetimeWrapper_57_io_in = _T_1232 & io_rPort_14_en_0; // @[package.scala 94:16:@17775.4]
  assign RetimeWrapper_58_clock = clock; // @[:@17781.4]
  assign RetimeWrapper_58_reset = reset; // @[:@17782.4]
  assign RetimeWrapper_58_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@17784.4]
  assign RetimeWrapper_58_io_in = _T_1375 & io_rPort_14_en_0; // @[package.scala 94:16:@17783.4]
  assign RetimeWrapper_59_clock = clock; // @[:@17789.4]
  assign RetimeWrapper_59_reset = reset; // @[:@17790.4]
  assign RetimeWrapper_59_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@17792.4]
  assign RetimeWrapper_59_io_in = _T_1518 & io_rPort_14_en_0; // @[package.scala 94:16:@17791.4]
endmodule
module RetimeWrapper_240( // @[:@17812.2]
  input         clock, // @[:@17813.4]
  input         reset, // @[:@17814.4]
  input         io_flow, // @[:@17815.4]
  input  [63:0] io_in, // @[:@17815.4]
  output [63:0] io_out // @[:@17815.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17817.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17817.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17817.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17817.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17817.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17817.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@17817.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17830.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17829.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@17828.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17827.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17826.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17824.4]
endmodule
module SimBlackBoxesfix2fixBox_2( // @[:@17832.2]
  input  [31:0] io_a, // @[:@17835.4]
  output [32:0] io_b // @[:@17835.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@17842.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@17842.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@17847.4]
endmodule
module __2( // @[:@17849.2]
  input  [31:0] io_b, // @[:@17852.4]
  output [32:0] io_result // @[:@17852.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@17857.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@17857.4]
  SimBlackBoxesfix2fixBox_2 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@17857.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@17870.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@17865.4]
endmodule
module RetimeWrapper_241( // @[:@17924.2]
  input         clock, // @[:@17925.4]
  input         reset, // @[:@17926.4]
  input         io_flow, // @[:@17927.4]
  input  [31:0] io_in, // @[:@17927.4]
  output [31:0] io_out // @[:@17927.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17929.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17929.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17929.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17929.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17929.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17929.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@17929.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17942.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17941.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17940.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17939.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17938.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17936.4]
endmodule
module fix2fixBox( // @[:@17944.2]
  input         clock, // @[:@17945.4]
  input         reset, // @[:@17946.4]
  input  [32:0] io_a, // @[:@17947.4]
  input         io_flow, // @[:@17947.4]
  output [31:0] io_b // @[:@17947.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@17957.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@17957.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@17957.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@17957.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@17957.4]
  RetimeWrapper_241 RetimeWrapper ( // @[package.scala 93:22:@17957.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@17964.4]
  assign RetimeWrapper_clock = clock; // @[:@17958.4]
  assign RetimeWrapper_reset = reset; // @[:@17959.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@17961.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@17960.4]
endmodule
module x539_sum( // @[:@17966.2]
  input         clock, // @[:@17967.4]
  input         reset, // @[:@17968.4]
  input  [31:0] io_a, // @[:@17969.4]
  input  [31:0] io_b, // @[:@17969.4]
  input         io_flow, // @[:@17969.4]
  output [31:0] io_result // @[:@17969.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@17977.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@17977.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@17984.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@17984.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@18002.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@18002.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@18002.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@18002.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@18002.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@17982.4 Math.scala 713:14:@17983.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@17989.4 Math.scala 713:14:@17990.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@17991.4]
  __2 _ ( // @[Math.scala 709:24:@17977.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@17984.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@18002.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@17982.4 Math.scala 713:14:@17983.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@17989.4 Math.scala 713:14:@17990.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@17991.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@18010.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@17980.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@17987.4]
  assign fix2fixBox_clock = clock; // @[:@18003.4]
  assign fix2fixBox_reset = reset; // @[:@18004.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@18005.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@18008.4]
endmodule
module RetimeWrapper_242( // @[:@18024.2]
  input   clock, // @[:@18025.4]
  input   reset, // @[:@18026.4]
  input   io_flow, // @[:@18027.4]
  input   io_in, // @[:@18027.4]
  output  io_out // @[:@18027.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@18029.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@18029.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@18029.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18029.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18029.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18029.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@18029.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18042.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18041.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@18040.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18039.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18038.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18036.4]
endmodule
module RetimeWrapper_243( // @[:@18056.2]
  input         clock, // @[:@18057.4]
  input         reset, // @[:@18058.4]
  input         io_flow, // @[:@18059.4]
  input  [31:0] io_in, // @[:@18059.4]
  output [31:0] io_out // @[:@18059.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18061.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18061.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18061.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18061.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18061.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18061.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@18061.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18074.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18073.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@18072.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18071.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18070.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18068.4]
endmodule
module RetimeWrapper_244( // @[:@18088.2]
  input        clock, // @[:@18089.4]
  input        reset, // @[:@18090.4]
  input        io_flow, // @[:@18091.4]
  input  [7:0] io_in, // @[:@18091.4]
  output [7:0] io_out // @[:@18091.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18093.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18093.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18093.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18093.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18093.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18093.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@18093.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18106.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18105.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@18104.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18103.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18102.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18100.4]
endmodule
module RetimeWrapper_246( // @[:@18152.2]
  input         clock, // @[:@18153.4]
  input         reset, // @[:@18154.4]
  input         io_flow, // @[:@18155.4]
  input  [31:0] io_in, // @[:@18155.4]
  output [31:0] io_out // @[:@18155.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18157.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18157.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18157.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18157.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18157.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18157.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@18157.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18170.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18169.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@18168.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18167.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18166.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18164.4]
endmodule
module RetimeWrapper_252( // @[:@18640.2]
  input         clock, // @[:@18641.4]
  input         reset, // @[:@18642.4]
  input         io_flow, // @[:@18643.4]
  input  [31:0] io_in, // @[:@18643.4]
  output [31:0] io_out // @[:@18643.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18645.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18645.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18645.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18645.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18645.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18645.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@18645.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18658.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18657.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@18656.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18655.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18654.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18652.4]
endmodule
module RetimeWrapper_283( // @[:@20964.2]
  input         clock, // @[:@20965.4]
  input         reset, // @[:@20966.4]
  input         io_flow, // @[:@20967.4]
  input  [31:0] io_in, // @[:@20967.4]
  output [31:0] io_out // @[:@20967.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20969.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20969.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20969.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20969.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20969.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20969.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(11)) sr ( // @[RetimeShiftRegister.scala 15:20:@20969.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20982.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20981.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@20980.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20979.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20978.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20976.4]
endmodule
module RetimeWrapper_287( // @[:@21240.2]
  input   clock, // @[:@21241.4]
  input   reset, // @[:@21242.4]
  input   io_flow, // @[:@21243.4]
  input   io_in, // @[:@21243.4]
  output  io_out // @[:@21243.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@21245.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@21245.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@21245.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21245.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21245.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21245.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(13)) sr ( // @[RetimeShiftRegister.scala 15:20:@21245.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21258.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21257.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@21256.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21255.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21254.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21252.4]
endmodule
module RetimeWrapper_304( // @[:@22080.2]
  input         clock, // @[:@22081.4]
  input         reset, // @[:@22082.4]
  input         io_flow, // @[:@22083.4]
  input  [31:0] io_in, // @[:@22083.4]
  output [31:0] io_out // @[:@22083.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22085.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22085.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22085.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22085.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22085.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22085.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(12)) sr ( // @[RetimeShiftRegister.scala 15:20:@22085.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22098.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22097.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22096.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22095.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22094.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22092.4]
endmodule
module RetimeWrapper_321( // @[:@23512.2]
  input         clock, // @[:@23513.4]
  input         reset, // @[:@23514.4]
  input         io_flow, // @[:@23515.4]
  input  [31:0] io_in, // @[:@23515.4]
  output [31:0] io_out // @[:@23515.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@23517.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@23517.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@23517.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@23517.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@23517.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@23517.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@23517.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@23530.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@23529.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@23528.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@23527.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@23526.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@23524.4]
endmodule
module SimBlackBoxesfix2fixBox_82( // @[:@28200.2]
  input  [7:0] io_a, // @[:@28203.4]
  output [8:0] io_b // @[:@28203.4]
);
  assign io_b = {1'h0,io_a}; // @[SimBlackBoxes.scala 99:40:@28214.4]
endmodule
module __82( // @[:@28216.2]
  input  [7:0] io_b, // @[:@28219.4]
  output [8:0] io_result // @[:@28219.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@28224.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@28224.4]
  SimBlackBoxesfix2fixBox_82 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@28224.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@28237.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@28232.4]
endmodule
module fix2fixBox_40( // @[:@28310.2]
  input        clock, // @[:@28311.4]
  input        reset, // @[:@28312.4]
  input  [8:0] io_a, // @[:@28313.4]
  input        io_flow, // @[:@28313.4]
  output [7:0] io_b // @[:@28313.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@28323.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@28323.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@28323.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@28323.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@28323.4]
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@28323.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@28330.4]
  assign RetimeWrapper_clock = clock; // @[:@28324.4]
  assign RetimeWrapper_reset = reset; // @[:@28325.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@28327.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@28326.4]
endmodule
module x811_x23( // @[:@28332.2]
  input        clock, // @[:@28333.4]
  input        reset, // @[:@28334.4]
  input  [7:0] io_a, // @[:@28335.4]
  input  [7:0] io_b, // @[:@28335.4]
  input        io_flow, // @[:@28335.4]
  output [7:0] io_result // @[:@28335.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@28343.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@28343.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@28350.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@28350.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@28360.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@28360.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@28360.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@28360.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@28360.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@28348.4 Math.scala 713:14:@28349.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@28355.4 Math.scala 713:14:@28356.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@28357.4]
  __82 _ ( // @[Math.scala 709:24:@28343.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __82 __1 ( // @[Math.scala 709:24:@28350.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_40 fix2fixBox ( // @[Math.scala 141:30:@28360.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@28348.4 Math.scala 713:14:@28349.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@28355.4 Math.scala 713:14:@28356.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@28357.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@28368.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@28346.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@28353.4]
  assign fix2fixBox_clock = clock; // @[:@28361.4]
  assign fix2fixBox_reset = reset; // @[:@28362.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@28363.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@28366.4]
endmodule
module fix2fixBox_44( // @[:@28958.2]
  input  [8:0] io_a, // @[:@28961.4]
  output [7:0] io_b // @[:@28961.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@28971.4]
endmodule
module x815_x23( // @[:@28973.2]
  input  [7:0] io_a, // @[:@28976.4]
  input  [7:0] io_b, // @[:@28976.4]
  output [7:0] io_result // @[:@28976.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@28984.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@28984.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@28991.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@28991.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@29001.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@29001.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@28989.4 Math.scala 713:14:@28990.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@28996.4 Math.scala 713:14:@28997.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@28998.4]
  __82 _ ( // @[Math.scala 709:24:@28984.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __82 __1 ( // @[Math.scala 709:24:@28991.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_44 fix2fixBox ( // @[Math.scala 141:30:@29001.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@28989.4 Math.scala 713:14:@28990.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@28996.4 Math.scala 713:14:@28997.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@28998.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@29009.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@28987.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@28994.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@29004.4]
endmodule
module RetimeWrapper_428( // @[:@38356.2]
  input   clock, // @[:@38357.4]
  input   reset, // @[:@38358.4]
  input   io_flow, // @[:@38359.4]
  input   io_in, // @[:@38359.4]
  output  io_out // @[:@38359.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@38361.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@38361.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@38361.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@38361.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@38361.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@38361.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@38361.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@38374.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@38373.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@38372.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@38371.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@38370.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@38368.4]
endmodule
module RetimeWrapper_429( // @[:@38388.2]
  input         clock, // @[:@38389.4]
  input         reset, // @[:@38390.4]
  input         io_flow, // @[:@38391.4]
  input  [31:0] io_in, // @[:@38391.4]
  output [31:0] io_out // @[:@38391.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@38393.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@38393.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@38393.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@38393.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@38393.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@38393.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@38393.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@38406.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@38405.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@38404.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@38403.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@38402.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@38400.4]
endmodule
module RetimeWrapper_432( // @[:@38484.2]
  input         clock, // @[:@38485.4]
  input         reset, // @[:@38486.4]
  input         io_flow, // @[:@38487.4]
  input  [31:0] io_in, // @[:@38487.4]
  output [31:0] io_out // @[:@38487.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@38489.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@38489.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@38489.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@38489.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@38489.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@38489.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(17)) sr ( // @[RetimeShiftRegister.scala 15:20:@38489.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@38502.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@38501.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@38500.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@38499.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@38498.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@38496.4]
endmodule
module RetimeWrapper_435( // @[:@38580.2]
  input         clock, // @[:@38581.4]
  input         reset, // @[:@38582.4]
  input         io_flow, // @[:@38583.4]
  input  [31:0] io_in, // @[:@38583.4]
  output [31:0] io_out // @[:@38583.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@38585.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@38585.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@38585.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@38585.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@38585.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@38585.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(16)) sr ( // @[RetimeShiftRegister.scala 15:20:@38585.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@38598.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@38597.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@38596.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@38595.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@38594.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@38592.4]
endmodule
module RetimeWrapper_456( // @[:@39252.2]
  input   clock, // @[:@39253.4]
  input   reset, // @[:@39254.4]
  input   io_flow, // @[:@39255.4]
  input   io_in, // @[:@39255.4]
  output  io_out // @[:@39255.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@39257.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@39257.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@39257.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@39257.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@39257.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@39257.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(19)) sr ( // @[RetimeShiftRegister.scala 15:20:@39257.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@39270.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@39269.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@39268.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@39267.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@39266.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@39264.4]
endmodule
module RetimeWrapper_457( // @[:@39284.2]
  input   clock, // @[:@39285.4]
  input   reset, // @[:@39286.4]
  input   io_flow, // @[:@39287.4]
  input   io_in, // @[:@39287.4]
  output  io_out // @[:@39287.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@39289.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@39289.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@39289.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@39289.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@39289.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@39289.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@39289.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@39302.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@39301.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@39300.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@39299.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@39298.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@39296.4]
endmodule
module RetimeWrapper_506( // @[:@41245.2]
  input        clock, // @[:@41246.4]
  input        reset, // @[:@41247.4]
  input        io_flow, // @[:@41248.4]
  input  [7:0] io_in, // @[:@41248.4]
  output [7:0] io_out // @[:@41248.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@41250.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@41250.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@41250.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@41250.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@41250.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@41250.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@41250.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@41263.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@41262.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@41261.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@41260.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@41259.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@41257.4]
endmodule
module SimBlackBoxesfix2fixBox_216( // @[:@41265.2]
  input  [7:0] io_a, // @[:@41268.4]
  output [7:0] io_b // @[:@41268.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@41278.4]
endmodule
module __216( // @[:@41280.2]
  input  [7:0] io_b, // @[:@41283.4]
  output [7:0] io_result // @[:@41283.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@41288.4]
  wire [7:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@41288.4]
  SimBlackBoxesfix2fixBox_216 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@41288.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@41301.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@41296.4]
endmodule
module x951_div( // @[:@41303.2]
  input        clock, // @[:@41304.4]
  input        reset, // @[:@41305.4]
  input  [7:0] io_a, // @[:@41306.4]
  input        io_flow, // @[:@41306.4]
  output [7:0] io_result // @[:@41306.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@41313.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@41313.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@41313.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@41313.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@41313.4]
  wire [7:0] __io_b; // @[Math.scala 709:24:@41323.4]
  wire [7:0] __io_result; // @[Math.scala 709:24:@41323.4]
  RetimeWrapper_506 RetimeWrapper ( // @[package.scala 93:22:@41313.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  __216 _ ( // @[Math.scala 709:24:@41323.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign io_result = __io_result; // @[Math.scala 291:34:@41331.4]
  assign RetimeWrapper_clock = clock; // @[:@41314.4]
  assign RetimeWrapper_reset = reset; // @[:@41315.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@41317.4]
  assign RetimeWrapper_io_in = io_a / 8'h6; // @[package.scala 94:16:@41316.4]
  assign __io_b = RetimeWrapper_io_out; // @[Math.scala 710:17:@41326.4]
endmodule
module RetimeWrapper_514( // @[:@44796.2]
  input         clock, // @[:@44797.4]
  input         reset, // @[:@44798.4]
  input         io_flow, // @[:@44799.4]
  input  [63:0] io_in, // @[:@44799.4]
  output [63:0] io_out // @[:@44799.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@44801.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@44801.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@44801.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@44801.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@44801.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@44801.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@44801.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@44814.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@44813.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@44812.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@44811.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@44810.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@44808.4]
endmodule
module RetimeWrapper_515( // @[:@44828.2]
  input   clock, // @[:@44829.4]
  input   reset, // @[:@44830.4]
  input   io_flow, // @[:@44831.4]
  input   io_in, // @[:@44831.4]
  output  io_out // @[:@44831.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@44833.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@44833.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@44833.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@44833.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@44833.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@44833.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(29)) sr ( // @[RetimeShiftRegister.scala 15:20:@44833.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@44846.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@44845.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@44844.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@44843.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@44842.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@44840.4]
endmodule
module x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@44912.2]
  input          clock, // @[:@44913.4]
  input          reset, // @[:@44914.4]
  output         io_in_x511_TREADY, // @[:@44915.4]
  input  [255:0] io_in_x511_TDATA, // @[:@44915.4]
  input  [7:0]   io_in_x511_TID, // @[:@44915.4]
  input  [7:0]   io_in_x511_TDEST, // @[:@44915.4]
  output         io_in_x512_TVALID, // @[:@44915.4]
  input          io_in_x512_TREADY, // @[:@44915.4]
  output [255:0] io_in_x512_TDATA, // @[:@44915.4]
  input          io_sigsIn_backpressure, // @[:@44915.4]
  input          io_sigsIn_datapathEn, // @[:@44915.4]
  input          io_sigsIn_break, // @[:@44915.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@44915.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@44915.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@44915.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@44915.4]
  input          io_rr // @[:@44915.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@44929.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@44929.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@44941.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@44941.4]
  wire  x524_lb_0_clock; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_reset; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_23_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_23_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_23_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_23_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_23_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_22_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_22_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_22_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_22_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_22_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_21_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_21_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_21_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_21_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_21_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_20_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_20_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_20_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_20_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_20_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_19_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_19_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_19_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_19_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_19_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_18_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_18_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_18_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_18_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_18_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_17_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_17_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_17_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_17_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_17_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_16_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_16_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_16_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_16_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_16_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_15_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_15_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_15_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_15_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_15_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_14_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_14_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_14_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_14_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_14_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_13_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_13_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_13_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_13_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_13_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_12_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_12_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_12_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_12_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_12_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_11_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_11_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_11_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_11_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_11_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_10_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_10_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_10_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_10_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_10_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_9_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_9_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_9_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_9_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_9_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_8_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_8_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_8_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_8_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_8_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_7_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_7_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_7_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_7_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_7_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_6_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_6_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_6_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_6_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_6_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_5_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_5_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_5_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_5_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_5_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_4_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_4_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_4_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_4_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_4_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_3_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_3_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_3_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_3_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_3_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_2_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_2_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_2_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_2_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_2_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_1_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_1_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_1_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_1_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_1_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_rPort_0_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_0_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_0_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_rPort_0_backpressure; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_rPort_0_output_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_wPort_7_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_7_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_wPort_7_data_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_7_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_wPort_6_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_6_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_wPort_6_data_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_6_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_wPort_5_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_5_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_wPort_5_data_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_5_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_wPort_4_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_4_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_wPort_4_data_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_4_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_wPort_3_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_3_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_wPort_3_data_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_3_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_wPort_2_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_2_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_wPort_2_data_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_2_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_wPort_1_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_1_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_wPort_1_data_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_1_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [2:0] x524_lb_0_io_wPort_0_banks_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_0_ofs_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire [7:0] x524_lb_0_io_wPort_0_data_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x524_lb_0_io_wPort_0_en_0; // @[m_x524_lb_0.scala 57:17:@44951.4]
  wire  x525_lb2_0_clock; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_reset; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_rPort_14_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_14_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_14_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_14_backpressure; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_rPort_14_output_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_rPort_13_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_13_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_13_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_13_backpressure; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_rPort_13_output_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_rPort_12_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_12_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_12_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_12_backpressure; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_rPort_12_output_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_rPort_11_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_11_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_11_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_11_backpressure; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_rPort_11_output_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_rPort_10_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_10_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_10_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_10_backpressure; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_rPort_10_output_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_rPort_9_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_9_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_9_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_9_backpressure; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_rPort_9_output_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_rPort_8_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_8_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_8_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_8_backpressure; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_rPort_8_output_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_rPort_7_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_7_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_7_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_7_backpressure; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_rPort_7_output_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_rPort_6_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_6_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_6_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_6_backpressure; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_rPort_6_output_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_rPort_5_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_5_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_5_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_5_backpressure; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_rPort_5_output_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_rPort_4_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_4_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_4_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_4_backpressure; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_rPort_4_output_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_rPort_3_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_3_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_3_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_3_backpressure; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_rPort_3_output_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_rPort_2_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_2_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_2_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_2_backpressure; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_rPort_2_output_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_rPort_1_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_1_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_1_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_1_backpressure; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_rPort_1_output_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_rPort_0_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_0_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_0_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_rPort_0_backpressure; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_rPort_0_output_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_wPort_7_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_7_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_wPort_7_data_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_7_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_wPort_6_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_6_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_wPort_6_data_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_6_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_wPort_5_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_5_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_wPort_5_data_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_5_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_wPort_4_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_4_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_wPort_4_data_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_4_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_wPort_3_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_3_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_wPort_3_data_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_3_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_wPort_2_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_2_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_wPort_2_data_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_2_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_wPort_1_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_1_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_wPort_1_data_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_1_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [2:0] x525_lb2_0_io_wPort_0_banks_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_0_ofs_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire [7:0] x525_lb2_0_io_wPort_0_data_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  x525_lb2_0_io_wPort_0_en_0; // @[m_x525_lb2_0.scala 48:17:@45164.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@45336.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@45336.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@45336.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@45336.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@45336.4]
  wire  x539_sum_1_clock; // @[Math.scala 150:24:@45444.4]
  wire  x539_sum_1_reset; // @[Math.scala 150:24:@45444.4]
  wire [31:0] x539_sum_1_io_a; // @[Math.scala 150:24:@45444.4]
  wire [31:0] x539_sum_1_io_b; // @[Math.scala 150:24:@45444.4]
  wire  x539_sum_1_io_flow; // @[Math.scala 150:24:@45444.4]
  wire [31:0] x539_sum_1_io_result; // @[Math.scala 150:24:@45444.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@45454.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@45454.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@45454.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@45454.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@45454.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@45463.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@45463.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@45463.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@45463.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@45463.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@45472.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@45472.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@45472.4]
  wire [7:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@45472.4]
  wire [7:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@45472.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@45481.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@45481.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@45481.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@45481.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@45481.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@45490.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@45490.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@45490.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@45490.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@45490.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@45503.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@45503.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@45503.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@45503.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@45503.4]
  wire  x545_rdcol_1_clock; // @[Math.scala 150:24:@45526.4]
  wire  x545_rdcol_1_reset; // @[Math.scala 150:24:@45526.4]
  wire [31:0] x545_rdcol_1_io_a; // @[Math.scala 150:24:@45526.4]
  wire [31:0] x545_rdcol_1_io_b; // @[Math.scala 150:24:@45526.4]
  wire  x545_rdcol_1_io_flow; // @[Math.scala 150:24:@45526.4]
  wire [31:0] x545_rdcol_1_io_result; // @[Math.scala 150:24:@45526.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@45547.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@45547.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@45547.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@45547.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@45547.4]
  wire  x549_sum_1_clock; // @[Math.scala 150:24:@45556.4]
  wire  x549_sum_1_reset; // @[Math.scala 150:24:@45556.4]
  wire [31:0] x549_sum_1_io_a; // @[Math.scala 150:24:@45556.4]
  wire [31:0] x549_sum_1_io_b; // @[Math.scala 150:24:@45556.4]
  wire  x549_sum_1_io_flow; // @[Math.scala 150:24:@45556.4]
  wire [31:0] x549_sum_1_io_result; // @[Math.scala 150:24:@45556.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@45566.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@45566.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@45566.4]
  wire [7:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@45566.4]
  wire [7:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@45566.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@45575.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@45575.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@45575.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@45575.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@45575.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@45588.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@45588.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@45588.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@45588.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@45588.4]
  wire  x554_rdcol_1_clock; // @[Math.scala 150:24:@45611.4]
  wire  x554_rdcol_1_reset; // @[Math.scala 150:24:@45611.4]
  wire [31:0] x554_rdcol_1_io_a; // @[Math.scala 150:24:@45611.4]
  wire [31:0] x554_rdcol_1_io_b; // @[Math.scala 150:24:@45611.4]
  wire  x554_rdcol_1_io_flow; // @[Math.scala 150:24:@45611.4]
  wire [31:0] x554_rdcol_1_io_result; // @[Math.scala 150:24:@45611.4]
  wire  x558_sum_1_clock; // @[Math.scala 150:24:@45632.4]
  wire  x558_sum_1_reset; // @[Math.scala 150:24:@45632.4]
  wire [31:0] x558_sum_1_io_a; // @[Math.scala 150:24:@45632.4]
  wire [31:0] x558_sum_1_io_b; // @[Math.scala 150:24:@45632.4]
  wire  x558_sum_1_io_flow; // @[Math.scala 150:24:@45632.4]
  wire [31:0] x558_sum_1_io_result; // @[Math.scala 150:24:@45632.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@45642.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@45642.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@45642.4]
  wire [7:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@45642.4]
  wire [7:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@45642.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@45651.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@45651.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@45651.4]
  wire [31:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@45651.4]
  wire [31:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@45651.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@45664.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@45664.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@45664.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@45664.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@45664.4]
  wire  x563_rdcol_1_clock; // @[Math.scala 150:24:@45687.4]
  wire  x563_rdcol_1_reset; // @[Math.scala 150:24:@45687.4]
  wire [31:0] x563_rdcol_1_io_a; // @[Math.scala 150:24:@45687.4]
  wire [31:0] x563_rdcol_1_io_b; // @[Math.scala 150:24:@45687.4]
  wire  x563_rdcol_1_io_flow; // @[Math.scala 150:24:@45687.4]
  wire [31:0] x563_rdcol_1_io_result; // @[Math.scala 150:24:@45687.4]
  wire  x567_sum_1_clock; // @[Math.scala 150:24:@45708.4]
  wire  x567_sum_1_reset; // @[Math.scala 150:24:@45708.4]
  wire [31:0] x567_sum_1_io_a; // @[Math.scala 150:24:@45708.4]
  wire [31:0] x567_sum_1_io_b; // @[Math.scala 150:24:@45708.4]
  wire  x567_sum_1_io_flow; // @[Math.scala 150:24:@45708.4]
  wire [31:0] x567_sum_1_io_result; // @[Math.scala 150:24:@45708.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@45718.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@45718.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@45718.4]
  wire [31:0] RetimeWrapper_14_io_in; // @[package.scala 93:22:@45718.4]
  wire [31:0] RetimeWrapper_14_io_out; // @[package.scala 93:22:@45718.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@45727.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@45727.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@45727.4]
  wire [7:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@45727.4]
  wire [7:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@45727.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@45740.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@45740.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@45740.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@45740.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@45740.4]
  wire  x572_rdrow_1_clock; // @[Math.scala 150:24:@45763.4]
  wire  x572_rdrow_1_reset; // @[Math.scala 150:24:@45763.4]
  wire [31:0] x572_rdrow_1_io_a; // @[Math.scala 150:24:@45763.4]
  wire [31:0] x572_rdrow_1_io_b; // @[Math.scala 150:24:@45763.4]
  wire  x572_rdrow_1_io_flow; // @[Math.scala 150:24:@45763.4]
  wire [31:0] x572_rdrow_1_io_result; // @[Math.scala 150:24:@45763.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@45844.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@45844.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@45844.4]
  wire [31:0] RetimeWrapper_17_io_in; // @[package.scala 93:22:@45844.4]
  wire [31:0] RetimeWrapper_17_io_out; // @[package.scala 93:22:@45844.4]
  wire  x581_sum_1_clock; // @[Math.scala 150:24:@45853.4]
  wire  x581_sum_1_reset; // @[Math.scala 150:24:@45853.4]
  wire [31:0] x581_sum_1_io_a; // @[Math.scala 150:24:@45853.4]
  wire [31:0] x581_sum_1_io_b; // @[Math.scala 150:24:@45853.4]
  wire  x581_sum_1_io_flow; // @[Math.scala 150:24:@45853.4]
  wire [31:0] x581_sum_1_io_result; // @[Math.scala 150:24:@45853.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@45863.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@45863.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@45863.4]
  wire [7:0] RetimeWrapper_18_io_in; // @[package.scala 93:22:@45863.4]
  wire [7:0] RetimeWrapper_18_io_out; // @[package.scala 93:22:@45863.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@45872.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@45872.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@45872.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@45872.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@45872.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@45881.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@45881.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@45881.4]
  wire [31:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@45881.4]
  wire [31:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@45881.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@45894.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@45894.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@45894.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@45894.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@45894.4]
  wire  x587_sum_1_clock; // @[Math.scala 150:24:@45917.4]
  wire  x587_sum_1_reset; // @[Math.scala 150:24:@45917.4]
  wire [31:0] x587_sum_1_io_a; // @[Math.scala 150:24:@45917.4]
  wire [31:0] x587_sum_1_io_b; // @[Math.scala 150:24:@45917.4]
  wire  x587_sum_1_io_flow; // @[Math.scala 150:24:@45917.4]
  wire [31:0] x587_sum_1_io_result; // @[Math.scala 150:24:@45917.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@45927.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@45927.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@45927.4]
  wire [31:0] RetimeWrapper_22_io_in; // @[package.scala 93:22:@45927.4]
  wire [31:0] RetimeWrapper_22_io_out; // @[package.scala 93:22:@45927.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@45936.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@45936.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@45936.4]
  wire [7:0] RetimeWrapper_23_io_in; // @[package.scala 93:22:@45936.4]
  wire [7:0] RetimeWrapper_23_io_out; // @[package.scala 93:22:@45936.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@45949.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@45949.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@45949.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@45949.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@45949.4]
  wire  x592_sum_1_clock; // @[Math.scala 150:24:@45972.4]
  wire  x592_sum_1_reset; // @[Math.scala 150:24:@45972.4]
  wire [31:0] x592_sum_1_io_a; // @[Math.scala 150:24:@45972.4]
  wire [31:0] x592_sum_1_io_b; // @[Math.scala 150:24:@45972.4]
  wire  x592_sum_1_io_flow; // @[Math.scala 150:24:@45972.4]
  wire [31:0] x592_sum_1_io_result; // @[Math.scala 150:24:@45972.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@45982.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@45982.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@45982.4]
  wire [7:0] RetimeWrapper_25_io_in; // @[package.scala 93:22:@45982.4]
  wire [7:0] RetimeWrapper_25_io_out; // @[package.scala 93:22:@45982.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@45991.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@45991.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@45991.4]
  wire [31:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@45991.4]
  wire [31:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@45991.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@46004.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@46004.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@46004.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@46004.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@46004.4]
  wire  x597_sum_1_clock; // @[Math.scala 150:24:@46027.4]
  wire  x597_sum_1_reset; // @[Math.scala 150:24:@46027.4]
  wire [31:0] x597_sum_1_io_a; // @[Math.scala 150:24:@46027.4]
  wire [31:0] x597_sum_1_io_b; // @[Math.scala 150:24:@46027.4]
  wire  x597_sum_1_io_flow; // @[Math.scala 150:24:@46027.4]
  wire [31:0] x597_sum_1_io_result; // @[Math.scala 150:24:@46027.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@46037.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@46037.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@46037.4]
  wire [31:0] RetimeWrapper_28_io_in; // @[package.scala 93:22:@46037.4]
  wire [31:0] RetimeWrapper_28_io_out; // @[package.scala 93:22:@46037.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@46046.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@46046.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@46046.4]
  wire [7:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@46046.4]
  wire [7:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@46046.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@46059.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@46059.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@46059.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@46059.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@46059.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@46080.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@46080.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@46080.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@46080.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@46080.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@46107.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@46107.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@46107.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@46107.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@46107.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@46149.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@46149.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@46149.4]
  wire [31:0] RetimeWrapper_33_io_in; // @[package.scala 93:22:@46149.4]
  wire [31:0] RetimeWrapper_33_io_out; // @[package.scala 93:22:@46149.4]
  wire  x609_sum_1_clock; // @[Math.scala 150:24:@46158.4]
  wire  x609_sum_1_reset; // @[Math.scala 150:24:@46158.4]
  wire [31:0] x609_sum_1_io_a; // @[Math.scala 150:24:@46158.4]
  wire [31:0] x609_sum_1_io_b; // @[Math.scala 150:24:@46158.4]
  wire  x609_sum_1_io_flow; // @[Math.scala 150:24:@46158.4]
  wire [31:0] x609_sum_1_io_result; // @[Math.scala 150:24:@46158.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@46168.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@46168.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@46168.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@46168.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@46168.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@46177.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@46177.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@46177.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@46177.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@46177.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@46186.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@46186.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@46186.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@46186.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@46186.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@46195.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@46195.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@46195.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@46195.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@46195.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@46209.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@46209.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@46209.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@46209.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@46209.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@46230.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@46230.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@46230.4]
  wire [31:0] RetimeWrapper_39_io_in; // @[package.scala 93:22:@46230.4]
  wire [31:0] RetimeWrapper_39_io_out; // @[package.scala 93:22:@46230.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@46252.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@46252.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@46252.4]
  wire [31:0] RetimeWrapper_40_io_in; // @[package.scala 93:22:@46252.4]
  wire [31:0] RetimeWrapper_40_io_out; // @[package.scala 93:22:@46252.4]
  wire  x618_sum_1_clock; // @[Math.scala 150:24:@46261.4]
  wire  x618_sum_1_reset; // @[Math.scala 150:24:@46261.4]
  wire [31:0] x618_sum_1_io_a; // @[Math.scala 150:24:@46261.4]
  wire [31:0] x618_sum_1_io_b; // @[Math.scala 150:24:@46261.4]
  wire  x618_sum_1_io_flow; // @[Math.scala 150:24:@46261.4]
  wire [31:0] x618_sum_1_io_result; // @[Math.scala 150:24:@46261.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@46271.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@46271.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@46271.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@46271.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@46271.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@46285.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@46285.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@46285.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@46285.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@46285.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@46306.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@46306.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@46306.4]
  wire [31:0] RetimeWrapper_43_io_in; // @[package.scala 93:22:@46306.4]
  wire [31:0] RetimeWrapper_43_io_out; // @[package.scala 93:22:@46306.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@46330.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@46330.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@46330.4]
  wire [31:0] RetimeWrapper_44_io_in; // @[package.scala 93:22:@46330.4]
  wire [31:0] RetimeWrapper_44_io_out; // @[package.scala 93:22:@46330.4]
  wire  x626_sum_1_clock; // @[Math.scala 150:24:@46339.4]
  wire  x626_sum_1_reset; // @[Math.scala 150:24:@46339.4]
  wire [31:0] x626_sum_1_io_a; // @[Math.scala 150:24:@46339.4]
  wire [31:0] x626_sum_1_io_b; // @[Math.scala 150:24:@46339.4]
  wire  x626_sum_1_io_flow; // @[Math.scala 150:24:@46339.4]
  wire [31:0] x626_sum_1_io_result; // @[Math.scala 150:24:@46339.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@46349.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@46349.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@46349.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@46349.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@46349.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@46363.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@46363.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@46363.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@46363.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@46363.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@46384.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@46384.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@46384.4]
  wire [31:0] RetimeWrapper_47_io_in; // @[package.scala 93:22:@46384.4]
  wire [31:0] RetimeWrapper_47_io_out; // @[package.scala 93:22:@46384.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@46400.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@46400.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@46400.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@46400.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@46400.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@46415.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@46415.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@46415.4]
  wire [31:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@46415.4]
  wire [31:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@46415.4]
  wire  x634_sum_1_clock; // @[Math.scala 150:24:@46424.4]
  wire  x634_sum_1_reset; // @[Math.scala 150:24:@46424.4]
  wire [31:0] x634_sum_1_io_a; // @[Math.scala 150:24:@46424.4]
  wire [31:0] x634_sum_1_io_b; // @[Math.scala 150:24:@46424.4]
  wire  x634_sum_1_io_flow; // @[Math.scala 150:24:@46424.4]
  wire [31:0] x634_sum_1_io_result; // @[Math.scala 150:24:@46424.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@46434.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@46434.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@46434.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@46434.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@46434.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@46448.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@46448.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@46448.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@46448.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@46448.4]
  wire  x639_rdcol_1_clock; // @[Math.scala 150:24:@46471.4]
  wire  x639_rdcol_1_reset; // @[Math.scala 150:24:@46471.4]
  wire [31:0] x639_rdcol_1_io_a; // @[Math.scala 150:24:@46471.4]
  wire [31:0] x639_rdcol_1_io_b; // @[Math.scala 150:24:@46471.4]
  wire  x639_rdcol_1_io_flow; // @[Math.scala 150:24:@46471.4]
  wire [31:0] x639_rdcol_1_io_result; // @[Math.scala 150:24:@46471.4]
  wire  x645_sum_1_clock; // @[Math.scala 150:24:@46503.4]
  wire  x645_sum_1_reset; // @[Math.scala 150:24:@46503.4]
  wire [31:0] x645_sum_1_io_a; // @[Math.scala 150:24:@46503.4]
  wire [31:0] x645_sum_1_io_b; // @[Math.scala 150:24:@46503.4]
  wire  x645_sum_1_io_flow; // @[Math.scala 150:24:@46503.4]
  wire [31:0] x645_sum_1_io_result; // @[Math.scala 150:24:@46503.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@46513.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@46513.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@46513.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@46513.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@46513.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@46527.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@46527.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@46527.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@46527.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@46527.4]
  wire  x651_rdcol_1_clock; // @[Math.scala 150:24:@46550.4]
  wire  x651_rdcol_1_reset; // @[Math.scala 150:24:@46550.4]
  wire [31:0] x651_rdcol_1_io_a; // @[Math.scala 150:24:@46550.4]
  wire [31:0] x651_rdcol_1_io_b; // @[Math.scala 150:24:@46550.4]
  wire  x651_rdcol_1_io_flow; // @[Math.scala 150:24:@46550.4]
  wire [31:0] x651_rdcol_1_io_result; // @[Math.scala 150:24:@46550.4]
  wire  x657_sum_1_clock; // @[Math.scala 150:24:@46582.4]
  wire  x657_sum_1_reset; // @[Math.scala 150:24:@46582.4]
  wire [31:0] x657_sum_1_io_a; // @[Math.scala 150:24:@46582.4]
  wire [31:0] x657_sum_1_io_b; // @[Math.scala 150:24:@46582.4]
  wire  x657_sum_1_io_flow; // @[Math.scala 150:24:@46582.4]
  wire [31:0] x657_sum_1_io_result; // @[Math.scala 150:24:@46582.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@46592.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@46592.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@46592.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@46592.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@46592.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@46606.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@46606.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@46606.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@46606.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@46606.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@46627.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@46627.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@46627.4]
  wire [31:0] RetimeWrapper_56_io_in; // @[package.scala 93:22:@46627.4]
  wire [31:0] RetimeWrapper_56_io_out; // @[package.scala 93:22:@46627.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@46654.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@46654.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@46654.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@46654.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@46654.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@46689.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@46689.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@46689.4]
  wire [31:0] RetimeWrapper_58_io_in; // @[package.scala 93:22:@46689.4]
  wire [31:0] RetimeWrapper_58_io_out; // @[package.scala 93:22:@46689.4]
  wire  x669_sum_1_clock; // @[Math.scala 150:24:@46700.4]
  wire  x669_sum_1_reset; // @[Math.scala 150:24:@46700.4]
  wire [31:0] x669_sum_1_io_a; // @[Math.scala 150:24:@46700.4]
  wire [31:0] x669_sum_1_io_b; // @[Math.scala 150:24:@46700.4]
  wire  x669_sum_1_io_flow; // @[Math.scala 150:24:@46700.4]
  wire [31:0] x669_sum_1_io_result; // @[Math.scala 150:24:@46700.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@46710.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@46710.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@46710.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@46710.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@46710.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@46719.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@46719.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@46719.4]
  wire [31:0] RetimeWrapper_60_io_in; // @[package.scala 93:22:@46719.4]
  wire [31:0] RetimeWrapper_60_io_out; // @[package.scala 93:22:@46719.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@46733.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@46733.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@46733.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@46733.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@46733.4]
  wire  x677_sum_1_clock; // @[Math.scala 150:24:@46760.4]
  wire  x677_sum_1_reset; // @[Math.scala 150:24:@46760.4]
  wire [31:0] x677_sum_1_io_a; // @[Math.scala 150:24:@46760.4]
  wire [31:0] x677_sum_1_io_b; // @[Math.scala 150:24:@46760.4]
  wire  x677_sum_1_io_flow; // @[Math.scala 150:24:@46760.4]
  wire [31:0] x677_sum_1_io_result; // @[Math.scala 150:24:@46760.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@46770.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@46770.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@46770.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@46770.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@46770.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@46784.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@46784.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@46784.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@46784.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@46784.4]
  wire  x684_sum_1_clock; // @[Math.scala 150:24:@46811.4]
  wire  x684_sum_1_reset; // @[Math.scala 150:24:@46811.4]
  wire [31:0] x684_sum_1_io_a; // @[Math.scala 150:24:@46811.4]
  wire [31:0] x684_sum_1_io_b; // @[Math.scala 150:24:@46811.4]
  wire  x684_sum_1_io_flow; // @[Math.scala 150:24:@46811.4]
  wire [31:0] x684_sum_1_io_result; // @[Math.scala 150:24:@46811.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@46821.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@46821.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@46821.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@46821.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@46821.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@46835.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@46835.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@46835.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@46835.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@46835.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@46862.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@46862.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@46862.4]
  wire [31:0] RetimeWrapper_66_io_in; // @[package.scala 93:22:@46862.4]
  wire [31:0] RetimeWrapper_66_io_out; // @[package.scala 93:22:@46862.4]
  wire  x691_sum_1_clock; // @[Math.scala 150:24:@46871.4]
  wire  x691_sum_1_reset; // @[Math.scala 150:24:@46871.4]
  wire [31:0] x691_sum_1_io_a; // @[Math.scala 150:24:@46871.4]
  wire [31:0] x691_sum_1_io_b; // @[Math.scala 150:24:@46871.4]
  wire  x691_sum_1_io_flow; // @[Math.scala 150:24:@46871.4]
  wire [31:0] x691_sum_1_io_result; // @[Math.scala 150:24:@46871.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@46881.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@46881.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@46881.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@46881.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@46881.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@46890.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@46890.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@46890.4]
  wire [31:0] RetimeWrapper_68_io_in; // @[package.scala 93:22:@46890.4]
  wire [31:0] RetimeWrapper_68_io_out; // @[package.scala 93:22:@46890.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@46904.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@46904.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@46904.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@46904.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@46904.4]
  wire  x698_sum_1_clock; // @[Math.scala 150:24:@46931.4]
  wire  x698_sum_1_reset; // @[Math.scala 150:24:@46931.4]
  wire [31:0] x698_sum_1_io_a; // @[Math.scala 150:24:@46931.4]
  wire [31:0] x698_sum_1_io_b; // @[Math.scala 150:24:@46931.4]
  wire  x698_sum_1_io_flow; // @[Math.scala 150:24:@46931.4]
  wire [31:0] x698_sum_1_io_result; // @[Math.scala 150:24:@46931.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@46941.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@46941.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@46941.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@46941.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@46941.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@46955.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@46955.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@46955.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@46955.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@46955.4]
  wire  x705_sum_1_clock; // @[Math.scala 150:24:@46982.4]
  wire  x705_sum_1_reset; // @[Math.scala 150:24:@46982.4]
  wire [31:0] x705_sum_1_io_a; // @[Math.scala 150:24:@46982.4]
  wire [31:0] x705_sum_1_io_b; // @[Math.scala 150:24:@46982.4]
  wire  x705_sum_1_io_flow; // @[Math.scala 150:24:@46982.4]
  wire [31:0] x705_sum_1_io_result; // @[Math.scala 150:24:@46982.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@46992.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@46992.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@46992.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@46992.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@46992.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@47006.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@47006.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@47006.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@47006.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@47006.4]
  wire  x710_rdrow_1_clock; // @[Math.scala 150:24:@47029.4]
  wire  x710_rdrow_1_reset; // @[Math.scala 150:24:@47029.4]
  wire [31:0] x710_rdrow_1_io_a; // @[Math.scala 150:24:@47029.4]
  wire [31:0] x710_rdrow_1_io_b; // @[Math.scala 150:24:@47029.4]
  wire  x710_rdrow_1_io_flow; // @[Math.scala 150:24:@47029.4]
  wire [31:0] x710_rdrow_1_io_result; // @[Math.scala 150:24:@47029.4]
  wire  x717_sum_1_clock; // @[Math.scala 150:24:@47083.4]
  wire  x717_sum_1_reset; // @[Math.scala 150:24:@47083.4]
  wire [31:0] x717_sum_1_io_a; // @[Math.scala 150:24:@47083.4]
  wire [31:0] x717_sum_1_io_b; // @[Math.scala 150:24:@47083.4]
  wire  x717_sum_1_io_flow; // @[Math.scala 150:24:@47083.4]
  wire [31:0] x717_sum_1_io_result; // @[Math.scala 150:24:@47083.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@47093.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@47093.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@47093.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@47093.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@47093.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@47102.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@47102.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@47102.4]
  wire [31:0] RetimeWrapper_75_io_in; // @[package.scala 93:22:@47102.4]
  wire [31:0] RetimeWrapper_75_io_out; // @[package.scala 93:22:@47102.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@47116.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@47116.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@47116.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@47116.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@47116.4]
  wire  x725_sum_1_clock; // @[Math.scala 150:24:@47145.4]
  wire  x725_sum_1_reset; // @[Math.scala 150:24:@47145.4]
  wire [31:0] x725_sum_1_io_a; // @[Math.scala 150:24:@47145.4]
  wire [31:0] x725_sum_1_io_b; // @[Math.scala 150:24:@47145.4]
  wire  x725_sum_1_io_flow; // @[Math.scala 150:24:@47145.4]
  wire [31:0] x725_sum_1_io_result; // @[Math.scala 150:24:@47145.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@47155.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@47155.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@47155.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@47155.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@47155.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@47169.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@47169.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@47169.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@47169.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@47169.4]
  wire  x732_sum_1_clock; // @[Math.scala 150:24:@47196.4]
  wire  x732_sum_1_reset; // @[Math.scala 150:24:@47196.4]
  wire [31:0] x732_sum_1_io_a; // @[Math.scala 150:24:@47196.4]
  wire [31:0] x732_sum_1_io_b; // @[Math.scala 150:24:@47196.4]
  wire  x732_sum_1_io_flow; // @[Math.scala 150:24:@47196.4]
  wire [31:0] x732_sum_1_io_result; // @[Math.scala 150:24:@47196.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@47206.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@47206.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@47206.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@47206.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@47206.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@47220.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@47220.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@47220.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@47220.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@47220.4]
  wire  x739_sum_1_clock; // @[Math.scala 150:24:@47247.4]
  wire  x739_sum_1_reset; // @[Math.scala 150:24:@47247.4]
  wire [31:0] x739_sum_1_io_a; // @[Math.scala 150:24:@47247.4]
  wire [31:0] x739_sum_1_io_b; // @[Math.scala 150:24:@47247.4]
  wire  x739_sum_1_io_flow; // @[Math.scala 150:24:@47247.4]
  wire [31:0] x739_sum_1_io_result; // @[Math.scala 150:24:@47247.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@47257.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@47257.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@47257.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@47257.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@47257.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@47271.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@47271.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@47271.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@47271.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@47271.4]
  wire  x746_sum_1_clock; // @[Math.scala 150:24:@47298.4]
  wire  x746_sum_1_reset; // @[Math.scala 150:24:@47298.4]
  wire [31:0] x746_sum_1_io_a; // @[Math.scala 150:24:@47298.4]
  wire [31:0] x746_sum_1_io_b; // @[Math.scala 150:24:@47298.4]
  wire  x746_sum_1_io_flow; // @[Math.scala 150:24:@47298.4]
  wire [31:0] x746_sum_1_io_result; // @[Math.scala 150:24:@47298.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@47308.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@47308.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@47308.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@47308.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@47308.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@47322.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@47322.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@47322.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@47322.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@47322.4]
  wire  x753_sum_1_clock; // @[Math.scala 150:24:@47349.4]
  wire  x753_sum_1_reset; // @[Math.scala 150:24:@47349.4]
  wire [31:0] x753_sum_1_io_a; // @[Math.scala 150:24:@47349.4]
  wire [31:0] x753_sum_1_io_b; // @[Math.scala 150:24:@47349.4]
  wire  x753_sum_1_io_flow; // @[Math.scala 150:24:@47349.4]
  wire [31:0] x753_sum_1_io_result; // @[Math.scala 150:24:@47349.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@47359.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@47359.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@47359.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@47359.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@47359.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@47373.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@47373.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@47373.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@47373.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@47373.4]
  wire  x758_rdrow_1_clock; // @[Math.scala 150:24:@47396.4]
  wire  x758_rdrow_1_reset; // @[Math.scala 150:24:@47396.4]
  wire [31:0] x758_rdrow_1_io_a; // @[Math.scala 150:24:@47396.4]
  wire [31:0] x758_rdrow_1_io_b; // @[Math.scala 150:24:@47396.4]
  wire  x758_rdrow_1_io_flow; // @[Math.scala 150:24:@47396.4]
  wire [31:0] x758_rdrow_1_io_result; // @[Math.scala 150:24:@47396.4]
  wire  x765_sum_1_clock; // @[Math.scala 150:24:@47450.4]
  wire  x765_sum_1_reset; // @[Math.scala 150:24:@47450.4]
  wire [31:0] x765_sum_1_io_a; // @[Math.scala 150:24:@47450.4]
  wire [31:0] x765_sum_1_io_b; // @[Math.scala 150:24:@47450.4]
  wire  x765_sum_1_io_flow; // @[Math.scala 150:24:@47450.4]
  wire [31:0] x765_sum_1_io_result; // @[Math.scala 150:24:@47450.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@47460.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@47460.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@47460.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@47460.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@47460.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@47469.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@47469.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@47469.4]
  wire [31:0] RetimeWrapper_88_io_in; // @[package.scala 93:22:@47469.4]
  wire [31:0] RetimeWrapper_88_io_out; // @[package.scala 93:22:@47469.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@47483.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@47483.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@47483.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@47483.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@47483.4]
  wire  x773_sum_1_clock; // @[Math.scala 150:24:@47510.4]
  wire  x773_sum_1_reset; // @[Math.scala 150:24:@47510.4]
  wire [31:0] x773_sum_1_io_a; // @[Math.scala 150:24:@47510.4]
  wire [31:0] x773_sum_1_io_b; // @[Math.scala 150:24:@47510.4]
  wire  x773_sum_1_io_flow; // @[Math.scala 150:24:@47510.4]
  wire [31:0] x773_sum_1_io_result; // @[Math.scala 150:24:@47510.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@47520.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@47520.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@47520.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@47520.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@47520.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@47534.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@47534.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@47534.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@47534.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@47534.4]
  wire  x780_sum_1_clock; // @[Math.scala 150:24:@47563.4]
  wire  x780_sum_1_reset; // @[Math.scala 150:24:@47563.4]
  wire [31:0] x780_sum_1_io_a; // @[Math.scala 150:24:@47563.4]
  wire [31:0] x780_sum_1_io_b; // @[Math.scala 150:24:@47563.4]
  wire  x780_sum_1_io_flow; // @[Math.scala 150:24:@47563.4]
  wire [31:0] x780_sum_1_io_result; // @[Math.scala 150:24:@47563.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@47573.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@47573.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@47573.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@47573.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@47573.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@47587.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@47587.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@47587.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@47587.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@47587.4]
  wire  x787_sum_1_clock; // @[Math.scala 150:24:@47614.4]
  wire  x787_sum_1_reset; // @[Math.scala 150:24:@47614.4]
  wire [31:0] x787_sum_1_io_a; // @[Math.scala 150:24:@47614.4]
  wire [31:0] x787_sum_1_io_b; // @[Math.scala 150:24:@47614.4]
  wire  x787_sum_1_io_flow; // @[Math.scala 150:24:@47614.4]
  wire [31:0] x787_sum_1_io_result; // @[Math.scala 150:24:@47614.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@47624.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@47624.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@47624.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@47624.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@47624.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@47638.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@47638.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@47638.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@47638.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@47638.4]
  wire  x794_sum_1_clock; // @[Math.scala 150:24:@47665.4]
  wire  x794_sum_1_reset; // @[Math.scala 150:24:@47665.4]
  wire [31:0] x794_sum_1_io_a; // @[Math.scala 150:24:@47665.4]
  wire [31:0] x794_sum_1_io_b; // @[Math.scala 150:24:@47665.4]
  wire  x794_sum_1_io_flow; // @[Math.scala 150:24:@47665.4]
  wire [31:0] x794_sum_1_io_result; // @[Math.scala 150:24:@47665.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@47675.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@47675.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@47675.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@47675.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@47675.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@47689.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@47689.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@47689.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@47689.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@47689.4]
  wire  x801_sum_1_clock; // @[Math.scala 150:24:@47716.4]
  wire  x801_sum_1_reset; // @[Math.scala 150:24:@47716.4]
  wire [31:0] x801_sum_1_io_a; // @[Math.scala 150:24:@47716.4]
  wire [31:0] x801_sum_1_io_b; // @[Math.scala 150:24:@47716.4]
  wire  x801_sum_1_io_flow; // @[Math.scala 150:24:@47716.4]
  wire [31:0] x801_sum_1_io_result; // @[Math.scala 150:24:@47716.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@47726.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@47726.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@47726.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@47726.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@47726.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@47740.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@47740.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@47740.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@47740.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@47740.4]
  wire  x811_x23_1_clock; // @[Math.scala 150:24:@47786.4]
  wire  x811_x23_1_reset; // @[Math.scala 150:24:@47786.4]
  wire [7:0] x811_x23_1_io_a; // @[Math.scala 150:24:@47786.4]
  wire [7:0] x811_x23_1_io_b; // @[Math.scala 150:24:@47786.4]
  wire  x811_x23_1_io_flow; // @[Math.scala 150:24:@47786.4]
  wire [7:0] x811_x23_1_io_result; // @[Math.scala 150:24:@47786.4]
  wire  x812_x24_1_clock; // @[Math.scala 150:24:@47796.4]
  wire  x812_x24_1_reset; // @[Math.scala 150:24:@47796.4]
  wire [7:0] x812_x24_1_io_a; // @[Math.scala 150:24:@47796.4]
  wire [7:0] x812_x24_1_io_b; // @[Math.scala 150:24:@47796.4]
  wire  x812_x24_1_io_flow; // @[Math.scala 150:24:@47796.4]
  wire [7:0] x812_x24_1_io_result; // @[Math.scala 150:24:@47796.4]
  wire  x813_x23_1_clock; // @[Math.scala 150:24:@47806.4]
  wire  x813_x23_1_reset; // @[Math.scala 150:24:@47806.4]
  wire [7:0] x813_x23_1_io_a; // @[Math.scala 150:24:@47806.4]
  wire [7:0] x813_x23_1_io_b; // @[Math.scala 150:24:@47806.4]
  wire  x813_x23_1_io_flow; // @[Math.scala 150:24:@47806.4]
  wire [7:0] x813_x23_1_io_result; // @[Math.scala 150:24:@47806.4]
  wire  x814_x24_1_clock; // @[Math.scala 150:24:@47816.4]
  wire  x814_x24_1_reset; // @[Math.scala 150:24:@47816.4]
  wire [7:0] x814_x24_1_io_a; // @[Math.scala 150:24:@47816.4]
  wire [7:0] x814_x24_1_io_b; // @[Math.scala 150:24:@47816.4]
  wire  x814_x24_1_io_flow; // @[Math.scala 150:24:@47816.4]
  wire [7:0] x814_x24_1_io_result; // @[Math.scala 150:24:@47816.4]
  wire [7:0] x815_x23_1_io_a; // @[Math.scala 150:24:@47826.4]
  wire [7:0] x815_x23_1_io_b; // @[Math.scala 150:24:@47826.4]
  wire [7:0] x815_x23_1_io_result; // @[Math.scala 150:24:@47826.4]
  wire [7:0] x816_x24_1_io_a; // @[Math.scala 150:24:@47836.4]
  wire [7:0] x816_x24_1_io_b; // @[Math.scala 150:24:@47836.4]
  wire [7:0] x816_x24_1_io_result; // @[Math.scala 150:24:@47836.4]
  wire [7:0] x817_x23_1_io_a; // @[Math.scala 150:24:@47846.4]
  wire [7:0] x817_x23_1_io_b; // @[Math.scala 150:24:@47846.4]
  wire [7:0] x817_x23_1_io_result; // @[Math.scala 150:24:@47846.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@47856.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@47856.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@47856.4]
  wire [7:0] RetimeWrapper_100_io_in; // @[package.scala 93:22:@47856.4]
  wire [7:0] RetimeWrapper_100_io_out; // @[package.scala 93:22:@47856.4]
  wire [7:0] x818_sum_1_io_a; // @[Math.scala 150:24:@47865.4]
  wire [7:0] x818_sum_1_io_b; // @[Math.scala 150:24:@47865.4]
  wire [7:0] x818_sum_1_io_result; // @[Math.scala 150:24:@47865.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@47879.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@47879.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@47879.4]
  wire [7:0] RetimeWrapper_101_io_in; // @[package.scala 93:22:@47879.4]
  wire [7:0] RetimeWrapper_101_io_out; // @[package.scala 93:22:@47879.4]
  wire  x825_x23_1_clock; // @[Math.scala 150:24:@47914.4]
  wire  x825_x23_1_reset; // @[Math.scala 150:24:@47914.4]
  wire [7:0] x825_x23_1_io_a; // @[Math.scala 150:24:@47914.4]
  wire [7:0] x825_x23_1_io_b; // @[Math.scala 150:24:@47914.4]
  wire  x825_x23_1_io_flow; // @[Math.scala 150:24:@47914.4]
  wire [7:0] x825_x23_1_io_result; // @[Math.scala 150:24:@47914.4]
  wire  x826_x24_1_clock; // @[Math.scala 150:24:@47924.4]
  wire  x826_x24_1_reset; // @[Math.scala 150:24:@47924.4]
  wire [7:0] x826_x24_1_io_a; // @[Math.scala 150:24:@47924.4]
  wire [7:0] x826_x24_1_io_b; // @[Math.scala 150:24:@47924.4]
  wire  x826_x24_1_io_flow; // @[Math.scala 150:24:@47924.4]
  wire [7:0] x826_x24_1_io_result; // @[Math.scala 150:24:@47924.4]
  wire  x827_x23_1_clock; // @[Math.scala 150:24:@47934.4]
  wire  x827_x23_1_reset; // @[Math.scala 150:24:@47934.4]
  wire [7:0] x827_x23_1_io_a; // @[Math.scala 150:24:@47934.4]
  wire [7:0] x827_x23_1_io_b; // @[Math.scala 150:24:@47934.4]
  wire  x827_x23_1_io_flow; // @[Math.scala 150:24:@47934.4]
  wire [7:0] x827_x23_1_io_result; // @[Math.scala 150:24:@47934.4]
  wire  x828_x24_1_clock; // @[Math.scala 150:24:@47944.4]
  wire  x828_x24_1_reset; // @[Math.scala 150:24:@47944.4]
  wire [7:0] x828_x24_1_io_a; // @[Math.scala 150:24:@47944.4]
  wire [7:0] x828_x24_1_io_b; // @[Math.scala 150:24:@47944.4]
  wire  x828_x24_1_io_flow; // @[Math.scala 150:24:@47944.4]
  wire [7:0] x828_x24_1_io_result; // @[Math.scala 150:24:@47944.4]
  wire [7:0] x829_x23_1_io_a; // @[Math.scala 150:24:@47954.4]
  wire [7:0] x829_x23_1_io_b; // @[Math.scala 150:24:@47954.4]
  wire [7:0] x829_x23_1_io_result; // @[Math.scala 150:24:@47954.4]
  wire [7:0] x830_x24_1_io_a; // @[Math.scala 150:24:@47964.4]
  wire [7:0] x830_x24_1_io_b; // @[Math.scala 150:24:@47964.4]
  wire [7:0] x830_x24_1_io_result; // @[Math.scala 150:24:@47964.4]
  wire [7:0] x831_x23_1_io_a; // @[Math.scala 150:24:@47976.4]
  wire [7:0] x831_x23_1_io_b; // @[Math.scala 150:24:@47976.4]
  wire [7:0] x831_x23_1_io_result; // @[Math.scala 150:24:@47976.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@47986.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@47986.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@47986.4]
  wire [7:0] RetimeWrapper_102_io_in; // @[package.scala 93:22:@47986.4]
  wire [7:0] RetimeWrapper_102_io_out; // @[package.scala 93:22:@47986.4]
  wire [7:0] x832_sum_1_io_a; // @[Math.scala 150:24:@47995.4]
  wire [7:0] x832_sum_1_io_b; // @[Math.scala 150:24:@47995.4]
  wire [7:0] x832_sum_1_io_result; // @[Math.scala 150:24:@47995.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@48009.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@48009.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@48009.4]
  wire [7:0] RetimeWrapper_103_io_in; // @[package.scala 93:22:@48009.4]
  wire [7:0] RetimeWrapper_103_io_out; // @[package.scala 93:22:@48009.4]
  wire  x838_x23_1_clock; // @[Math.scala 150:24:@48039.4]
  wire  x838_x23_1_reset; // @[Math.scala 150:24:@48039.4]
  wire [7:0] x838_x23_1_io_a; // @[Math.scala 150:24:@48039.4]
  wire [7:0] x838_x23_1_io_b; // @[Math.scala 150:24:@48039.4]
  wire  x838_x23_1_io_flow; // @[Math.scala 150:24:@48039.4]
  wire [7:0] x838_x23_1_io_result; // @[Math.scala 150:24:@48039.4]
  wire  x839_x24_1_clock; // @[Math.scala 150:24:@48049.4]
  wire  x839_x24_1_reset; // @[Math.scala 150:24:@48049.4]
  wire [7:0] x839_x24_1_io_a; // @[Math.scala 150:24:@48049.4]
  wire [7:0] x839_x24_1_io_b; // @[Math.scala 150:24:@48049.4]
  wire  x839_x24_1_io_flow; // @[Math.scala 150:24:@48049.4]
  wire [7:0] x839_x24_1_io_result; // @[Math.scala 150:24:@48049.4]
  wire  x840_x23_1_clock; // @[Math.scala 150:24:@48059.4]
  wire  x840_x23_1_reset; // @[Math.scala 150:24:@48059.4]
  wire [7:0] x840_x23_1_io_a; // @[Math.scala 150:24:@48059.4]
  wire [7:0] x840_x23_1_io_b; // @[Math.scala 150:24:@48059.4]
  wire  x840_x23_1_io_flow; // @[Math.scala 150:24:@48059.4]
  wire [7:0] x840_x23_1_io_result; // @[Math.scala 150:24:@48059.4]
  wire  x841_x24_1_clock; // @[Math.scala 150:24:@48069.4]
  wire  x841_x24_1_reset; // @[Math.scala 150:24:@48069.4]
  wire [7:0] x841_x24_1_io_a; // @[Math.scala 150:24:@48069.4]
  wire [7:0] x841_x24_1_io_b; // @[Math.scala 150:24:@48069.4]
  wire  x841_x24_1_io_flow; // @[Math.scala 150:24:@48069.4]
  wire [7:0] x841_x24_1_io_result; // @[Math.scala 150:24:@48069.4]
  wire [7:0] x842_x23_1_io_a; // @[Math.scala 150:24:@48079.4]
  wire [7:0] x842_x23_1_io_b; // @[Math.scala 150:24:@48079.4]
  wire [7:0] x842_x23_1_io_result; // @[Math.scala 150:24:@48079.4]
  wire [7:0] x843_x24_1_io_a; // @[Math.scala 150:24:@48089.4]
  wire [7:0] x843_x24_1_io_b; // @[Math.scala 150:24:@48089.4]
  wire [7:0] x843_x24_1_io_result; // @[Math.scala 150:24:@48089.4]
  wire [7:0] x844_x23_1_io_a; // @[Math.scala 150:24:@48099.4]
  wire [7:0] x844_x23_1_io_b; // @[Math.scala 150:24:@48099.4]
  wire [7:0] x844_x23_1_io_result; // @[Math.scala 150:24:@48099.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@48109.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@48109.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@48109.4]
  wire [7:0] RetimeWrapper_104_io_in; // @[package.scala 93:22:@48109.4]
  wire [7:0] RetimeWrapper_104_io_out; // @[package.scala 93:22:@48109.4]
  wire [7:0] x845_sum_1_io_a; // @[Math.scala 150:24:@48118.4]
  wire [7:0] x845_sum_1_io_b; // @[Math.scala 150:24:@48118.4]
  wire [7:0] x845_sum_1_io_result; // @[Math.scala 150:24:@48118.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@48132.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@48132.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@48132.4]
  wire [7:0] RetimeWrapper_105_io_in; // @[package.scala 93:22:@48132.4]
  wire [7:0] RetimeWrapper_105_io_out; // @[package.scala 93:22:@48132.4]
  wire  x851_x23_1_clock; // @[Math.scala 150:24:@48162.4]
  wire  x851_x23_1_reset; // @[Math.scala 150:24:@48162.4]
  wire [7:0] x851_x23_1_io_a; // @[Math.scala 150:24:@48162.4]
  wire [7:0] x851_x23_1_io_b; // @[Math.scala 150:24:@48162.4]
  wire  x851_x23_1_io_flow; // @[Math.scala 150:24:@48162.4]
  wire [7:0] x851_x23_1_io_result; // @[Math.scala 150:24:@48162.4]
  wire  x852_x24_1_clock; // @[Math.scala 150:24:@48172.4]
  wire  x852_x24_1_reset; // @[Math.scala 150:24:@48172.4]
  wire [7:0] x852_x24_1_io_a; // @[Math.scala 150:24:@48172.4]
  wire [7:0] x852_x24_1_io_b; // @[Math.scala 150:24:@48172.4]
  wire  x852_x24_1_io_flow; // @[Math.scala 150:24:@48172.4]
  wire [7:0] x852_x24_1_io_result; // @[Math.scala 150:24:@48172.4]
  wire  x853_x23_1_clock; // @[Math.scala 150:24:@48182.4]
  wire  x853_x23_1_reset; // @[Math.scala 150:24:@48182.4]
  wire [7:0] x853_x23_1_io_a; // @[Math.scala 150:24:@48182.4]
  wire [7:0] x853_x23_1_io_b; // @[Math.scala 150:24:@48182.4]
  wire  x853_x23_1_io_flow; // @[Math.scala 150:24:@48182.4]
  wire [7:0] x853_x23_1_io_result; // @[Math.scala 150:24:@48182.4]
  wire  x854_x24_1_clock; // @[Math.scala 150:24:@48192.4]
  wire  x854_x24_1_reset; // @[Math.scala 150:24:@48192.4]
  wire [7:0] x854_x24_1_io_a; // @[Math.scala 150:24:@48192.4]
  wire [7:0] x854_x24_1_io_b; // @[Math.scala 150:24:@48192.4]
  wire  x854_x24_1_io_flow; // @[Math.scala 150:24:@48192.4]
  wire [7:0] x854_x24_1_io_result; // @[Math.scala 150:24:@48192.4]
  wire [7:0] x855_x23_1_io_a; // @[Math.scala 150:24:@48202.4]
  wire [7:0] x855_x23_1_io_b; // @[Math.scala 150:24:@48202.4]
  wire [7:0] x855_x23_1_io_result; // @[Math.scala 150:24:@48202.4]
  wire [7:0] x856_x24_1_io_a; // @[Math.scala 150:24:@48212.4]
  wire [7:0] x856_x24_1_io_b; // @[Math.scala 150:24:@48212.4]
  wire [7:0] x856_x24_1_io_result; // @[Math.scala 150:24:@48212.4]
  wire [7:0] x857_x23_1_io_a; // @[Math.scala 150:24:@48222.4]
  wire [7:0] x857_x23_1_io_b; // @[Math.scala 150:24:@48222.4]
  wire [7:0] x857_x23_1_io_result; // @[Math.scala 150:24:@48222.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@48232.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@48232.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@48232.4]
  wire [7:0] RetimeWrapper_106_io_in; // @[package.scala 93:22:@48232.4]
  wire [7:0] RetimeWrapper_106_io_out; // @[package.scala 93:22:@48232.4]
  wire [7:0] x858_sum_1_io_a; // @[Math.scala 150:24:@48241.4]
  wire [7:0] x858_sum_1_io_b; // @[Math.scala 150:24:@48241.4]
  wire [7:0] x858_sum_1_io_result; // @[Math.scala 150:24:@48241.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@48255.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@48255.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@48255.4]
  wire [7:0] RetimeWrapper_107_io_in; // @[package.scala 93:22:@48255.4]
  wire [7:0] RetimeWrapper_107_io_out; // @[package.scala 93:22:@48255.4]
  wire  x863_x23_1_clock; // @[Math.scala 150:24:@48280.4]
  wire  x863_x23_1_reset; // @[Math.scala 150:24:@48280.4]
  wire [7:0] x863_x23_1_io_a; // @[Math.scala 150:24:@48280.4]
  wire [7:0] x863_x23_1_io_b; // @[Math.scala 150:24:@48280.4]
  wire  x863_x23_1_io_flow; // @[Math.scala 150:24:@48280.4]
  wire [7:0] x863_x23_1_io_result; // @[Math.scala 150:24:@48280.4]
  wire  x864_x24_1_clock; // @[Math.scala 150:24:@48290.4]
  wire  x864_x24_1_reset; // @[Math.scala 150:24:@48290.4]
  wire [7:0] x864_x24_1_io_a; // @[Math.scala 150:24:@48290.4]
  wire [7:0] x864_x24_1_io_b; // @[Math.scala 150:24:@48290.4]
  wire  x864_x24_1_io_flow; // @[Math.scala 150:24:@48290.4]
  wire [7:0] x864_x24_1_io_result; // @[Math.scala 150:24:@48290.4]
  wire  x865_x23_1_clock; // @[Math.scala 150:24:@48300.4]
  wire  x865_x23_1_reset; // @[Math.scala 150:24:@48300.4]
  wire [7:0] x865_x23_1_io_a; // @[Math.scala 150:24:@48300.4]
  wire [7:0] x865_x23_1_io_b; // @[Math.scala 150:24:@48300.4]
  wire  x865_x23_1_io_flow; // @[Math.scala 150:24:@48300.4]
  wire [7:0] x865_x23_1_io_result; // @[Math.scala 150:24:@48300.4]
  wire  x866_x24_1_clock; // @[Math.scala 150:24:@48310.4]
  wire  x866_x24_1_reset; // @[Math.scala 150:24:@48310.4]
  wire [7:0] x866_x24_1_io_a; // @[Math.scala 150:24:@48310.4]
  wire [7:0] x866_x24_1_io_b; // @[Math.scala 150:24:@48310.4]
  wire  x866_x24_1_io_flow; // @[Math.scala 150:24:@48310.4]
  wire [7:0] x866_x24_1_io_result; // @[Math.scala 150:24:@48310.4]
  wire [7:0] x867_x23_1_io_a; // @[Math.scala 150:24:@48320.4]
  wire [7:0] x867_x23_1_io_b; // @[Math.scala 150:24:@48320.4]
  wire [7:0] x867_x23_1_io_result; // @[Math.scala 150:24:@48320.4]
  wire [7:0] x868_x24_1_io_a; // @[Math.scala 150:24:@48330.4]
  wire [7:0] x868_x24_1_io_b; // @[Math.scala 150:24:@48330.4]
  wire [7:0] x868_x24_1_io_result; // @[Math.scala 150:24:@48330.4]
  wire [7:0] x869_x23_1_io_a; // @[Math.scala 150:24:@48340.4]
  wire [7:0] x869_x23_1_io_b; // @[Math.scala 150:24:@48340.4]
  wire [7:0] x869_x23_1_io_result; // @[Math.scala 150:24:@48340.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@48350.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@48350.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@48350.4]
  wire [7:0] RetimeWrapper_108_io_in; // @[package.scala 93:22:@48350.4]
  wire [7:0] RetimeWrapper_108_io_out; // @[package.scala 93:22:@48350.4]
  wire [7:0] x870_sum_1_io_a; // @[Math.scala 150:24:@48359.4]
  wire [7:0] x870_sum_1_io_b; // @[Math.scala 150:24:@48359.4]
  wire [7:0] x870_sum_1_io_result; // @[Math.scala 150:24:@48359.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@48373.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@48373.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@48373.4]
  wire [7:0] RetimeWrapper_109_io_in; // @[package.scala 93:22:@48373.4]
  wire [7:0] RetimeWrapper_109_io_out; // @[package.scala 93:22:@48373.4]
  wire  x874_x23_1_clock; // @[Math.scala 150:24:@48393.4]
  wire  x874_x23_1_reset; // @[Math.scala 150:24:@48393.4]
  wire [7:0] x874_x23_1_io_a; // @[Math.scala 150:24:@48393.4]
  wire [7:0] x874_x23_1_io_b; // @[Math.scala 150:24:@48393.4]
  wire  x874_x23_1_io_flow; // @[Math.scala 150:24:@48393.4]
  wire [7:0] x874_x23_1_io_result; // @[Math.scala 150:24:@48393.4]
  wire  x875_x24_1_clock; // @[Math.scala 150:24:@48403.4]
  wire  x875_x24_1_reset; // @[Math.scala 150:24:@48403.4]
  wire [7:0] x875_x24_1_io_a; // @[Math.scala 150:24:@48403.4]
  wire [7:0] x875_x24_1_io_b; // @[Math.scala 150:24:@48403.4]
  wire  x875_x24_1_io_flow; // @[Math.scala 150:24:@48403.4]
  wire [7:0] x875_x24_1_io_result; // @[Math.scala 150:24:@48403.4]
  wire  x876_x23_1_clock; // @[Math.scala 150:24:@48415.4]
  wire  x876_x23_1_reset; // @[Math.scala 150:24:@48415.4]
  wire [7:0] x876_x23_1_io_a; // @[Math.scala 150:24:@48415.4]
  wire [7:0] x876_x23_1_io_b; // @[Math.scala 150:24:@48415.4]
  wire  x876_x23_1_io_flow; // @[Math.scala 150:24:@48415.4]
  wire [7:0] x876_x23_1_io_result; // @[Math.scala 150:24:@48415.4]
  wire  x877_x24_1_clock; // @[Math.scala 150:24:@48425.4]
  wire  x877_x24_1_reset; // @[Math.scala 150:24:@48425.4]
  wire [7:0] x877_x24_1_io_a; // @[Math.scala 150:24:@48425.4]
  wire [7:0] x877_x24_1_io_b; // @[Math.scala 150:24:@48425.4]
  wire  x877_x24_1_io_flow; // @[Math.scala 150:24:@48425.4]
  wire [7:0] x877_x24_1_io_result; // @[Math.scala 150:24:@48425.4]
  wire [7:0] x878_x23_1_io_a; // @[Math.scala 150:24:@48435.4]
  wire [7:0] x878_x23_1_io_b; // @[Math.scala 150:24:@48435.4]
  wire [7:0] x878_x23_1_io_result; // @[Math.scala 150:24:@48435.4]
  wire [7:0] x879_x24_1_io_a; // @[Math.scala 150:24:@48445.4]
  wire [7:0] x879_x24_1_io_b; // @[Math.scala 150:24:@48445.4]
  wire [7:0] x879_x24_1_io_result; // @[Math.scala 150:24:@48445.4]
  wire [7:0] x880_x23_1_io_a; // @[Math.scala 150:24:@48455.4]
  wire [7:0] x880_x23_1_io_b; // @[Math.scala 150:24:@48455.4]
  wire [7:0] x880_x23_1_io_result; // @[Math.scala 150:24:@48455.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@48465.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@48465.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@48465.4]
  wire [7:0] RetimeWrapper_110_io_in; // @[package.scala 93:22:@48465.4]
  wire [7:0] RetimeWrapper_110_io_out; // @[package.scala 93:22:@48465.4]
  wire [7:0] x881_sum_1_io_a; // @[Math.scala 150:24:@48474.4]
  wire [7:0] x881_sum_1_io_b; // @[Math.scala 150:24:@48474.4]
  wire [7:0] x881_sum_1_io_result; // @[Math.scala 150:24:@48474.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@48488.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@48488.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@48488.4]
  wire [7:0] RetimeWrapper_111_io_in; // @[package.scala 93:22:@48488.4]
  wire [7:0] RetimeWrapper_111_io_out; // @[package.scala 93:22:@48488.4]
  wire  x885_x23_1_clock; // @[Math.scala 150:24:@48508.4]
  wire  x885_x23_1_reset; // @[Math.scala 150:24:@48508.4]
  wire [7:0] x885_x23_1_io_a; // @[Math.scala 150:24:@48508.4]
  wire [7:0] x885_x23_1_io_b; // @[Math.scala 150:24:@48508.4]
  wire  x885_x23_1_io_flow; // @[Math.scala 150:24:@48508.4]
  wire [7:0] x885_x23_1_io_result; // @[Math.scala 150:24:@48508.4]
  wire  x886_x24_1_clock; // @[Math.scala 150:24:@48518.4]
  wire  x886_x24_1_reset; // @[Math.scala 150:24:@48518.4]
  wire [7:0] x886_x24_1_io_a; // @[Math.scala 150:24:@48518.4]
  wire [7:0] x886_x24_1_io_b; // @[Math.scala 150:24:@48518.4]
  wire  x886_x24_1_io_flow; // @[Math.scala 150:24:@48518.4]
  wire [7:0] x886_x24_1_io_result; // @[Math.scala 150:24:@48518.4]
  wire  x887_x23_1_clock; // @[Math.scala 150:24:@48528.4]
  wire  x887_x23_1_reset; // @[Math.scala 150:24:@48528.4]
  wire [7:0] x887_x23_1_io_a; // @[Math.scala 150:24:@48528.4]
  wire [7:0] x887_x23_1_io_b; // @[Math.scala 150:24:@48528.4]
  wire  x887_x23_1_io_flow; // @[Math.scala 150:24:@48528.4]
  wire [7:0] x887_x23_1_io_result; // @[Math.scala 150:24:@48528.4]
  wire  x888_x24_1_clock; // @[Math.scala 150:24:@48538.4]
  wire  x888_x24_1_reset; // @[Math.scala 150:24:@48538.4]
  wire [7:0] x888_x24_1_io_a; // @[Math.scala 150:24:@48538.4]
  wire [7:0] x888_x24_1_io_b; // @[Math.scala 150:24:@48538.4]
  wire  x888_x24_1_io_flow; // @[Math.scala 150:24:@48538.4]
  wire [7:0] x888_x24_1_io_result; // @[Math.scala 150:24:@48538.4]
  wire [7:0] x889_x23_1_io_a; // @[Math.scala 150:24:@48548.4]
  wire [7:0] x889_x23_1_io_b; // @[Math.scala 150:24:@48548.4]
  wire [7:0] x889_x23_1_io_result; // @[Math.scala 150:24:@48548.4]
  wire [7:0] x890_x24_1_io_a; // @[Math.scala 150:24:@48558.4]
  wire [7:0] x890_x24_1_io_b; // @[Math.scala 150:24:@48558.4]
  wire [7:0] x890_x24_1_io_result; // @[Math.scala 150:24:@48558.4]
  wire [7:0] x891_x23_1_io_a; // @[Math.scala 150:24:@48568.4]
  wire [7:0] x891_x23_1_io_b; // @[Math.scala 150:24:@48568.4]
  wire [7:0] x891_x23_1_io_result; // @[Math.scala 150:24:@48568.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@48578.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@48578.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@48578.4]
  wire [7:0] RetimeWrapper_112_io_in; // @[package.scala 93:22:@48578.4]
  wire [7:0] RetimeWrapper_112_io_out; // @[package.scala 93:22:@48578.4]
  wire [7:0] x892_sum_1_io_a; // @[Math.scala 150:24:@48587.4]
  wire [7:0] x892_sum_1_io_b; // @[Math.scala 150:24:@48587.4]
  wire [7:0] x892_sum_1_io_result; // @[Math.scala 150:24:@48587.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@48601.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@48601.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@48601.4]
  wire [7:0] RetimeWrapper_113_io_in; // @[package.scala 93:22:@48601.4]
  wire [7:0] RetimeWrapper_113_io_out; // @[package.scala 93:22:@48601.4]
  wire  x897_x23_1_clock; // @[Math.scala 150:24:@48626.4]
  wire  x897_x23_1_reset; // @[Math.scala 150:24:@48626.4]
  wire [7:0] x897_x23_1_io_a; // @[Math.scala 150:24:@48626.4]
  wire [7:0] x897_x23_1_io_b; // @[Math.scala 150:24:@48626.4]
  wire  x897_x23_1_io_flow; // @[Math.scala 150:24:@48626.4]
  wire [7:0] x897_x23_1_io_result; // @[Math.scala 150:24:@48626.4]
  wire  x898_x24_1_clock; // @[Math.scala 150:24:@48636.4]
  wire  x898_x24_1_reset; // @[Math.scala 150:24:@48636.4]
  wire [7:0] x898_x24_1_io_a; // @[Math.scala 150:24:@48636.4]
  wire [7:0] x898_x24_1_io_b; // @[Math.scala 150:24:@48636.4]
  wire  x898_x24_1_io_flow; // @[Math.scala 150:24:@48636.4]
  wire [7:0] x898_x24_1_io_result; // @[Math.scala 150:24:@48636.4]
  wire  x899_x23_1_clock; // @[Math.scala 150:24:@48646.4]
  wire  x899_x23_1_reset; // @[Math.scala 150:24:@48646.4]
  wire [7:0] x899_x23_1_io_a; // @[Math.scala 150:24:@48646.4]
  wire [7:0] x899_x23_1_io_b; // @[Math.scala 150:24:@48646.4]
  wire  x899_x23_1_io_flow; // @[Math.scala 150:24:@48646.4]
  wire [7:0] x899_x23_1_io_result; // @[Math.scala 150:24:@48646.4]
  wire  x900_x24_1_clock; // @[Math.scala 150:24:@48656.4]
  wire  x900_x24_1_reset; // @[Math.scala 150:24:@48656.4]
  wire [7:0] x900_x24_1_io_a; // @[Math.scala 150:24:@48656.4]
  wire [7:0] x900_x24_1_io_b; // @[Math.scala 150:24:@48656.4]
  wire  x900_x24_1_io_flow; // @[Math.scala 150:24:@48656.4]
  wire [7:0] x900_x24_1_io_result; // @[Math.scala 150:24:@48656.4]
  wire [7:0] x901_x23_1_io_a; // @[Math.scala 150:24:@48666.4]
  wire [7:0] x901_x23_1_io_b; // @[Math.scala 150:24:@48666.4]
  wire [7:0] x901_x23_1_io_result; // @[Math.scala 150:24:@48666.4]
  wire [7:0] x902_x24_1_io_a; // @[Math.scala 150:24:@48676.4]
  wire [7:0] x902_x24_1_io_b; // @[Math.scala 150:24:@48676.4]
  wire [7:0] x902_x24_1_io_result; // @[Math.scala 150:24:@48676.4]
  wire [7:0] x903_x23_1_io_a; // @[Math.scala 150:24:@48686.4]
  wire [7:0] x903_x23_1_io_b; // @[Math.scala 150:24:@48686.4]
  wire [7:0] x903_x23_1_io_result; // @[Math.scala 150:24:@48686.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@48696.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@48696.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@48696.4]
  wire [7:0] RetimeWrapper_114_io_in; // @[package.scala 93:22:@48696.4]
  wire [7:0] RetimeWrapper_114_io_out; // @[package.scala 93:22:@48696.4]
  wire [7:0] x904_sum_1_io_a; // @[Math.scala 150:24:@48705.4]
  wire [7:0] x904_sum_1_io_b; // @[Math.scala 150:24:@48705.4]
  wire [7:0] x904_sum_1_io_result; // @[Math.scala 150:24:@48705.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@48719.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@48719.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@48719.4]
  wire [7:0] RetimeWrapper_115_io_in; // @[package.scala 93:22:@48719.4]
  wire [7:0] RetimeWrapper_115_io_out; // @[package.scala 93:22:@48719.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@48729.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@48729.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@48729.4]
  wire  RetimeWrapper_116_io_in; // @[package.scala 93:22:@48729.4]
  wire  RetimeWrapper_116_io_out; // @[package.scala 93:22:@48729.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@48738.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@48738.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@48738.4]
  wire [31:0] RetimeWrapper_117_io_in; // @[package.scala 93:22:@48738.4]
  wire [31:0] RetimeWrapper_117_io_out; // @[package.scala 93:22:@48738.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@48747.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@48747.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@48747.4]
  wire [7:0] RetimeWrapper_118_io_in; // @[package.scala 93:22:@48747.4]
  wire [7:0] RetimeWrapper_118_io_out; // @[package.scala 93:22:@48747.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@48756.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@48756.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@48756.4]
  wire  RetimeWrapper_119_io_in; // @[package.scala 93:22:@48756.4]
  wire  RetimeWrapper_119_io_out; // @[package.scala 93:22:@48756.4]
  wire  RetimeWrapper_120_clock; // @[package.scala 93:22:@48765.4]
  wire  RetimeWrapper_120_reset; // @[package.scala 93:22:@48765.4]
  wire  RetimeWrapper_120_io_flow; // @[package.scala 93:22:@48765.4]
  wire [31:0] RetimeWrapper_120_io_in; // @[package.scala 93:22:@48765.4]
  wire [31:0] RetimeWrapper_120_io_out; // @[package.scala 93:22:@48765.4]
  wire  RetimeWrapper_121_clock; // @[package.scala 93:22:@48778.4]
  wire  RetimeWrapper_121_reset; // @[package.scala 93:22:@48778.4]
  wire  RetimeWrapper_121_io_flow; // @[package.scala 93:22:@48778.4]
  wire  RetimeWrapper_121_io_in; // @[package.scala 93:22:@48778.4]
  wire  RetimeWrapper_121_io_out; // @[package.scala 93:22:@48778.4]
  wire  RetimeWrapper_122_clock; // @[package.scala 93:22:@48799.4]
  wire  RetimeWrapper_122_reset; // @[package.scala 93:22:@48799.4]
  wire  RetimeWrapper_122_io_flow; // @[package.scala 93:22:@48799.4]
  wire [7:0] RetimeWrapper_122_io_in; // @[package.scala 93:22:@48799.4]
  wire [7:0] RetimeWrapper_122_io_out; // @[package.scala 93:22:@48799.4]
  wire  RetimeWrapper_123_clock; // @[package.scala 93:22:@48808.4]
  wire  RetimeWrapper_123_reset; // @[package.scala 93:22:@48808.4]
  wire  RetimeWrapper_123_io_flow; // @[package.scala 93:22:@48808.4]
  wire [31:0] RetimeWrapper_123_io_in; // @[package.scala 93:22:@48808.4]
  wire [31:0] RetimeWrapper_123_io_out; // @[package.scala 93:22:@48808.4]
  wire  RetimeWrapper_124_clock; // @[package.scala 93:22:@48821.4]
  wire  RetimeWrapper_124_reset; // @[package.scala 93:22:@48821.4]
  wire  RetimeWrapper_124_io_flow; // @[package.scala 93:22:@48821.4]
  wire  RetimeWrapper_124_io_in; // @[package.scala 93:22:@48821.4]
  wire  RetimeWrapper_124_io_out; // @[package.scala 93:22:@48821.4]
  wire  RetimeWrapper_125_clock; // @[package.scala 93:22:@48842.4]
  wire  RetimeWrapper_125_reset; // @[package.scala 93:22:@48842.4]
  wire  RetimeWrapper_125_io_flow; // @[package.scala 93:22:@48842.4]
  wire [31:0] RetimeWrapper_125_io_in; // @[package.scala 93:22:@48842.4]
  wire [31:0] RetimeWrapper_125_io_out; // @[package.scala 93:22:@48842.4]
  wire  RetimeWrapper_126_clock; // @[package.scala 93:22:@48851.4]
  wire  RetimeWrapper_126_reset; // @[package.scala 93:22:@48851.4]
  wire  RetimeWrapper_126_io_flow; // @[package.scala 93:22:@48851.4]
  wire [7:0] RetimeWrapper_126_io_in; // @[package.scala 93:22:@48851.4]
  wire [7:0] RetimeWrapper_126_io_out; // @[package.scala 93:22:@48851.4]
  wire  RetimeWrapper_127_clock; // @[package.scala 93:22:@48864.4]
  wire  RetimeWrapper_127_reset; // @[package.scala 93:22:@48864.4]
  wire  RetimeWrapper_127_io_flow; // @[package.scala 93:22:@48864.4]
  wire  RetimeWrapper_127_io_in; // @[package.scala 93:22:@48864.4]
  wire  RetimeWrapper_127_io_out; // @[package.scala 93:22:@48864.4]
  wire  RetimeWrapper_128_clock; // @[package.scala 93:22:@48885.4]
  wire  RetimeWrapper_128_reset; // @[package.scala 93:22:@48885.4]
  wire  RetimeWrapper_128_io_flow; // @[package.scala 93:22:@48885.4]
  wire [31:0] RetimeWrapper_128_io_in; // @[package.scala 93:22:@48885.4]
  wire [31:0] RetimeWrapper_128_io_out; // @[package.scala 93:22:@48885.4]
  wire  RetimeWrapper_129_clock; // @[package.scala 93:22:@48894.4]
  wire  RetimeWrapper_129_reset; // @[package.scala 93:22:@48894.4]
  wire  RetimeWrapper_129_io_flow; // @[package.scala 93:22:@48894.4]
  wire [7:0] RetimeWrapper_129_io_in; // @[package.scala 93:22:@48894.4]
  wire [7:0] RetimeWrapper_129_io_out; // @[package.scala 93:22:@48894.4]
  wire  RetimeWrapper_130_clock; // @[package.scala 93:22:@48907.4]
  wire  RetimeWrapper_130_reset; // @[package.scala 93:22:@48907.4]
  wire  RetimeWrapper_130_io_flow; // @[package.scala 93:22:@48907.4]
  wire  RetimeWrapper_130_io_in; // @[package.scala 93:22:@48907.4]
  wire  RetimeWrapper_130_io_out; // @[package.scala 93:22:@48907.4]
  wire  RetimeWrapper_131_clock; // @[package.scala 93:22:@48928.4]
  wire  RetimeWrapper_131_reset; // @[package.scala 93:22:@48928.4]
  wire  RetimeWrapper_131_io_flow; // @[package.scala 93:22:@48928.4]
  wire [31:0] RetimeWrapper_131_io_in; // @[package.scala 93:22:@48928.4]
  wire [31:0] RetimeWrapper_131_io_out; // @[package.scala 93:22:@48928.4]
  wire  RetimeWrapper_132_clock; // @[package.scala 93:22:@48937.4]
  wire  RetimeWrapper_132_reset; // @[package.scala 93:22:@48937.4]
  wire  RetimeWrapper_132_io_flow; // @[package.scala 93:22:@48937.4]
  wire [7:0] RetimeWrapper_132_io_in; // @[package.scala 93:22:@48937.4]
  wire [7:0] RetimeWrapper_132_io_out; // @[package.scala 93:22:@48937.4]
  wire  RetimeWrapper_133_clock; // @[package.scala 93:22:@48946.4]
  wire  RetimeWrapper_133_reset; // @[package.scala 93:22:@48946.4]
  wire  RetimeWrapper_133_io_flow; // @[package.scala 93:22:@48946.4]
  wire [31:0] RetimeWrapper_133_io_in; // @[package.scala 93:22:@48946.4]
  wire [31:0] RetimeWrapper_133_io_out; // @[package.scala 93:22:@48946.4]
  wire  RetimeWrapper_134_clock; // @[package.scala 93:22:@48959.4]
  wire  RetimeWrapper_134_reset; // @[package.scala 93:22:@48959.4]
  wire  RetimeWrapper_134_io_flow; // @[package.scala 93:22:@48959.4]
  wire  RetimeWrapper_134_io_in; // @[package.scala 93:22:@48959.4]
  wire  RetimeWrapper_134_io_out; // @[package.scala 93:22:@48959.4]
  wire  RetimeWrapper_135_clock; // @[package.scala 93:22:@48980.4]
  wire  RetimeWrapper_135_reset; // @[package.scala 93:22:@48980.4]
  wire  RetimeWrapper_135_io_flow; // @[package.scala 93:22:@48980.4]
  wire [7:0] RetimeWrapper_135_io_in; // @[package.scala 93:22:@48980.4]
  wire [7:0] RetimeWrapper_135_io_out; // @[package.scala 93:22:@48980.4]
  wire  RetimeWrapper_136_clock; // @[package.scala 93:22:@48989.4]
  wire  RetimeWrapper_136_reset; // @[package.scala 93:22:@48989.4]
  wire  RetimeWrapper_136_io_flow; // @[package.scala 93:22:@48989.4]
  wire [31:0] RetimeWrapper_136_io_in; // @[package.scala 93:22:@48989.4]
  wire [31:0] RetimeWrapper_136_io_out; // @[package.scala 93:22:@48989.4]
  wire  RetimeWrapper_137_clock; // @[package.scala 93:22:@49002.4]
  wire  RetimeWrapper_137_reset; // @[package.scala 93:22:@49002.4]
  wire  RetimeWrapper_137_io_flow; // @[package.scala 93:22:@49002.4]
  wire  RetimeWrapper_137_io_in; // @[package.scala 93:22:@49002.4]
  wire  RetimeWrapper_137_io_out; // @[package.scala 93:22:@49002.4]
  wire  RetimeWrapper_138_clock; // @[package.scala 93:22:@49023.4]
  wire  RetimeWrapper_138_reset; // @[package.scala 93:22:@49023.4]
  wire  RetimeWrapper_138_io_flow; // @[package.scala 93:22:@49023.4]
  wire [7:0] RetimeWrapper_138_io_in; // @[package.scala 93:22:@49023.4]
  wire [7:0] RetimeWrapper_138_io_out; // @[package.scala 93:22:@49023.4]
  wire  RetimeWrapper_139_clock; // @[package.scala 93:22:@49032.4]
  wire  RetimeWrapper_139_reset; // @[package.scala 93:22:@49032.4]
  wire  RetimeWrapper_139_io_flow; // @[package.scala 93:22:@49032.4]
  wire [31:0] RetimeWrapper_139_io_in; // @[package.scala 93:22:@49032.4]
  wire [31:0] RetimeWrapper_139_io_out; // @[package.scala 93:22:@49032.4]
  wire  RetimeWrapper_140_clock; // @[package.scala 93:22:@49045.4]
  wire  RetimeWrapper_140_reset; // @[package.scala 93:22:@49045.4]
  wire  RetimeWrapper_140_io_flow; // @[package.scala 93:22:@49045.4]
  wire  RetimeWrapper_140_io_in; // @[package.scala 93:22:@49045.4]
  wire  RetimeWrapper_140_io_out; // @[package.scala 93:22:@49045.4]
  wire  RetimeWrapper_141_clock; // @[package.scala 93:22:@49066.4]
  wire  RetimeWrapper_141_reset; // @[package.scala 93:22:@49066.4]
  wire  RetimeWrapper_141_io_flow; // @[package.scala 93:22:@49066.4]
  wire [31:0] RetimeWrapper_141_io_in; // @[package.scala 93:22:@49066.4]
  wire [31:0] RetimeWrapper_141_io_out; // @[package.scala 93:22:@49066.4]
  wire  RetimeWrapper_142_clock; // @[package.scala 93:22:@49075.4]
  wire  RetimeWrapper_142_reset; // @[package.scala 93:22:@49075.4]
  wire  RetimeWrapper_142_io_flow; // @[package.scala 93:22:@49075.4]
  wire [7:0] RetimeWrapper_142_io_in; // @[package.scala 93:22:@49075.4]
  wire [7:0] RetimeWrapper_142_io_out; // @[package.scala 93:22:@49075.4]
  wire  RetimeWrapper_143_clock; // @[package.scala 93:22:@49088.4]
  wire  RetimeWrapper_143_reset; // @[package.scala 93:22:@49088.4]
  wire  RetimeWrapper_143_io_flow; // @[package.scala 93:22:@49088.4]
  wire  RetimeWrapper_143_io_in; // @[package.scala 93:22:@49088.4]
  wire  RetimeWrapper_143_io_out; // @[package.scala 93:22:@49088.4]
  wire  RetimeWrapper_144_clock; // @[package.scala 93:22:@49109.4]
  wire  RetimeWrapper_144_reset; // @[package.scala 93:22:@49109.4]
  wire  RetimeWrapper_144_io_flow; // @[package.scala 93:22:@49109.4]
  wire  RetimeWrapper_144_io_in; // @[package.scala 93:22:@49109.4]
  wire  RetimeWrapper_144_io_out; // @[package.scala 93:22:@49109.4]
  wire  RetimeWrapper_145_clock; // @[package.scala 93:22:@49118.4]
  wire  RetimeWrapper_145_reset; // @[package.scala 93:22:@49118.4]
  wire  RetimeWrapper_145_io_flow; // @[package.scala 93:22:@49118.4]
  wire  RetimeWrapper_145_io_in; // @[package.scala 93:22:@49118.4]
  wire  RetimeWrapper_145_io_out; // @[package.scala 93:22:@49118.4]
  wire  RetimeWrapper_146_clock; // @[package.scala 93:22:@49127.4]
  wire  RetimeWrapper_146_reset; // @[package.scala 93:22:@49127.4]
  wire  RetimeWrapper_146_io_flow; // @[package.scala 93:22:@49127.4]
  wire  RetimeWrapper_146_io_in; // @[package.scala 93:22:@49127.4]
  wire  RetimeWrapper_146_io_out; // @[package.scala 93:22:@49127.4]
  wire  RetimeWrapper_147_clock; // @[package.scala 93:22:@49136.4]
  wire  RetimeWrapper_147_reset; // @[package.scala 93:22:@49136.4]
  wire  RetimeWrapper_147_io_flow; // @[package.scala 93:22:@49136.4]
  wire [31:0] RetimeWrapper_147_io_in; // @[package.scala 93:22:@49136.4]
  wire [31:0] RetimeWrapper_147_io_out; // @[package.scala 93:22:@49136.4]
  wire  RetimeWrapper_148_clock; // @[package.scala 93:22:@49145.4]
  wire  RetimeWrapper_148_reset; // @[package.scala 93:22:@49145.4]
  wire  RetimeWrapper_148_io_flow; // @[package.scala 93:22:@49145.4]
  wire [31:0] RetimeWrapper_148_io_in; // @[package.scala 93:22:@49145.4]
  wire [31:0] RetimeWrapper_148_io_out; // @[package.scala 93:22:@49145.4]
  wire  RetimeWrapper_149_clock; // @[package.scala 93:22:@49159.4]
  wire  RetimeWrapper_149_reset; // @[package.scala 93:22:@49159.4]
  wire  RetimeWrapper_149_io_flow; // @[package.scala 93:22:@49159.4]
  wire  RetimeWrapper_149_io_in; // @[package.scala 93:22:@49159.4]
  wire  RetimeWrapper_149_io_out; // @[package.scala 93:22:@49159.4]
  wire  RetimeWrapper_150_clock; // @[package.scala 93:22:@49180.4]
  wire  RetimeWrapper_150_reset; // @[package.scala 93:22:@49180.4]
  wire  RetimeWrapper_150_io_flow; // @[package.scala 93:22:@49180.4]
  wire [31:0] RetimeWrapper_150_io_in; // @[package.scala 93:22:@49180.4]
  wire [31:0] RetimeWrapper_150_io_out; // @[package.scala 93:22:@49180.4]
  wire  RetimeWrapper_151_clock; // @[package.scala 93:22:@49189.4]
  wire  RetimeWrapper_151_reset; // @[package.scala 93:22:@49189.4]
  wire  RetimeWrapper_151_io_flow; // @[package.scala 93:22:@49189.4]
  wire  RetimeWrapper_151_io_in; // @[package.scala 93:22:@49189.4]
  wire  RetimeWrapper_151_io_out; // @[package.scala 93:22:@49189.4]
  wire  RetimeWrapper_152_clock; // @[package.scala 93:22:@49203.4]
  wire  RetimeWrapper_152_reset; // @[package.scala 93:22:@49203.4]
  wire  RetimeWrapper_152_io_flow; // @[package.scala 93:22:@49203.4]
  wire  RetimeWrapper_152_io_in; // @[package.scala 93:22:@49203.4]
  wire  RetimeWrapper_152_io_out; // @[package.scala 93:22:@49203.4]
  wire  RetimeWrapper_153_clock; // @[package.scala 93:22:@49224.4]
  wire  RetimeWrapper_153_reset; // @[package.scala 93:22:@49224.4]
  wire  RetimeWrapper_153_io_flow; // @[package.scala 93:22:@49224.4]
  wire  RetimeWrapper_153_io_in; // @[package.scala 93:22:@49224.4]
  wire  RetimeWrapper_153_io_out; // @[package.scala 93:22:@49224.4]
  wire  RetimeWrapper_154_clock; // @[package.scala 93:22:@49233.4]
  wire  RetimeWrapper_154_reset; // @[package.scala 93:22:@49233.4]
  wire  RetimeWrapper_154_io_flow; // @[package.scala 93:22:@49233.4]
  wire [31:0] RetimeWrapper_154_io_in; // @[package.scala 93:22:@49233.4]
  wire [31:0] RetimeWrapper_154_io_out; // @[package.scala 93:22:@49233.4]
  wire  RetimeWrapper_155_clock; // @[package.scala 93:22:@49247.4]
  wire  RetimeWrapper_155_reset; // @[package.scala 93:22:@49247.4]
  wire  RetimeWrapper_155_io_flow; // @[package.scala 93:22:@49247.4]
  wire  RetimeWrapper_155_io_in; // @[package.scala 93:22:@49247.4]
  wire  RetimeWrapper_155_io_out; // @[package.scala 93:22:@49247.4]
  wire  RetimeWrapper_156_clock; // @[package.scala 93:22:@49268.4]
  wire  RetimeWrapper_156_reset; // @[package.scala 93:22:@49268.4]
  wire  RetimeWrapper_156_io_flow; // @[package.scala 93:22:@49268.4]
  wire [31:0] RetimeWrapper_156_io_in; // @[package.scala 93:22:@49268.4]
  wire [31:0] RetimeWrapper_156_io_out; // @[package.scala 93:22:@49268.4]
  wire  RetimeWrapper_157_clock; // @[package.scala 93:22:@49277.4]
  wire  RetimeWrapper_157_reset; // @[package.scala 93:22:@49277.4]
  wire  RetimeWrapper_157_io_flow; // @[package.scala 93:22:@49277.4]
  wire  RetimeWrapper_157_io_in; // @[package.scala 93:22:@49277.4]
  wire  RetimeWrapper_157_io_out; // @[package.scala 93:22:@49277.4]
  wire  RetimeWrapper_158_clock; // @[package.scala 93:22:@49291.4]
  wire  RetimeWrapper_158_reset; // @[package.scala 93:22:@49291.4]
  wire  RetimeWrapper_158_io_flow; // @[package.scala 93:22:@49291.4]
  wire  RetimeWrapper_158_io_in; // @[package.scala 93:22:@49291.4]
  wire  RetimeWrapper_158_io_out; // @[package.scala 93:22:@49291.4]
  wire  RetimeWrapper_159_clock; // @[package.scala 93:22:@49312.4]
  wire  RetimeWrapper_159_reset; // @[package.scala 93:22:@49312.4]
  wire  RetimeWrapper_159_io_flow; // @[package.scala 93:22:@49312.4]
  wire [31:0] RetimeWrapper_159_io_in; // @[package.scala 93:22:@49312.4]
  wire [31:0] RetimeWrapper_159_io_out; // @[package.scala 93:22:@49312.4]
  wire  RetimeWrapper_160_clock; // @[package.scala 93:22:@49321.4]
  wire  RetimeWrapper_160_reset; // @[package.scala 93:22:@49321.4]
  wire  RetimeWrapper_160_io_flow; // @[package.scala 93:22:@49321.4]
  wire  RetimeWrapper_160_io_in; // @[package.scala 93:22:@49321.4]
  wire  RetimeWrapper_160_io_out; // @[package.scala 93:22:@49321.4]
  wire  RetimeWrapper_161_clock; // @[package.scala 93:22:@49335.4]
  wire  RetimeWrapper_161_reset; // @[package.scala 93:22:@49335.4]
  wire  RetimeWrapper_161_io_flow; // @[package.scala 93:22:@49335.4]
  wire  RetimeWrapper_161_io_in; // @[package.scala 93:22:@49335.4]
  wire  RetimeWrapper_161_io_out; // @[package.scala 93:22:@49335.4]
  wire  RetimeWrapper_162_clock; // @[package.scala 93:22:@49356.4]
  wire  RetimeWrapper_162_reset; // @[package.scala 93:22:@49356.4]
  wire  RetimeWrapper_162_io_flow; // @[package.scala 93:22:@49356.4]
  wire  RetimeWrapper_162_io_in; // @[package.scala 93:22:@49356.4]
  wire  RetimeWrapper_162_io_out; // @[package.scala 93:22:@49356.4]
  wire  RetimeWrapper_163_clock; // @[package.scala 93:22:@49365.4]
  wire  RetimeWrapper_163_reset; // @[package.scala 93:22:@49365.4]
  wire  RetimeWrapper_163_io_flow; // @[package.scala 93:22:@49365.4]
  wire [31:0] RetimeWrapper_163_io_in; // @[package.scala 93:22:@49365.4]
  wire [31:0] RetimeWrapper_163_io_out; // @[package.scala 93:22:@49365.4]
  wire  RetimeWrapper_164_clock; // @[package.scala 93:22:@49374.4]
  wire  RetimeWrapper_164_reset; // @[package.scala 93:22:@49374.4]
  wire  RetimeWrapper_164_io_flow; // @[package.scala 93:22:@49374.4]
  wire [31:0] RetimeWrapper_164_io_in; // @[package.scala 93:22:@49374.4]
  wire [31:0] RetimeWrapper_164_io_out; // @[package.scala 93:22:@49374.4]
  wire  RetimeWrapper_165_clock; // @[package.scala 93:22:@49388.4]
  wire  RetimeWrapper_165_reset; // @[package.scala 93:22:@49388.4]
  wire  RetimeWrapper_165_io_flow; // @[package.scala 93:22:@49388.4]
  wire  RetimeWrapper_165_io_in; // @[package.scala 93:22:@49388.4]
  wire  RetimeWrapper_165_io_out; // @[package.scala 93:22:@49388.4]
  wire  RetimeWrapper_166_clock; // @[package.scala 93:22:@49409.4]
  wire  RetimeWrapper_166_reset; // @[package.scala 93:22:@49409.4]
  wire  RetimeWrapper_166_io_flow; // @[package.scala 93:22:@49409.4]
  wire [31:0] RetimeWrapper_166_io_in; // @[package.scala 93:22:@49409.4]
  wire [31:0] RetimeWrapper_166_io_out; // @[package.scala 93:22:@49409.4]
  wire  RetimeWrapper_167_clock; // @[package.scala 93:22:@49418.4]
  wire  RetimeWrapper_167_reset; // @[package.scala 93:22:@49418.4]
  wire  RetimeWrapper_167_io_flow; // @[package.scala 93:22:@49418.4]
  wire  RetimeWrapper_167_io_in; // @[package.scala 93:22:@49418.4]
  wire  RetimeWrapper_167_io_out; // @[package.scala 93:22:@49418.4]
  wire  RetimeWrapper_168_clock; // @[package.scala 93:22:@49432.4]
  wire  RetimeWrapper_168_reset; // @[package.scala 93:22:@49432.4]
  wire  RetimeWrapper_168_io_flow; // @[package.scala 93:22:@49432.4]
  wire  RetimeWrapper_168_io_in; // @[package.scala 93:22:@49432.4]
  wire  RetimeWrapper_168_io_out; // @[package.scala 93:22:@49432.4]
  wire  RetimeWrapper_169_clock; // @[package.scala 93:22:@49453.4]
  wire  RetimeWrapper_169_reset; // @[package.scala 93:22:@49453.4]
  wire  RetimeWrapper_169_io_flow; // @[package.scala 93:22:@49453.4]
  wire  RetimeWrapper_169_io_in; // @[package.scala 93:22:@49453.4]
  wire  RetimeWrapper_169_io_out; // @[package.scala 93:22:@49453.4]
  wire  RetimeWrapper_170_clock; // @[package.scala 93:22:@49462.4]
  wire  RetimeWrapper_170_reset; // @[package.scala 93:22:@49462.4]
  wire  RetimeWrapper_170_io_flow; // @[package.scala 93:22:@49462.4]
  wire [31:0] RetimeWrapper_170_io_in; // @[package.scala 93:22:@49462.4]
  wire [31:0] RetimeWrapper_170_io_out; // @[package.scala 93:22:@49462.4]
  wire  RetimeWrapper_171_clock; // @[package.scala 93:22:@49476.4]
  wire  RetimeWrapper_171_reset; // @[package.scala 93:22:@49476.4]
  wire  RetimeWrapper_171_io_flow; // @[package.scala 93:22:@49476.4]
  wire  RetimeWrapper_171_io_in; // @[package.scala 93:22:@49476.4]
  wire  RetimeWrapper_171_io_out; // @[package.scala 93:22:@49476.4]
  wire  RetimeWrapper_172_clock; // @[package.scala 93:22:@49497.4]
  wire  RetimeWrapper_172_reset; // @[package.scala 93:22:@49497.4]
  wire  RetimeWrapper_172_io_flow; // @[package.scala 93:22:@49497.4]
  wire  RetimeWrapper_172_io_in; // @[package.scala 93:22:@49497.4]
  wire  RetimeWrapper_172_io_out; // @[package.scala 93:22:@49497.4]
  wire  RetimeWrapper_173_clock; // @[package.scala 93:22:@49506.4]
  wire  RetimeWrapper_173_reset; // @[package.scala 93:22:@49506.4]
  wire  RetimeWrapper_173_io_flow; // @[package.scala 93:22:@49506.4]
  wire [31:0] RetimeWrapper_173_io_in; // @[package.scala 93:22:@49506.4]
  wire [31:0] RetimeWrapper_173_io_out; // @[package.scala 93:22:@49506.4]
  wire  RetimeWrapper_174_clock; // @[package.scala 93:22:@49520.4]
  wire  RetimeWrapper_174_reset; // @[package.scala 93:22:@49520.4]
  wire  RetimeWrapper_174_io_flow; // @[package.scala 93:22:@49520.4]
  wire  RetimeWrapper_174_io_in; // @[package.scala 93:22:@49520.4]
  wire  RetimeWrapper_174_io_out; // @[package.scala 93:22:@49520.4]
  wire  RetimeWrapper_175_clock; // @[package.scala 93:22:@49541.4]
  wire  RetimeWrapper_175_reset; // @[package.scala 93:22:@49541.4]
  wire  RetimeWrapper_175_io_flow; // @[package.scala 93:22:@49541.4]
  wire [31:0] RetimeWrapper_175_io_in; // @[package.scala 93:22:@49541.4]
  wire [31:0] RetimeWrapper_175_io_out; // @[package.scala 93:22:@49541.4]
  wire  RetimeWrapper_176_clock; // @[package.scala 93:22:@49550.4]
  wire  RetimeWrapper_176_reset; // @[package.scala 93:22:@49550.4]
  wire  RetimeWrapper_176_io_flow; // @[package.scala 93:22:@49550.4]
  wire  RetimeWrapper_176_io_in; // @[package.scala 93:22:@49550.4]
  wire  RetimeWrapper_176_io_out; // @[package.scala 93:22:@49550.4]
  wire  RetimeWrapper_177_clock; // @[package.scala 93:22:@49564.4]
  wire  RetimeWrapper_177_reset; // @[package.scala 93:22:@49564.4]
  wire  RetimeWrapper_177_io_flow; // @[package.scala 93:22:@49564.4]
  wire  RetimeWrapper_177_io_in; // @[package.scala 93:22:@49564.4]
  wire  RetimeWrapper_177_io_out; // @[package.scala 93:22:@49564.4]
  wire  RetimeWrapper_178_clock; // @[package.scala 93:22:@49585.4]
  wire  RetimeWrapper_178_reset; // @[package.scala 93:22:@49585.4]
  wire  RetimeWrapper_178_io_flow; // @[package.scala 93:22:@49585.4]
  wire  RetimeWrapper_178_io_in; // @[package.scala 93:22:@49585.4]
  wire  RetimeWrapper_178_io_out; // @[package.scala 93:22:@49585.4]
  wire  RetimeWrapper_179_clock; // @[package.scala 93:22:@49594.4]
  wire  RetimeWrapper_179_reset; // @[package.scala 93:22:@49594.4]
  wire  RetimeWrapper_179_io_flow; // @[package.scala 93:22:@49594.4]
  wire [31:0] RetimeWrapper_179_io_in; // @[package.scala 93:22:@49594.4]
  wire [31:0] RetimeWrapper_179_io_out; // @[package.scala 93:22:@49594.4]
  wire  RetimeWrapper_180_clock; // @[package.scala 93:22:@49603.4]
  wire  RetimeWrapper_180_reset; // @[package.scala 93:22:@49603.4]
  wire  RetimeWrapper_180_io_flow; // @[package.scala 93:22:@49603.4]
  wire [31:0] RetimeWrapper_180_io_in; // @[package.scala 93:22:@49603.4]
  wire [31:0] RetimeWrapper_180_io_out; // @[package.scala 93:22:@49603.4]
  wire  RetimeWrapper_181_clock; // @[package.scala 93:22:@49617.4]
  wire  RetimeWrapper_181_reset; // @[package.scala 93:22:@49617.4]
  wire  RetimeWrapper_181_io_flow; // @[package.scala 93:22:@49617.4]
  wire  RetimeWrapper_181_io_in; // @[package.scala 93:22:@49617.4]
  wire  RetimeWrapper_181_io_out; // @[package.scala 93:22:@49617.4]
  wire  RetimeWrapper_182_clock; // @[package.scala 93:22:@49638.4]
  wire  RetimeWrapper_182_reset; // @[package.scala 93:22:@49638.4]
  wire  RetimeWrapper_182_io_flow; // @[package.scala 93:22:@49638.4]
  wire  RetimeWrapper_182_io_in; // @[package.scala 93:22:@49638.4]
  wire  RetimeWrapper_182_io_out; // @[package.scala 93:22:@49638.4]
  wire  RetimeWrapper_183_clock; // @[package.scala 93:22:@49647.4]
  wire  RetimeWrapper_183_reset; // @[package.scala 93:22:@49647.4]
  wire  RetimeWrapper_183_io_flow; // @[package.scala 93:22:@49647.4]
  wire [31:0] RetimeWrapper_183_io_in; // @[package.scala 93:22:@49647.4]
  wire [31:0] RetimeWrapper_183_io_out; // @[package.scala 93:22:@49647.4]
  wire  RetimeWrapper_184_clock; // @[package.scala 93:22:@49661.4]
  wire  RetimeWrapper_184_reset; // @[package.scala 93:22:@49661.4]
  wire  RetimeWrapper_184_io_flow; // @[package.scala 93:22:@49661.4]
  wire  RetimeWrapper_184_io_in; // @[package.scala 93:22:@49661.4]
  wire  RetimeWrapper_184_io_out; // @[package.scala 93:22:@49661.4]
  wire  RetimeWrapper_185_clock; // @[package.scala 93:22:@49682.4]
  wire  RetimeWrapper_185_reset; // @[package.scala 93:22:@49682.4]
  wire  RetimeWrapper_185_io_flow; // @[package.scala 93:22:@49682.4]
  wire [31:0] RetimeWrapper_185_io_in; // @[package.scala 93:22:@49682.4]
  wire [31:0] RetimeWrapper_185_io_out; // @[package.scala 93:22:@49682.4]
  wire  RetimeWrapper_186_clock; // @[package.scala 93:22:@49691.4]
  wire  RetimeWrapper_186_reset; // @[package.scala 93:22:@49691.4]
  wire  RetimeWrapper_186_io_flow; // @[package.scala 93:22:@49691.4]
  wire  RetimeWrapper_186_io_in; // @[package.scala 93:22:@49691.4]
  wire  RetimeWrapper_186_io_out; // @[package.scala 93:22:@49691.4]
  wire  RetimeWrapper_187_clock; // @[package.scala 93:22:@49705.4]
  wire  RetimeWrapper_187_reset; // @[package.scala 93:22:@49705.4]
  wire  RetimeWrapper_187_io_flow; // @[package.scala 93:22:@49705.4]
  wire  RetimeWrapper_187_io_in; // @[package.scala 93:22:@49705.4]
  wire  RetimeWrapper_187_io_out; // @[package.scala 93:22:@49705.4]
  wire  RetimeWrapper_188_clock; // @[package.scala 93:22:@49726.4]
  wire  RetimeWrapper_188_reset; // @[package.scala 93:22:@49726.4]
  wire  RetimeWrapper_188_io_flow; // @[package.scala 93:22:@49726.4]
  wire  RetimeWrapper_188_io_in; // @[package.scala 93:22:@49726.4]
  wire  RetimeWrapper_188_io_out; // @[package.scala 93:22:@49726.4]
  wire  RetimeWrapper_189_clock; // @[package.scala 93:22:@49735.4]
  wire  RetimeWrapper_189_reset; // @[package.scala 93:22:@49735.4]
  wire  RetimeWrapper_189_io_flow; // @[package.scala 93:22:@49735.4]
  wire [31:0] RetimeWrapper_189_io_in; // @[package.scala 93:22:@49735.4]
  wire [31:0] RetimeWrapper_189_io_out; // @[package.scala 93:22:@49735.4]
  wire  RetimeWrapper_190_clock; // @[package.scala 93:22:@49749.4]
  wire  RetimeWrapper_190_reset; // @[package.scala 93:22:@49749.4]
  wire  RetimeWrapper_190_io_flow; // @[package.scala 93:22:@49749.4]
  wire  RetimeWrapper_190_io_in; // @[package.scala 93:22:@49749.4]
  wire  RetimeWrapper_190_io_out; // @[package.scala 93:22:@49749.4]
  wire  RetimeWrapper_191_clock; // @[package.scala 93:22:@49770.4]
  wire  RetimeWrapper_191_reset; // @[package.scala 93:22:@49770.4]
  wire  RetimeWrapper_191_io_flow; // @[package.scala 93:22:@49770.4]
  wire [31:0] RetimeWrapper_191_io_in; // @[package.scala 93:22:@49770.4]
  wire [31:0] RetimeWrapper_191_io_out; // @[package.scala 93:22:@49770.4]
  wire  RetimeWrapper_192_clock; // @[package.scala 93:22:@49779.4]
  wire  RetimeWrapper_192_reset; // @[package.scala 93:22:@49779.4]
  wire  RetimeWrapper_192_io_flow; // @[package.scala 93:22:@49779.4]
  wire  RetimeWrapper_192_io_in; // @[package.scala 93:22:@49779.4]
  wire  RetimeWrapper_192_io_out; // @[package.scala 93:22:@49779.4]
  wire  RetimeWrapper_193_clock; // @[package.scala 93:22:@49793.4]
  wire  RetimeWrapper_193_reset; // @[package.scala 93:22:@49793.4]
  wire  RetimeWrapper_193_io_flow; // @[package.scala 93:22:@49793.4]
  wire  RetimeWrapper_193_io_in; // @[package.scala 93:22:@49793.4]
  wire  RetimeWrapper_193_io_out; // @[package.scala 93:22:@49793.4]
  wire [7:0] x948_x25_1_io_a; // @[Math.scala 150:24:@49826.4]
  wire [7:0] x948_x25_1_io_b; // @[Math.scala 150:24:@49826.4]
  wire [7:0] x948_x25_1_io_result; // @[Math.scala 150:24:@49826.4]
  wire [7:0] x949_x26_1_io_a; // @[Math.scala 150:24:@49836.4]
  wire [7:0] x949_x26_1_io_b; // @[Math.scala 150:24:@49836.4]
  wire [7:0] x949_x26_1_io_result; // @[Math.scala 150:24:@49836.4]
  wire [7:0] x950_sum_1_io_a; // @[Math.scala 150:24:@49846.4]
  wire [7:0] x950_sum_1_io_b; // @[Math.scala 150:24:@49846.4]
  wire [7:0] x950_sum_1_io_result; // @[Math.scala 150:24:@49846.4]
  wire  x951_div_1_clock; // @[Math.scala 327:24:@49858.4]
  wire  x951_div_1_reset; // @[Math.scala 327:24:@49858.4]
  wire [7:0] x951_div_1_io_a; // @[Math.scala 327:24:@49858.4]
  wire  x951_div_1_io_flow; // @[Math.scala 327:24:@49858.4]
  wire [7:0] x951_div_1_io_result; // @[Math.scala 327:24:@49858.4]
  wire [7:0] x954_x25_1_io_a; // @[Math.scala 150:24:@49878.4]
  wire [7:0] x954_x25_1_io_b; // @[Math.scala 150:24:@49878.4]
  wire [7:0] x954_x25_1_io_result; // @[Math.scala 150:24:@49878.4]
  wire [7:0] x955_x26_1_io_a; // @[Math.scala 150:24:@49888.4]
  wire [7:0] x955_x26_1_io_b; // @[Math.scala 150:24:@49888.4]
  wire [7:0] x955_x26_1_io_result; // @[Math.scala 150:24:@49888.4]
  wire [7:0] x956_sum_1_io_a; // @[Math.scala 150:24:@49898.4]
  wire [7:0] x956_sum_1_io_b; // @[Math.scala 150:24:@49898.4]
  wire [7:0] x956_sum_1_io_result; // @[Math.scala 150:24:@49898.4]
  wire  x957_div_1_clock; // @[Math.scala 327:24:@49910.4]
  wire  x957_div_1_reset; // @[Math.scala 327:24:@49910.4]
  wire [7:0] x957_div_1_io_a; // @[Math.scala 327:24:@49910.4]
  wire  x957_div_1_io_flow; // @[Math.scala 327:24:@49910.4]
  wire [7:0] x957_div_1_io_result; // @[Math.scala 327:24:@49910.4]
  wire [7:0] x960_x25_1_io_a; // @[Math.scala 150:24:@49930.4]
  wire [7:0] x960_x25_1_io_b; // @[Math.scala 150:24:@49930.4]
  wire [7:0] x960_x25_1_io_result; // @[Math.scala 150:24:@49930.4]
  wire [7:0] x961_x26_1_io_a; // @[Math.scala 150:24:@49940.4]
  wire [7:0] x961_x26_1_io_b; // @[Math.scala 150:24:@49940.4]
  wire [7:0] x961_x26_1_io_result; // @[Math.scala 150:24:@49940.4]
  wire [7:0] x962_sum_1_io_a; // @[Math.scala 150:24:@49950.4]
  wire [7:0] x962_sum_1_io_b; // @[Math.scala 150:24:@49950.4]
  wire [7:0] x962_sum_1_io_result; // @[Math.scala 150:24:@49950.4]
  wire  x963_div_1_clock; // @[Math.scala 327:24:@49962.4]
  wire  x963_div_1_reset; // @[Math.scala 327:24:@49962.4]
  wire [7:0] x963_div_1_io_a; // @[Math.scala 327:24:@49962.4]
  wire  x963_div_1_io_flow; // @[Math.scala 327:24:@49962.4]
  wire [7:0] x963_div_1_io_result; // @[Math.scala 327:24:@49962.4]
  wire [7:0] x966_x25_1_io_a; // @[Math.scala 150:24:@49984.4]
  wire [7:0] x966_x25_1_io_b; // @[Math.scala 150:24:@49984.4]
  wire [7:0] x966_x25_1_io_result; // @[Math.scala 150:24:@49984.4]
  wire [7:0] x967_x26_1_io_a; // @[Math.scala 150:24:@49994.4]
  wire [7:0] x967_x26_1_io_b; // @[Math.scala 150:24:@49994.4]
  wire [7:0] x967_x26_1_io_result; // @[Math.scala 150:24:@49994.4]
  wire [7:0] x968_sum_1_io_a; // @[Math.scala 150:24:@50004.4]
  wire [7:0] x968_sum_1_io_b; // @[Math.scala 150:24:@50004.4]
  wire [7:0] x968_sum_1_io_result; // @[Math.scala 150:24:@50004.4]
  wire  x969_div_1_clock; // @[Math.scala 327:24:@50016.4]
  wire  x969_div_1_reset; // @[Math.scala 327:24:@50016.4]
  wire [7:0] x969_div_1_io_a; // @[Math.scala 327:24:@50016.4]
  wire  x969_div_1_io_flow; // @[Math.scala 327:24:@50016.4]
  wire [7:0] x969_div_1_io_result; // @[Math.scala 327:24:@50016.4]
  wire [7:0] x971_x25_1_io_a; // @[Math.scala 150:24:@50031.4]
  wire [7:0] x971_x25_1_io_b; // @[Math.scala 150:24:@50031.4]
  wire [7:0] x971_x25_1_io_result; // @[Math.scala 150:24:@50031.4]
  wire [7:0] x972_x26_1_io_a; // @[Math.scala 150:24:@50041.4]
  wire [7:0] x972_x26_1_io_b; // @[Math.scala 150:24:@50041.4]
  wire [7:0] x972_x26_1_io_result; // @[Math.scala 150:24:@50041.4]
  wire [7:0] x973_sum_1_io_a; // @[Math.scala 150:24:@50051.4]
  wire [7:0] x973_sum_1_io_b; // @[Math.scala 150:24:@50051.4]
  wire [7:0] x973_sum_1_io_result; // @[Math.scala 150:24:@50051.4]
  wire  x974_div_1_clock; // @[Math.scala 327:24:@50063.4]
  wire  x974_div_1_reset; // @[Math.scala 327:24:@50063.4]
  wire [7:0] x974_div_1_io_a; // @[Math.scala 327:24:@50063.4]
  wire  x974_div_1_io_flow; // @[Math.scala 327:24:@50063.4]
  wire [7:0] x974_div_1_io_result; // @[Math.scala 327:24:@50063.4]
  wire [7:0] x976_x25_1_io_a; // @[Math.scala 150:24:@50078.4]
  wire [7:0] x976_x25_1_io_b; // @[Math.scala 150:24:@50078.4]
  wire [7:0] x976_x25_1_io_result; // @[Math.scala 150:24:@50078.4]
  wire [7:0] x977_x26_1_io_a; // @[Math.scala 150:24:@50088.4]
  wire [7:0] x977_x26_1_io_b; // @[Math.scala 150:24:@50088.4]
  wire [7:0] x977_x26_1_io_result; // @[Math.scala 150:24:@50088.4]
  wire [7:0] x978_sum_1_io_a; // @[Math.scala 150:24:@50098.4]
  wire [7:0] x978_sum_1_io_b; // @[Math.scala 150:24:@50098.4]
  wire [7:0] x978_sum_1_io_result; // @[Math.scala 150:24:@50098.4]
  wire  x979_div_1_clock; // @[Math.scala 327:24:@50110.4]
  wire  x979_div_1_reset; // @[Math.scala 327:24:@50110.4]
  wire [7:0] x979_div_1_io_a; // @[Math.scala 327:24:@50110.4]
  wire  x979_div_1_io_flow; // @[Math.scala 327:24:@50110.4]
  wire [7:0] x979_div_1_io_result; // @[Math.scala 327:24:@50110.4]
  wire [7:0] x981_x25_1_io_a; // @[Math.scala 150:24:@50125.4]
  wire [7:0] x981_x25_1_io_b; // @[Math.scala 150:24:@50125.4]
  wire [7:0] x981_x25_1_io_result; // @[Math.scala 150:24:@50125.4]
  wire [7:0] x982_x26_1_io_a; // @[Math.scala 150:24:@50135.4]
  wire [7:0] x982_x26_1_io_b; // @[Math.scala 150:24:@50135.4]
  wire [7:0] x982_x26_1_io_result; // @[Math.scala 150:24:@50135.4]
  wire [7:0] x983_sum_1_io_a; // @[Math.scala 150:24:@50145.4]
  wire [7:0] x983_sum_1_io_b; // @[Math.scala 150:24:@50145.4]
  wire [7:0] x983_sum_1_io_result; // @[Math.scala 150:24:@50145.4]
  wire  x984_div_1_clock; // @[Math.scala 327:24:@50157.4]
  wire  x984_div_1_reset; // @[Math.scala 327:24:@50157.4]
  wire [7:0] x984_div_1_io_a; // @[Math.scala 327:24:@50157.4]
  wire  x984_div_1_io_flow; // @[Math.scala 327:24:@50157.4]
  wire [7:0] x984_div_1_io_result; // @[Math.scala 327:24:@50157.4]
  wire [7:0] x987_x25_1_io_a; // @[Math.scala 150:24:@50177.4]
  wire [7:0] x987_x25_1_io_b; // @[Math.scala 150:24:@50177.4]
  wire [7:0] x987_x25_1_io_result; // @[Math.scala 150:24:@50177.4]
  wire [7:0] x988_x26_1_io_a; // @[Math.scala 150:24:@50187.4]
  wire [7:0] x988_x26_1_io_b; // @[Math.scala 150:24:@50187.4]
  wire [7:0] x988_x26_1_io_result; // @[Math.scala 150:24:@50187.4]
  wire [7:0] x989_sum_1_io_a; // @[Math.scala 150:24:@50197.4]
  wire [7:0] x989_sum_1_io_b; // @[Math.scala 150:24:@50197.4]
  wire [7:0] x989_sum_1_io_result; // @[Math.scala 150:24:@50197.4]
  wire  x990_div_1_clock; // @[Math.scala 327:24:@50209.4]
  wire  x990_div_1_reset; // @[Math.scala 327:24:@50209.4]
  wire [7:0] x990_div_1_io_a; // @[Math.scala 327:24:@50209.4]
  wire  x990_div_1_io_flow; // @[Math.scala 327:24:@50209.4]
  wire [7:0] x990_div_1_io_result; // @[Math.scala 327:24:@50209.4]
  wire  RetimeWrapper_194_clock; // @[package.scala 93:22:@50237.4]
  wire  RetimeWrapper_194_reset; // @[package.scala 93:22:@50237.4]
  wire  RetimeWrapper_194_io_flow; // @[package.scala 93:22:@50237.4]
  wire [63:0] RetimeWrapper_194_io_in; // @[package.scala 93:22:@50237.4]
  wire [63:0] RetimeWrapper_194_io_out; // @[package.scala 93:22:@50237.4]
  wire  RetimeWrapper_195_clock; // @[package.scala 93:22:@50246.4]
  wire  RetimeWrapper_195_reset; // @[package.scala 93:22:@50246.4]
  wire  RetimeWrapper_195_io_flow; // @[package.scala 93:22:@50246.4]
  wire  RetimeWrapper_195_io_in; // @[package.scala 93:22:@50246.4]
  wire  RetimeWrapper_195_io_out; // @[package.scala 93:22:@50246.4]
  wire  RetimeWrapper_196_clock; // @[package.scala 93:22:@50255.4]
  wire  RetimeWrapper_196_reset; // @[package.scala 93:22:@50255.4]
  wire  RetimeWrapper_196_io_flow; // @[package.scala 93:22:@50255.4]
  wire  RetimeWrapper_196_io_in; // @[package.scala 93:22:@50255.4]
  wire  RetimeWrapper_196_io_out; // @[package.scala 93:22:@50255.4]
  wire  RetimeWrapper_197_clock; // @[package.scala 93:22:@50264.4]
  wire  RetimeWrapper_197_reset; // @[package.scala 93:22:@50264.4]
  wire  RetimeWrapper_197_io_flow; // @[package.scala 93:22:@50264.4]
  wire  RetimeWrapper_197_io_in; // @[package.scala 93:22:@50264.4]
  wire  RetimeWrapper_197_io_out; // @[package.scala 93:22:@50264.4]
  wire  b522; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 62:18:@44949.4]
  wire  b523; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 63:18:@44950.4]
  wire  _T_207; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 69:30:@45324.4]
  wire  _T_208; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 69:37:@45325.4]
  wire  _T_212; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 71:76:@45330.4]
  wire  _T_213; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 71:62:@45331.4]
  wire  _T_215; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 71:101:@45332.4]
  wire [63:0] x1061_x526_D1_0_number; // @[package.scala 96:25:@45341.4 package.scala 96:25:@45342.4]
  wire [31:0] b520_number; // @[Math.scala 712:22:@44934.4 Math.scala 713:14:@44935.4]
  wire [31:0] _T_255; // @[Math.scala 499:52:@45369.4]
  wire  x530; // @[Math.scala 499:44:@45377.4]
  wire  x531; // @[Math.scala 499:44:@45384.4]
  wire  x532; // @[Math.scala 499:44:@45391.4]
  wire [31:0] _T_302; // @[Mux.scala 19:72:@45403.4]
  wire [31:0] _T_304; // @[Mux.scala 19:72:@45404.4]
  wire [31:0] _T_306; // @[Mux.scala 19:72:@45405.4]
  wire [31:0] _T_308; // @[Mux.scala 19:72:@45407.4]
  wire [31:0] x533_number; // @[Mux.scala 19:72:@45408.4]
  wire [31:0] _T_320; // @[Math.scala 406:49:@45418.4]
  wire [31:0] _T_322; // @[Math.scala 406:56:@45420.4]
  wire [31:0] _T_323; // @[Math.scala 406:56:@45421.4]
  wire  _T_328; // @[FixedPoint.scala 50:25:@45427.4]
  wire [1:0] _T_332; // @[Bitwise.scala 72:12:@45429.4]
  wire [29:0] _T_333; // @[FixedPoint.scala 18:52:@45430.4]
  wire [31:0] b521_number; // @[Math.scala 712:22:@44946.4 Math.scala 713:14:@44947.4]
  wire  _T_338; // @[FixedPoint.scala 50:25:@45436.4]
  wire [1:0] _T_342; // @[Bitwise.scala 72:12:@45438.4]
  wire [29:0] _T_343; // @[FixedPoint.scala 18:52:@45439.4]
  wire  _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 114:101:@45500.4]
  wire  _T_372; // @[package.scala 96:25:@45508.4 package.scala 96:25:@45509.4]
  wire  _T_374; // @[implicits.scala 55:10:@45510.4]
  wire  _T_375; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 114:118:@45511.4]
  wire  _T_377; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 114:205:@45513.4]
  wire  _T_378; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 114:224:@45514.4]
  wire  x1065_b522_D8; // @[package.scala 96:25:@45486.4 package.scala 96:25:@45487.4]
  wire  _T_379; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 114:250:@45515.4]
  wire  x1062_b523_D8; // @[package.scala 96:25:@45459.4 package.scala 96:25:@45460.4]
  wire [31:0] x545_rdcol_number; // @[Math.scala 154:22:@45532.4 Math.scala 155:14:@45533.4]
  wire  _T_392; // @[FixedPoint.scala 50:25:@45539.4]
  wire [1:0] _T_396; // @[Bitwise.scala 72:12:@45541.4]
  wire [29:0] _T_397; // @[FixedPoint.scala 18:52:@45542.4]
  wire  _T_420; // @[package.scala 96:25:@45593.4 package.scala 96:25:@45594.4]
  wire  _T_422; // @[implicits.scala 55:10:@45595.4]
  wire  _T_423; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 133:118:@45596.4]
  wire  _T_425; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 133:205:@45598.4]
  wire  _T_426; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 133:224:@45599.4]
  wire  _T_427; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 133:250:@45600.4]
  wire [31:0] x554_rdcol_number; // @[Math.scala 154:22:@45617.4 Math.scala 155:14:@45618.4]
  wire  _T_440; // @[FixedPoint.scala 50:25:@45624.4]
  wire [1:0] _T_444; // @[Bitwise.scala 72:12:@45626.4]
  wire [29:0] _T_445; // @[FixedPoint.scala 18:52:@45627.4]
  wire  _T_465; // @[package.scala 96:25:@45669.4 package.scala 96:25:@45670.4]
  wire  _T_467; // @[implicits.scala 55:10:@45671.4]
  wire  _T_468; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 150:118:@45672.4]
  wire  _T_470; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 150:205:@45674.4]
  wire  _T_471; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 150:224:@45675.4]
  wire  _T_472; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 150:250:@45676.4]
  wire [31:0] x563_rdcol_number; // @[Math.scala 154:22:@45693.4 Math.scala 155:14:@45694.4]
  wire  _T_485; // @[FixedPoint.scala 50:25:@45700.4]
  wire [1:0] _T_489; // @[Bitwise.scala 72:12:@45702.4]
  wire [29:0] _T_490; // @[FixedPoint.scala 18:52:@45703.4]
  wire  _T_510; // @[package.scala 96:25:@45745.4 package.scala 96:25:@45746.4]
  wire  _T_512; // @[implicits.scala 55:10:@45747.4]
  wire  _T_513; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 167:118:@45748.4]
  wire  _T_515; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 167:205:@45750.4]
  wire  _T_516; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 167:224:@45751.4]
  wire  _T_517; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 167:250:@45752.4]
  wire [31:0] x572_rdrow_number; // @[Math.scala 154:22:@45769.4 Math.scala 155:14:@45770.4]
  wire [31:0] _T_532; // @[Math.scala 499:52:@45776.4]
  wire  x574; // @[Math.scala 499:44:@45784.4]
  wire  x575; // @[Math.scala 499:44:@45791.4]
  wire  x576; // @[Math.scala 499:44:@45798.4]
  wire [31:0] _T_579; // @[Mux.scala 19:72:@45810.4]
  wire [31:0] _T_581; // @[Mux.scala 19:72:@45811.4]
  wire [31:0] _T_583; // @[Mux.scala 19:72:@45812.4]
  wire [31:0] _T_585; // @[Mux.scala 19:72:@45814.4]
  wire [31:0] x577_number; // @[Mux.scala 19:72:@45815.4]
  wire [31:0] _T_599; // @[Math.scala 406:49:@45827.4]
  wire [31:0] _T_601; // @[Math.scala 406:56:@45829.4]
  wire [31:0] _T_602; // @[Math.scala 406:56:@45830.4]
  wire  _T_607; // @[FixedPoint.scala 50:25:@45836.4]
  wire [1:0] _T_611; // @[Bitwise.scala 72:12:@45838.4]
  wire [29:0] _T_612; // @[FixedPoint.scala 18:52:@45839.4]
  wire  _T_638; // @[package.scala 96:25:@45899.4 package.scala 96:25:@45900.4]
  wire  _T_640; // @[implicits.scala 55:10:@45901.4]
  wire  _T_641; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 208:166:@45902.4]
  wire  _T_643; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 208:253:@45904.4]
  wire  _T_644; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 208:272:@45905.4]
  wire  _T_645; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 208:298:@45906.4]
  wire  _T_666; // @[package.scala 96:25:@45954.4 package.scala 96:25:@45955.4]
  wire  _T_668; // @[implicits.scala 55:10:@45956.4]
  wire  _T_669; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 221:166:@45957.4]
  wire  _T_671; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 221:253:@45959.4]
  wire  _T_672; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 221:272:@45960.4]
  wire  _T_673; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 221:298:@45961.4]
  wire  _T_694; // @[package.scala 96:25:@46009.4 package.scala 96:25:@46010.4]
  wire  _T_696; // @[implicits.scala 55:10:@46011.4]
  wire  _T_697; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 234:166:@46012.4]
  wire  _T_699; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 234:253:@46014.4]
  wire  _T_700; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 234:272:@46015.4]
  wire  _T_701; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 234:298:@46016.4]
  wire  _T_722; // @[package.scala 96:25:@46064.4 package.scala 96:25:@46065.4]
  wire  _T_724; // @[implicits.scala 55:10:@46066.4]
  wire  _T_725; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 247:166:@46067.4]
  wire  _T_727; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 247:253:@46069.4]
  wire  _T_728; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 247:272:@46070.4]
  wire  _T_729; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 247:298:@46071.4]
  wire [31:0] x1084_x572_rdrow_D11_number; // @[package.scala 96:25:@46085.4 package.scala 96:25:@46086.4]
  wire [31:0] _T_741; // @[Math.scala 406:49:@46092.4]
  wire [31:0] _T_743; // @[Math.scala 406:56:@46094.4]
  wire [31:0] _T_744; // @[Math.scala 406:56:@46095.4]
  wire [31:0] x1053_number; // @[implicits.scala 133:21:@46096.4]
  wire  x603; // @[Math.scala 465:44:@46104.4]
  wire [31:0] x1085_x563_rdcol_D11_number; // @[package.scala 96:25:@46112.4 package.scala 96:25:@46113.4]
  wire [31:0] _T_762; // @[Math.scala 465:37:@46118.4]
  wire  x604; // @[Math.scala 465:44:@46120.4]
  wire  x605; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 260:24:@46123.4]
  wire [31:0] _T_776; // @[Math.scala 406:49:@46132.4]
  wire [31:0] _T_778; // @[Math.scala 406:56:@46134.4]
  wire [31:0] _T_779; // @[Math.scala 406:56:@46135.4]
  wire  _T_784; // @[FixedPoint.scala 50:25:@46141.4]
  wire [1:0] _T_788; // @[Bitwise.scala 72:12:@46143.4]
  wire [29:0] _T_789; // @[FixedPoint.scala 18:52:@46144.4]
  wire  _T_824; // @[package.scala 96:25:@46214.4 package.scala 96:25:@46215.4]
  wire  _T_826; // @[implicits.scala 55:10:@46216.4]
  wire  _T_827; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 283:194:@46217.4]
  wire  x1088_x606_D1; // @[package.scala 96:25:@46182.4 package.scala 96:25:@46183.4]
  wire  _T_828; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 283:282:@46218.4]
  wire  x1089_b522_D13; // @[package.scala 96:25:@46191.4 package.scala 96:25:@46192.4]
  wire  _T_829; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 283:291:@46219.4]
  wire  x1087_b523_D13; // @[package.scala 96:25:@46173.4 package.scala 96:25:@46174.4]
  wire [31:0] x1091_x554_rdcol_D11_number; // @[package.scala 96:25:@46235.4 package.scala 96:25:@46236.4]
  wire [31:0] _T_840; // @[Math.scala 465:37:@46241.4]
  wire  x615; // @[Math.scala 465:44:@46243.4]
  wire  x616; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 291:24:@46246.4]
  wire  _T_871; // @[package.scala 96:25:@46290.4 package.scala 96:25:@46291.4]
  wire  _T_873; // @[implicits.scala 55:10:@46292.4]
  wire  _T_874; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 310:194:@46293.4]
  wire  x1093_x617_D1; // @[package.scala 96:25:@46276.4 package.scala 96:25:@46277.4]
  wire  _T_875; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 310:282:@46294.4]
  wire  _T_876; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 310:291:@46295.4]
  wire [31:0] x1094_x545_rdcol_D11_number; // @[package.scala 96:25:@46311.4 package.scala 96:25:@46312.4]
  wire [31:0] _T_889; // @[Math.scala 465:37:@46319.4]
  wire  x623; // @[Math.scala 465:44:@46321.4]
  wire  x624; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 320:59:@46324.4]
  wire  _T_920; // @[package.scala 96:25:@46368.4 package.scala 96:25:@46369.4]
  wire  _T_922; // @[implicits.scala 55:10:@46370.4]
  wire  _T_923; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 333:194:@46371.4]
  wire  x1096_x625_D1; // @[package.scala 96:25:@46354.4 package.scala 96:25:@46355.4]
  wire  _T_924; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 333:282:@46372.4]
  wire  _T_925; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 333:291:@46373.4]
  wire [31:0] x1097_b521_D11_number; // @[package.scala 96:25:@46389.4 package.scala 96:25:@46390.4]
  wire [31:0] _T_936; // @[Math.scala 465:37:@46395.4]
  wire  x631; // @[Math.scala 465:44:@46397.4]
  wire  x1098_x631_D1; // @[package.scala 96:25:@46405.4 package.scala 96:25:@46406.4]
  wire  x632; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 343:59:@46409.4]
  wire  _T_970; // @[package.scala 96:25:@46453.4 package.scala 96:25:@46454.4]
  wire  _T_972; // @[implicits.scala 55:10:@46455.4]
  wire  _T_973; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 356:194:@46456.4]
  wire  x1100_x633_D1; // @[package.scala 96:25:@46439.4 package.scala 96:25:@46440.4]
  wire  _T_974; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 356:282:@46457.4]
  wire  _T_975; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 356:291:@46458.4]
  wire [31:0] x639_rdcol_number; // @[Math.scala 154:22:@46477.4 Math.scala 155:14:@46478.4]
  wire [31:0] _T_990; // @[Math.scala 465:37:@46483.4]
  wire  x640; // @[Math.scala 465:44:@46485.4]
  wire  x641; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 364:59:@46488.4]
  wire  _T_1000; // @[FixedPoint.scala 50:25:@46495.4]
  wire [1:0] _T_1004; // @[Bitwise.scala 72:12:@46497.4]
  wire [29:0] _T_1005; // @[FixedPoint.scala 18:52:@46498.4]
  wire  _T_1028; // @[package.scala 96:25:@46532.4 package.scala 96:25:@46533.4]
  wire  _T_1030; // @[implicits.scala 55:10:@46534.4]
  wire  _T_1031; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 377:194:@46535.4]
  wire  x1101_x642_D1; // @[package.scala 96:25:@46518.4 package.scala 96:25:@46519.4]
  wire  _T_1032; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 377:282:@46536.4]
  wire  _T_1033; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 377:291:@46537.4]
  wire [31:0] x651_rdcol_number; // @[Math.scala 154:22:@46556.4 Math.scala 155:14:@46557.4]
  wire [31:0] _T_1048; // @[Math.scala 465:37:@46562.4]
  wire  x652; // @[Math.scala 465:44:@46564.4]
  wire  x653; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 385:59:@46567.4]
  wire  _T_1058; // @[FixedPoint.scala 50:25:@46574.4]
  wire [1:0] _T_1062; // @[Bitwise.scala 72:12:@46576.4]
  wire [29:0] _T_1063; // @[FixedPoint.scala 18:52:@46577.4]
  wire  _T_1086; // @[package.scala 96:25:@46611.4 package.scala 96:25:@46612.4]
  wire  _T_1088; // @[implicits.scala 55:10:@46613.4]
  wire  _T_1089; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 398:194:@46614.4]
  wire  x1102_x654_D1; // @[package.scala 96:25:@46597.4 package.scala 96:25:@46598.4]
  wire  _T_1090; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 398:282:@46615.4]
  wire  _T_1091; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 398:291:@46616.4]
  wire [31:0] x1103_b520_D11_number; // @[package.scala 96:25:@46632.4 package.scala 96:25:@46633.4]
  wire [31:0] _T_1104; // @[Math.scala 406:49:@46639.4]
  wire [31:0] _T_1106; // @[Math.scala 406:56:@46641.4]
  wire [31:0] _T_1107; // @[Math.scala 406:56:@46642.4]
  wire [31:0] x1055_number; // @[implicits.scala 133:21:@46643.4]
  wire  x664; // @[Math.scala 465:44:@46651.4]
  wire  x1104_x664_D1; // @[package.scala 96:25:@46659.4 package.scala 96:25:@46660.4]
  wire  x665; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 410:25:@46663.4]
  wire [31:0] _T_1131; // @[Math.scala 406:49:@46672.4]
  wire [31:0] _T_1133; // @[Math.scala 406:56:@46674.4]
  wire [31:0] _T_1134; // @[Math.scala 406:56:@46675.4]
  wire  _T_1139; // @[FixedPoint.scala 50:25:@46681.4]
  wire [1:0] _T_1143; // @[Bitwise.scala 72:12:@46683.4]
  wire [29:0] _T_1144; // @[FixedPoint.scala 18:52:@46684.4]
  wire  _T_1175; // @[package.scala 96:25:@46738.4 package.scala 96:25:@46739.4]
  wire  _T_1177; // @[implicits.scala 55:10:@46740.4]
  wire  _T_1178; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 437:194:@46741.4]
  wire  x1106_x666_D1; // @[package.scala 96:25:@46715.4 package.scala 96:25:@46716.4]
  wire  _T_1179; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 437:282:@46742.4]
  wire  _T_1180; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 437:291:@46743.4]
  wire  x675; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 441:60:@46754.4]
  wire  _T_1208; // @[package.scala 96:25:@46789.4 package.scala 96:25:@46790.4]
  wire  _T_1210; // @[implicits.scala 55:10:@46791.4]
  wire  _T_1211; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 452:194:@46792.4]
  wire  x1108_x676_D1; // @[package.scala 96:25:@46775.4 package.scala 96:25:@46776.4]
  wire  _T_1212; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 452:282:@46793.4]
  wire  _T_1213; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 452:291:@46794.4]
  wire  x682; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 456:60:@46805.4]
  wire  _T_1241; // @[package.scala 96:25:@46840.4 package.scala 96:25:@46841.4]
  wire  _T_1243; // @[implicits.scala 55:10:@46842.4]
  wire  _T_1244; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 467:194:@46843.4]
  wire  x1109_x683_D1; // @[package.scala 96:25:@46826.4 package.scala 96:25:@46827.4]
  wire  _T_1245; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 467:282:@46844.4]
  wire  _T_1246; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 467:291:@46845.4]
  wire  x689; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 471:59:@46856.4]
  wire  _T_1280; // @[package.scala 96:25:@46909.4 package.scala 96:25:@46910.4]
  wire  _T_1282; // @[implicits.scala 55:10:@46911.4]
  wire  _T_1283; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 486:194:@46912.4]
  wire  x1111_x690_D2; // @[package.scala 96:25:@46886.4 package.scala 96:25:@46887.4]
  wire  _T_1284; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 486:282:@46913.4]
  wire  _T_1285; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 486:291:@46914.4]
  wire  x696; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 490:60:@46925.4]
  wire  _T_1313; // @[package.scala 96:25:@46960.4 package.scala 96:25:@46961.4]
  wire  _T_1315; // @[implicits.scala 55:10:@46962.4]
  wire  _T_1316; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 501:194:@46963.4]
  wire  x1113_x697_D1; // @[package.scala 96:25:@46946.4 package.scala 96:25:@46947.4]
  wire  _T_1317; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 501:282:@46964.4]
  wire  _T_1318; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 501:291:@46965.4]
  wire  x703; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 505:60:@46976.4]
  wire  _T_1346; // @[package.scala 96:25:@47011.4 package.scala 96:25:@47012.4]
  wire  _T_1348; // @[implicits.scala 55:10:@47013.4]
  wire  _T_1349; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 516:194:@47014.4]
  wire  x1114_x704_D1; // @[package.scala 96:25:@46997.4 package.scala 96:25:@46998.4]
  wire  _T_1350; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 516:282:@47015.4]
  wire  _T_1351; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 516:291:@47016.4]
  wire [31:0] x710_rdrow_number; // @[Math.scala 154:22:@47035.4 Math.scala 155:14:@47036.4]
  wire [31:0] _T_1368; // @[Math.scala 406:49:@47042.4]
  wire [31:0] _T_1370; // @[Math.scala 406:56:@47044.4]
  wire [31:0] _T_1371; // @[Math.scala 406:56:@47045.4]
  wire [31:0] x1057_number; // @[implicits.scala 133:21:@47046.4]
  wire  x712; // @[Math.scala 465:44:@47054.4]
  wire  x713; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 526:24:@47057.4]
  wire [31:0] _T_1392; // @[Math.scala 406:49:@47066.4]
  wire [31:0] _T_1394; // @[Math.scala 406:56:@47068.4]
  wire [31:0] _T_1395; // @[Math.scala 406:56:@47069.4]
  wire  _T_1400; // @[FixedPoint.scala 50:25:@47075.4]
  wire [1:0] _T_1404; // @[Bitwise.scala 72:12:@47077.4]
  wire [29:0] _T_1405; // @[FixedPoint.scala 18:52:@47078.4]
  wire  _T_1431; // @[package.scala 96:25:@47121.4 package.scala 96:25:@47122.4]
  wire  _T_1433; // @[implicits.scala 55:10:@47123.4]
  wire  _T_1434; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 543:194:@47124.4]
  wire  x1115_x714_D1; // @[package.scala 96:25:@47098.4 package.scala 96:25:@47099.4]
  wire  _T_1435; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 543:282:@47125.4]
  wire  _T_1436; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 543:291:@47126.4]
  wire  x723; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 553:59:@47137.4]
  wire  _T_1466; // @[package.scala 96:25:@47174.4 package.scala 96:25:@47175.4]
  wire  _T_1468; // @[implicits.scala 55:10:@47176.4]
  wire  _T_1469; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 566:194:@47177.4]
  wire  x1117_x724_D1; // @[package.scala 96:25:@47160.4 package.scala 96:25:@47161.4]
  wire  _T_1470; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 566:282:@47178.4]
  wire  _T_1471; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 566:291:@47179.4]
  wire  x730; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 570:59:@47190.4]
  wire  _T_1499; // @[package.scala 96:25:@47225.4 package.scala 96:25:@47226.4]
  wire  _T_1501; // @[implicits.scala 55:10:@47227.4]
  wire  _T_1502; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 581:194:@47228.4]
  wire  x1118_x731_D1; // @[package.scala 96:25:@47211.4 package.scala 96:25:@47212.4]
  wire  _T_1503; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 581:282:@47229.4]
  wire  _T_1504; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 581:291:@47230.4]
  wire  x737; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 585:59:@47241.4]
  wire  _T_1532; // @[package.scala 96:25:@47276.4 package.scala 96:25:@47277.4]
  wire  _T_1534; // @[implicits.scala 55:10:@47278.4]
  wire  _T_1535; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 596:194:@47279.4]
  wire  x1119_x738_D1; // @[package.scala 96:25:@47262.4 package.scala 96:25:@47263.4]
  wire  _T_1536; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 596:282:@47280.4]
  wire  _T_1537; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 596:291:@47281.4]
  wire  x744; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 600:59:@47292.4]
  wire  _T_1565; // @[package.scala 96:25:@47327.4 package.scala 96:25:@47328.4]
  wire  _T_1567; // @[implicits.scala 55:10:@47329.4]
  wire  _T_1568; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 611:194:@47330.4]
  wire  x1120_x745_D1; // @[package.scala 96:25:@47313.4 package.scala 96:25:@47314.4]
  wire  _T_1569; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 611:282:@47331.4]
  wire  _T_1570; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 611:291:@47332.4]
  wire  x751; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 615:59:@47343.4]
  wire  _T_1598; // @[package.scala 96:25:@47378.4 package.scala 96:25:@47379.4]
  wire  _T_1600; // @[implicits.scala 55:10:@47380.4]
  wire  _T_1601; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 626:194:@47381.4]
  wire  x1121_x752_D1; // @[package.scala 96:25:@47364.4 package.scala 96:25:@47365.4]
  wire  _T_1602; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 626:282:@47382.4]
  wire  _T_1603; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 626:291:@47383.4]
  wire [31:0] x758_rdrow_number; // @[Math.scala 154:22:@47402.4 Math.scala 155:14:@47403.4]
  wire [31:0] _T_1620; // @[Math.scala 406:49:@47409.4]
  wire [31:0] _T_1622; // @[Math.scala 406:56:@47411.4]
  wire [31:0] _T_1623; // @[Math.scala 406:56:@47412.4]
  wire [31:0] x1059_number; // @[implicits.scala 133:21:@47413.4]
  wire  x760; // @[Math.scala 465:44:@47421.4]
  wire  x761; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 636:24:@47424.4]
  wire [31:0] _T_1644; // @[Math.scala 406:49:@47433.4]
  wire [31:0] _T_1646; // @[Math.scala 406:56:@47435.4]
  wire [31:0] _T_1647; // @[Math.scala 406:56:@47436.4]
  wire  _T_1652; // @[FixedPoint.scala 50:25:@47442.4]
  wire [1:0] _T_1656; // @[Bitwise.scala 72:12:@47444.4]
  wire [29:0] _T_1657; // @[FixedPoint.scala 18:52:@47445.4]
  wire  _T_1683; // @[package.scala 96:25:@47488.4 package.scala 96:25:@47489.4]
  wire  _T_1685; // @[implicits.scala 55:10:@47490.4]
  wire  _T_1686; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 653:194:@47491.4]
  wire  x1122_x762_D1; // @[package.scala 96:25:@47465.4 package.scala 96:25:@47466.4]
  wire  _T_1687; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 653:282:@47492.4]
  wire  _T_1688; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 653:291:@47493.4]
  wire  x771; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 657:24:@47504.4]
  wire  _T_1716; // @[package.scala 96:25:@47539.4 package.scala 96:25:@47540.4]
  wire  _T_1718; // @[implicits.scala 55:10:@47541.4]
  wire  _T_1719; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 668:194:@47542.4]
  wire  x1124_x772_D1; // @[package.scala 96:25:@47525.4 package.scala 96:25:@47526.4]
  wire  _T_1720; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 668:282:@47543.4]
  wire  _T_1721; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 668:291:@47544.4]
  wire  x778; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 672:24:@47555.4]
  wire  _T_1751; // @[package.scala 96:25:@47592.4 package.scala 96:25:@47593.4]
  wire  _T_1753; // @[implicits.scala 55:10:@47594.4]
  wire  _T_1754; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 691:194:@47595.4]
  wire  x1125_x779_D1; // @[package.scala 96:25:@47578.4 package.scala 96:25:@47579.4]
  wire  _T_1755; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 691:282:@47596.4]
  wire  _T_1756; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 691:291:@47597.4]
  wire  x785; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 695:59:@47608.4]
  wire  _T_1784; // @[package.scala 96:25:@47643.4 package.scala 96:25:@47644.4]
  wire  _T_1786; // @[implicits.scala 55:10:@47645.4]
  wire  _T_1787; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 706:194:@47646.4]
  wire  x1126_x786_D1; // @[package.scala 96:25:@47629.4 package.scala 96:25:@47630.4]
  wire  _T_1788; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 706:282:@47647.4]
  wire  _T_1789; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 706:291:@47648.4]
  wire  x792; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 710:59:@47659.4]
  wire  _T_1817; // @[package.scala 96:25:@47694.4 package.scala 96:25:@47695.4]
  wire  _T_1819; // @[implicits.scala 55:10:@47696.4]
  wire  _T_1820; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 721:194:@47697.4]
  wire  x1127_x793_D1; // @[package.scala 96:25:@47680.4 package.scala 96:25:@47681.4]
  wire  _T_1821; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 721:282:@47698.4]
  wire  _T_1822; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 721:291:@47699.4]
  wire  x799; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 725:59:@47710.4]
  wire  _T_1850; // @[package.scala 96:25:@47745.4 package.scala 96:25:@47746.4]
  wire  _T_1852; // @[implicits.scala 55:10:@47747.4]
  wire  _T_1853; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 736:194:@47748.4]
  wire  x1128_x800_D1; // @[package.scala 96:25:@47731.4 package.scala 96:25:@47732.4]
  wire  _T_1854; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 736:282:@47749.4]
  wire  _T_1855; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 736:291:@47750.4]
  wire [7:0] x621_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 306:29:@46279.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 310:410:@46302.4]
  wire [8:0] _GEN_0; // @[Math.scala 450:32:@47762.4]
  wire [8:0] _T_1861; // @[Math.scala 450:32:@47762.4]
  wire [7:0] x673_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 433:29:@46727.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 437:410:@46750.4]
  wire [8:0] _GEN_1; // @[Math.scala 450:32:@47767.4]
  wire [8:0] _T_1865; // @[Math.scala 450:32:@47767.4]
  wire [7:0] x680_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 448:29:@46778.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 452:410:@46801.4]
  wire [9:0] _GEN_2; // @[Math.scala 450:32:@47772.4]
  wire [9:0] _T_1869; // @[Math.scala 450:32:@47772.4]
  wire [7:0] x687_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 463:29:@46829.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 467:410:@46852.4]
  wire [8:0] _GEN_3; // @[Math.scala 450:32:@47777.4]
  wire [8:0] _T_1873; // @[Math.scala 450:32:@47777.4]
  wire [7:0] x728_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 562:29:@47163.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 566:410:@47186.4]
  wire [8:0] _GEN_4; // @[Math.scala 450:32:@47782.4]
  wire [8:0] _T_1877; // @[Math.scala 450:32:@47782.4]
  wire [7:0] x818_sum_number; // @[Math.scala 154:22:@47871.4 Math.scala 155:14:@47872.4]
  wire [3:0] _T_1913; // @[FixedPoint.scala 18:52:@47877.4]
  wire [7:0] x629_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 329:29:@46357.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 333:410:@46380.4]
  wire [8:0] _GEN_5; // @[Math.scala 450:32:@47890.4]
  wire [8:0] _T_1920; // @[Math.scala 450:32:@47890.4]
  wire [8:0] _GEN_6; // @[Math.scala 450:32:@47895.4]
  wire [8:0] _T_1924; // @[Math.scala 450:32:@47895.4]
  wire [9:0] _GEN_7; // @[Math.scala 450:32:@47900.4]
  wire [9:0] _T_1928; // @[Math.scala 450:32:@47900.4]
  wire [7:0] x694_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 482:29:@46898.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 486:410:@46921.4]
  wire [8:0] _GEN_8; // @[Math.scala 450:32:@47905.4]
  wire [8:0] _T_1932; // @[Math.scala 450:32:@47905.4]
  wire [7:0] x735_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 577:29:@47214.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 581:410:@47237.4]
  wire [8:0] _GEN_9; // @[Math.scala 450:32:@47910.4]
  wire [8:0] _T_1936; // @[Math.scala 450:32:@47910.4]
  wire [7:0] x832_sum_number; // @[Math.scala 154:22:@48001.4 Math.scala 155:14:@48002.4]
  wire [3:0] _T_1974; // @[FixedPoint.scala 18:52:@48007.4]
  wire [7:0] x637_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 352:29:@46442.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 356:410:@46465.4]
  wire [8:0] _GEN_10; // @[Math.scala 450:32:@48020.4]
  wire [8:0] _T_1981; // @[Math.scala 450:32:@48020.4]
  wire [9:0] _GEN_11; // @[Math.scala 450:32:@48025.4]
  wire [9:0] _T_1985; // @[Math.scala 450:32:@48025.4]
  wire [7:0] x701_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 497:29:@46949.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 501:410:@46972.4]
  wire [8:0] _GEN_12; // @[Math.scala 450:32:@48030.4]
  wire [8:0] _T_1989; // @[Math.scala 450:32:@48030.4]
  wire [7:0] x742_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 592:29:@47265.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 596:410:@47288.4]
  wire [8:0] _GEN_13; // @[Math.scala 450:32:@48035.4]
  wire [8:0] _T_1993; // @[Math.scala 450:32:@48035.4]
  wire [7:0] x845_sum_number; // @[Math.scala 154:22:@48124.4 Math.scala 155:14:@48125.4]
  wire [3:0] _T_2029; // @[FixedPoint.scala 18:52:@48130.4]
  wire [7:0] x649_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 373:29:@46521.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 377:410:@46544.4]
  wire [8:0] _GEN_14; // @[Math.scala 450:32:@48143.4]
  wire [8:0] _T_2036; // @[Math.scala 450:32:@48143.4]
  wire [9:0] _GEN_15; // @[Math.scala 450:32:@48148.4]
  wire [9:0] _T_2040; // @[Math.scala 450:32:@48148.4]
  wire [7:0] x708_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 512:29:@47000.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 516:410:@47023.4]
  wire [8:0] _GEN_16; // @[Math.scala 450:32:@48153.4]
  wire [8:0] _T_2044; // @[Math.scala 450:32:@48153.4]
  wire [7:0] x749_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 607:29:@47316.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 611:410:@47339.4]
  wire [8:0] _GEN_17; // @[Math.scala 450:32:@48158.4]
  wire [8:0] _T_2048; // @[Math.scala 450:32:@48158.4]
  wire [7:0] x858_sum_number; // @[Math.scala 154:22:@48247.4 Math.scala 155:14:@48248.4]
  wire [3:0] _T_2084; // @[FixedPoint.scala 18:52:@48253.4]
  wire [7:0] x721_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 539:29:@47110.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 543:410:@47133.4]
  wire [8:0] _GEN_18; // @[Math.scala 450:32:@48266.4]
  wire [8:0] _T_2091; // @[Math.scala 450:32:@48266.4]
  wire [9:0] _GEN_19; // @[Math.scala 450:32:@48271.4]
  wire [9:0] _T_2095; // @[Math.scala 450:32:@48271.4]
  wire [7:0] x776_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 664:29:@47528.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 668:410:@47551.4]
  wire [8:0] _GEN_20; // @[Math.scala 450:32:@48276.4]
  wire [8:0] _T_2099; // @[Math.scala 450:32:@48276.4]
  wire [7:0] x870_sum_number; // @[Math.scala 154:22:@48365.4 Math.scala 155:14:@48366.4]
  wire [3:0] _T_2135; // @[FixedPoint.scala 18:52:@48371.4]
  wire [9:0] _GEN_21; // @[Math.scala 450:32:@48384.4]
  wire [9:0] _T_2142; // @[Math.scala 450:32:@48384.4]
  wire [7:0] x783_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 687:29:@47581.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 691:410:@47604.4]
  wire [8:0] _GEN_22; // @[Math.scala 450:32:@48389.4]
  wire [8:0] _T_2146; // @[Math.scala 450:32:@48389.4]
  wire [7:0] x881_sum_number; // @[Math.scala 154:22:@48480.4 Math.scala 155:14:@48481.4]
  wire [3:0] _T_2184; // @[FixedPoint.scala 18:52:@48486.4]
  wire [9:0] _GEN_23; // @[Math.scala 450:32:@48499.4]
  wire [9:0] _T_2191; // @[Math.scala 450:32:@48499.4]
  wire [7:0] x790_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 702:29:@47632.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 706:410:@47655.4]
  wire [8:0] _GEN_24; // @[Math.scala 450:32:@48504.4]
  wire [8:0] _T_2195; // @[Math.scala 450:32:@48504.4]
  wire [7:0] x892_sum_number; // @[Math.scala 154:22:@48593.4 Math.scala 155:14:@48594.4]
  wire [3:0] _T_2231; // @[FixedPoint.scala 18:52:@48599.4]
  wire [9:0] _GEN_25; // @[Math.scala 450:32:@48612.4]
  wire [9:0] _T_2238; // @[Math.scala 450:32:@48612.4]
  wire [7:0] x756_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 622:29:@47367.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 626:410:@47390.4]
  wire [8:0] _GEN_26; // @[Math.scala 450:32:@48617.4]
  wire [8:0] _T_2242; // @[Math.scala 450:32:@48617.4]
  wire [7:0] x797_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 717:29:@47683.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 721:410:@47706.4]
  wire [8:0] _GEN_27; // @[Math.scala 450:32:@48622.4]
  wire [8:0] _T_2246; // @[Math.scala 450:32:@48622.4]
  wire [7:0] x904_sum_number; // @[Math.scala 154:22:@48711.4 Math.scala 155:14:@48712.4]
  wire [3:0] _T_2282; // @[FixedPoint.scala 18:52:@48717.4]
  wire  _T_2310; // @[package.scala 96:25:@48783.4 package.scala 96:25:@48784.4]
  wire  _T_2312; // @[implicits.scala 55:10:@48785.4]
  wire  _T_2313; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 986:167:@48786.4]
  wire  _T_2315; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 986:255:@48788.4]
  wire  _T_2316; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 986:274:@48789.4]
  wire  x1140_b522_D18; // @[package.scala 96:25:@48761.4 package.scala 96:25:@48762.4]
  wire  _T_2317; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 986:300:@48790.4]
  wire  x1137_b523_D18; // @[package.scala 96:25:@48734.4 package.scala 96:25:@48735.4]
  wire  _T_2334; // @[package.scala 96:25:@48826.4 package.scala 96:25:@48827.4]
  wire  _T_2336; // @[implicits.scala 55:10:@48828.4]
  wire  _T_2337; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 995:167:@48829.4]
  wire  _T_2339; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 995:255:@48831.4]
  wire  _T_2340; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 995:274:@48832.4]
  wire  _T_2341; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 995:300:@48833.4]
  wire  _T_2358; // @[package.scala 96:25:@48869.4 package.scala 96:25:@48870.4]
  wire  _T_2360; // @[implicits.scala 55:10:@48871.4]
  wire  _T_2361; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1004:167:@48872.4]
  wire  _T_2363; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1004:255:@48874.4]
  wire  _T_2364; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1004:274:@48875.4]
  wire  _T_2365; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1004:300:@48876.4]
  wire  _T_2382; // @[package.scala 96:25:@48912.4 package.scala 96:25:@48913.4]
  wire  _T_2384; // @[implicits.scala 55:10:@48914.4]
  wire  _T_2385; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1013:167:@48915.4]
  wire  _T_2387; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1013:255:@48917.4]
  wire  _T_2388; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1013:274:@48918.4]
  wire  _T_2389; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1013:300:@48919.4]
  wire  _T_2409; // @[package.scala 96:25:@48964.4 package.scala 96:25:@48965.4]
  wire  _T_2411; // @[implicits.scala 55:10:@48966.4]
  wire  _T_2412; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1030:167:@48967.4]
  wire  _T_2414; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1030:255:@48969.4]
  wire  _T_2415; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1030:274:@48970.4]
  wire  _T_2416; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1030:300:@48971.4]
  wire  _T_2433; // @[package.scala 96:25:@49007.4 package.scala 96:25:@49008.4]
  wire  _T_2435; // @[implicits.scala 55:10:@49009.4]
  wire  _T_2436; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1039:167:@49010.4]
  wire  _T_2438; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1039:255:@49012.4]
  wire  _T_2439; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1039:274:@49013.4]
  wire  _T_2440; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1039:300:@49014.4]
  wire  _T_2457; // @[package.scala 96:25:@49050.4 package.scala 96:25:@49051.4]
  wire  _T_2459; // @[implicits.scala 55:10:@49052.4]
  wire  _T_2460; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1048:167:@49053.4]
  wire  _T_2462; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1048:255:@49055.4]
  wire  _T_2463; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1048:274:@49056.4]
  wire  _T_2464; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1048:300:@49057.4]
  wire  _T_2481; // @[package.scala 96:25:@49093.4 package.scala 96:25:@49094.4]
  wire  _T_2483; // @[implicits.scala 55:10:@49095.4]
  wire  _T_2484; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1057:167:@49096.4]
  wire  _T_2486; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1057:255:@49098.4]
  wire  _T_2487; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1057:274:@49099.4]
  wire  _T_2488; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1057:300:@49100.4]
  wire  _T_2520; // @[package.scala 96:25:@49164.4 package.scala 96:25:@49165.4]
  wire  _T_2522; // @[implicits.scala 55:10:@49166.4]
  wire  _T_2523; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1073:195:@49167.4]
  wire  x1158_x606_D7; // @[package.scala 96:25:@49123.4 package.scala 96:25:@49124.4]
  wire  _T_2524; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1073:283:@49168.4]
  wire  x1159_b522_D19; // @[package.scala 96:25:@49132.4 package.scala 96:25:@49133.4]
  wire  _T_2525; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1073:292:@49169.4]
  wire  x1157_b523_D19; // @[package.scala 96:25:@49114.4 package.scala 96:25:@49115.4]
  wire  _T_2549; // @[package.scala 96:25:@49208.4 package.scala 96:25:@49209.4]
  wire  _T_2551; // @[implicits.scala 55:10:@49210.4]
  wire  _T_2552; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1084:195:@49211.4]
  wire  x1163_x617_D7; // @[package.scala 96:25:@49194.4 package.scala 96:25:@49195.4]
  wire  _T_2553; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1084:283:@49212.4]
  wire  _T_2554; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1084:292:@49213.4]
  wire  _T_2578; // @[package.scala 96:25:@49252.4 package.scala 96:25:@49253.4]
  wire  _T_2580; // @[implicits.scala 55:10:@49254.4]
  wire  _T_2581; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1095:195:@49255.4]
  wire  x1164_x625_D7; // @[package.scala 96:25:@49229.4 package.scala 96:25:@49230.4]
  wire  _T_2582; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1095:283:@49256.4]
  wire  _T_2583; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1095:292:@49257.4]
  wire  _T_2607; // @[package.scala 96:25:@49296.4 package.scala 96:25:@49297.4]
  wire  _T_2609; // @[implicits.scala 55:10:@49298.4]
  wire  _T_2610; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1106:195:@49299.4]
  wire  x1167_x633_D7; // @[package.scala 96:25:@49282.4 package.scala 96:25:@49283.4]
  wire  _T_2611; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1106:283:@49300.4]
  wire  _T_2612; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1106:292:@49301.4]
  wire  _T_2636; // @[package.scala 96:25:@49340.4 package.scala 96:25:@49341.4]
  wire  _T_2638; // @[implicits.scala 55:10:@49342.4]
  wire  _T_2639; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1117:195:@49343.4]
  wire  x1169_x642_D7; // @[package.scala 96:25:@49326.4 package.scala 96:25:@49327.4]
  wire  _T_2640; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1117:283:@49344.4]
  wire  _T_2641; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1117:292:@49345.4]
  wire  _T_2668; // @[package.scala 96:25:@49393.4 package.scala 96:25:@49394.4]
  wire  _T_2670; // @[implicits.scala 55:10:@49395.4]
  wire  _T_2671; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1130:195:@49396.4]
  wire  x1170_x666_D7; // @[package.scala 96:25:@49361.4 package.scala 96:25:@49362.4]
  wire  _T_2672; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1130:283:@49397.4]
  wire  _T_2673; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1130:292:@49398.4]
  wire  _T_2697; // @[package.scala 96:25:@49437.4 package.scala 96:25:@49438.4]
  wire  _T_2699; // @[implicits.scala 55:10:@49439.4]
  wire  _T_2700; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1141:195:@49440.4]
  wire  x1174_x676_D7; // @[package.scala 96:25:@49423.4 package.scala 96:25:@49424.4]
  wire  _T_2701; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1141:283:@49441.4]
  wire  _T_2702; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1141:292:@49442.4]
  wire  _T_2726; // @[package.scala 96:25:@49481.4 package.scala 96:25:@49482.4]
  wire  _T_2728; // @[implicits.scala 55:10:@49483.4]
  wire  _T_2729; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1152:195:@49484.4]
  wire  x1175_x683_D7; // @[package.scala 96:25:@49458.4 package.scala 96:25:@49459.4]
  wire  _T_2730; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1152:283:@49485.4]
  wire  _T_2731; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1152:292:@49486.4]
  wire  _T_2755; // @[package.scala 96:25:@49525.4 package.scala 96:25:@49526.4]
  wire  _T_2757; // @[implicits.scala 55:10:@49527.4]
  wire  _T_2758; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1169:195:@49528.4]
  wire  x1177_x690_D8; // @[package.scala 96:25:@49502.4 package.scala 96:25:@49503.4]
  wire  _T_2759; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1169:283:@49529.4]
  wire  _T_2760; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1169:292:@49530.4]
  wire  _T_2784; // @[package.scala 96:25:@49569.4 package.scala 96:25:@49570.4]
  wire  _T_2786; // @[implicits.scala 55:10:@49571.4]
  wire  _T_2787; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1180:195:@49572.4]
  wire  x1180_x697_D7; // @[package.scala 96:25:@49555.4 package.scala 96:25:@49556.4]
  wire  _T_2788; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1180:283:@49573.4]
  wire  _T_2789; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1180:292:@49574.4]
  wire  _T_2816; // @[package.scala 96:25:@49622.4 package.scala 96:25:@49623.4]
  wire  _T_2818; // @[implicits.scala 55:10:@49624.4]
  wire  _T_2819; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1193:195:@49625.4]
  wire  x1181_x714_D7; // @[package.scala 96:25:@49590.4 package.scala 96:25:@49591.4]
  wire  _T_2820; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1193:283:@49626.4]
  wire  _T_2821; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1193:292:@49627.4]
  wire  _T_2845; // @[package.scala 96:25:@49666.4 package.scala 96:25:@49667.4]
  wire  _T_2847; // @[implicits.scala 55:10:@49668.4]
  wire  _T_2848; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1204:195:@49669.4]
  wire  x1184_x724_D7; // @[package.scala 96:25:@49643.4 package.scala 96:25:@49644.4]
  wire  _T_2849; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1204:283:@49670.4]
  wire  _T_2850; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1204:292:@49671.4]
  wire  _T_2874; // @[package.scala 96:25:@49710.4 package.scala 96:25:@49711.4]
  wire  _T_2876; // @[implicits.scala 55:10:@49712.4]
  wire  _T_2877; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1215:195:@49713.4]
  wire  x1187_x731_D7; // @[package.scala 96:25:@49696.4 package.scala 96:25:@49697.4]
  wire  _T_2878; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1215:283:@49714.4]
  wire  _T_2879; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1215:292:@49715.4]
  wire  _T_2903; // @[package.scala 96:25:@49754.4 package.scala 96:25:@49755.4]
  wire  _T_2905; // @[implicits.scala 55:10:@49756.4]
  wire  _T_2906; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1226:195:@49757.4]
  wire  x1188_x738_D7; // @[package.scala 96:25:@49731.4 package.scala 96:25:@49732.4]
  wire  _T_2907; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1226:283:@49758.4]
  wire  _T_2908; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1226:292:@49759.4]
  wire  _T_2932; // @[package.scala 96:25:@49798.4 package.scala 96:25:@49799.4]
  wire  _T_2934; // @[implicits.scala 55:10:@49800.4]
  wire  _T_2935; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1237:195:@49801.4]
  wire  x1191_x745_D7; // @[package.scala 96:25:@49784.4 package.scala 96:25:@49785.4]
  wire  _T_2936; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1237:283:@49802.4]
  wire  _T_2937; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1237:292:@49803.4]
  wire [7:0] x918_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1080:29:@49197.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1084:341:@49220.4]
  wire [8:0] _GEN_28; // @[Math.scala 450:32:@49817.4]
  wire [8:0] _T_2945; // @[Math.scala 450:32:@49817.4]
  wire [7:0] x926_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1126:29:@49382.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1130:341:@49405.4]
  wire [8:0] _GEN_29; // @[Math.scala 450:32:@49822.4]
  wire [8:0] _T_2949; // @[Math.scala 450:32:@49822.4]
  wire [7:0] x920_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1091:29:@49241.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1095:341:@49264.4]
  wire [8:0] _GEN_30; // @[Math.scala 450:32:@49869.4]
  wire [8:0] _T_2969; // @[Math.scala 450:32:@49869.4]
  wire [7:0] x928_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1137:29:@49426.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1141:341:@49449.4]
  wire [8:0] _GEN_31; // @[Math.scala 450:32:@49874.4]
  wire [8:0] _T_2973; // @[Math.scala 450:32:@49874.4]
  wire [7:0] x922_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1102:29:@49285.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1106:341:@49308.4]
  wire [8:0] _GEN_32; // @[Math.scala 450:32:@49921.4]
  wire [8:0] _T_2993; // @[Math.scala 450:32:@49921.4]
  wire [7:0] x930_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1148:29:@49470.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1152:341:@49493.4]
  wire [8:0] _GEN_33; // @[Math.scala 450:32:@49926.4]
  wire [8:0] _T_2997; // @[Math.scala 450:32:@49926.4]
  wire [7:0] x924_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1113:29:@49329.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1117:341:@49352.4]
  wire [8:0] _GEN_34; // @[Math.scala 450:32:@49973.4]
  wire [8:0] _T_3017; // @[Math.scala 450:32:@49973.4]
  wire [7:0] x932_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1165:29:@49514.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1169:411:@49537.4]
  wire [8:0] _GEN_35; // @[Math.scala 450:32:@49980.4]
  wire [8:0] _T_3023; // @[Math.scala 450:32:@49980.4]
  wire [7:0] x936_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1189:29:@49611.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1193:411:@49634.4]
  wire [8:0] _GEN_36; // @[Math.scala 450:32:@50027.4]
  wire [8:0] _T_3043; // @[Math.scala 450:32:@50027.4]
  wire [7:0] x938_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1200:29:@49655.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1204:411:@49678.4]
  wire [8:0] _GEN_37; // @[Math.scala 450:32:@50074.4]
  wire [8:0] _T_3063; // @[Math.scala 450:32:@50074.4]
  wire [7:0] x940_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1211:29:@49699.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1215:411:@49722.4]
  wire [8:0] _GEN_38; // @[Math.scala 450:32:@50121.4]
  wire [8:0] _T_3083; // @[Math.scala 450:32:@50121.4]
  wire [7:0] x934_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1176:29:@49558.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1180:411:@49581.4]
  wire [8:0] _GEN_39; // @[Math.scala 450:32:@50168.4]
  wire [8:0] _T_3103; // @[Math.scala 450:32:@50168.4]
  wire [7:0] x942_rd_0_number; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1222:29:@49743.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1226:411:@49766.4]
  wire [8:0] _GEN_40; // @[Math.scala 450:32:@50173.4]
  wire [8:0] _T_3107; // @[Math.scala 450:32:@50173.4]
  wire [7:0] x984_div_number; // @[Math.scala 331:22:@50163.4 Math.scala 332:14:@50164.4]
  wire [7:0] x990_div_number; // @[Math.scala 331:22:@50215.4 Math.scala 332:14:@50216.4]
  wire [7:0] x974_div_number; // @[Math.scala 331:22:@50069.4 Math.scala 332:14:@50070.4]
  wire [7:0] x979_div_number; // @[Math.scala 331:22:@50116.4 Math.scala 332:14:@50117.4]
  wire [31:0] _T_3141; // @[Cat.scala 30:58:@50230.4]
  wire [7:0] x963_div_number; // @[Math.scala 331:22:@49968.4 Math.scala 332:14:@49969.4]
  wire [7:0] x969_div_number; // @[Math.scala 331:22:@50022.4 Math.scala 332:14:@50023.4]
  wire [7:0] x951_div_number; // @[Math.scala 331:22:@49864.4 Math.scala 332:14:@49865.4]
  wire [7:0] x957_div_number; // @[Math.scala 331:22:@49916.4 Math.scala 332:14:@49917.4]
  wire [31:0] _T_3144; // @[Cat.scala 30:58:@50233.4]
  wire  _T_3157; // @[package.scala 96:25:@50269.4 package.scala 96:25:@50270.4]
  wire  _T_3159; // @[implicits.scala 55:10:@50271.4]
  wire  x1192_b522_D29; // @[package.scala 96:25:@50251.4 package.scala 96:25:@50252.4]
  wire  _T_3160; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1349:116:@50272.4]
  wire  x1193_b523_D29; // @[package.scala 96:25:@50260.4 package.scala 96:25:@50261.4]
  wire  _T_3161; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1349:123:@50273.4]
  wire [31:0] x1063_x1051_D8_number; // @[package.scala 96:25:@45468.4 package.scala 96:25:@45469.4]
  wire [31:0] x1066_x539_sum_D7_number; // @[package.scala 96:25:@45495.4 package.scala 96:25:@45496.4]
  wire [31:0] x1069_x549_sum_D6_number; // @[package.scala 96:25:@45580.4 package.scala 96:25:@45581.4]
  wire [31:0] x1071_x558_sum_D6_number; // @[package.scala 96:25:@45656.4 package.scala 96:25:@45657.4]
  wire [31:0] x1072_x567_sum_D6_number; // @[package.scala 96:25:@45723.4 package.scala 96:25:@45724.4]
  wire [31:0] x1076_x1052_D7_number; // @[package.scala 96:25:@45877.4 package.scala 96:25:@45878.4]
  wire [31:0] x1077_x581_sum_D6_number; // @[package.scala 96:25:@45886.4 package.scala 96:25:@45887.4]
  wire [31:0] x1078_x587_sum_D6_number; // @[package.scala 96:25:@45932.4 package.scala 96:25:@45933.4]
  wire [31:0] x1081_x592_sum_D6_number; // @[package.scala 96:25:@45996.4 package.scala 96:25:@45997.4]
  wire [31:0] x1082_x597_sum_D6_number; // @[package.scala 96:25:@46042.4 package.scala 96:25:@46043.4]
  wire [31:0] x609_sum_number; // @[Math.scala 154:22:@46164.4 Math.scala 155:14:@46165.4]
  wire [31:0] x1090_x1054_D1_number; // @[package.scala 96:25:@46200.4 package.scala 96:25:@46201.4]
  wire [31:0] x618_sum_number; // @[Math.scala 154:22:@46267.4 Math.scala 155:14:@46268.4]
  wire [31:0] x626_sum_number; // @[Math.scala 154:22:@46345.4 Math.scala 155:14:@46346.4]
  wire [31:0] x634_sum_number; // @[Math.scala 154:22:@46430.4 Math.scala 155:14:@46431.4]
  wire [31:0] x645_sum_number; // @[Math.scala 154:22:@46509.4 Math.scala 155:14:@46510.4]
  wire [31:0] x657_sum_number; // @[Math.scala 154:22:@46588.4 Math.scala 155:14:@46589.4]
  wire [31:0] x669_sum_number; // @[Math.scala 154:22:@46706.4 Math.scala 155:14:@46707.4]
  wire [31:0] x1107_x1056_D2_number; // @[package.scala 96:25:@46724.4 package.scala 96:25:@46725.4]
  wire [31:0] x677_sum_number; // @[Math.scala 154:22:@46766.4 Math.scala 155:14:@46767.4]
  wire [31:0] x684_sum_number; // @[Math.scala 154:22:@46817.4 Math.scala 155:14:@46818.4]
  wire [31:0] x1112_x691_sum_D1_number; // @[package.scala 96:25:@46895.4 package.scala 96:25:@46896.4]
  wire [31:0] x698_sum_number; // @[Math.scala 154:22:@46937.4 Math.scala 155:14:@46938.4]
  wire [31:0] x705_sum_number; // @[Math.scala 154:22:@46988.4 Math.scala 155:14:@46989.4]
  wire [31:0] x717_sum_number; // @[Math.scala 154:22:@47089.4 Math.scala 155:14:@47090.4]
  wire [31:0] x1116_x1058_D1_number; // @[package.scala 96:25:@47107.4 package.scala 96:25:@47108.4]
  wire [31:0] x725_sum_number; // @[Math.scala 154:22:@47151.4 Math.scala 155:14:@47152.4]
  wire [31:0] x732_sum_number; // @[Math.scala 154:22:@47202.4 Math.scala 155:14:@47203.4]
  wire [31:0] x739_sum_number; // @[Math.scala 154:22:@47253.4 Math.scala 155:14:@47254.4]
  wire [31:0] x746_sum_number; // @[Math.scala 154:22:@47304.4 Math.scala 155:14:@47305.4]
  wire [31:0] x753_sum_number; // @[Math.scala 154:22:@47355.4 Math.scala 155:14:@47356.4]
  wire [31:0] x765_sum_number; // @[Math.scala 154:22:@47456.4 Math.scala 155:14:@47457.4]
  wire [31:0] x1123_x1060_D1_number; // @[package.scala 96:25:@47474.4 package.scala 96:25:@47475.4]
  wire [31:0] x773_sum_number; // @[Math.scala 154:22:@47516.4 Math.scala 155:14:@47517.4]
  wire [31:0] x780_sum_number; // @[Math.scala 154:22:@47569.4 Math.scala 155:14:@47570.4]
  wire [31:0] x787_sum_number; // @[Math.scala 154:22:@47620.4 Math.scala 155:14:@47621.4]
  wire [31:0] x794_sum_number; // @[Math.scala 154:22:@47671.4 Math.scala 155:14:@47672.4]
  wire [31:0] x801_sum_number; // @[Math.scala 154:22:@47722.4 Math.scala 155:14:@47723.4]
  wire [31:0] x1138_x1051_D18_number; // @[package.scala 96:25:@48743.4 package.scala 96:25:@48744.4]
  wire [31:0] x1141_x539_sum_D17_number; // @[package.scala 96:25:@48770.4 package.scala 96:25:@48771.4]
  wire [31:0] x1143_x549_sum_D16_number; // @[package.scala 96:25:@48813.4 package.scala 96:25:@48814.4]
  wire [31:0] x1144_x558_sum_D16_number; // @[package.scala 96:25:@48847.4 package.scala 96:25:@48848.4]
  wire [31:0] x1146_x567_sum_D16_number; // @[package.scala 96:25:@48890.4 package.scala 96:25:@48891.4]
  wire [31:0] x1148_x1052_D17_number; // @[package.scala 96:25:@48933.4 package.scala 96:25:@48934.4]
  wire [31:0] x1150_x581_sum_D16_number; // @[package.scala 96:25:@48951.4 package.scala 96:25:@48952.4]
  wire [31:0] x1152_x587_sum_D16_number; // @[package.scala 96:25:@48994.4 package.scala 96:25:@48995.4]
  wire [31:0] x1154_x592_sum_D16_number; // @[package.scala 96:25:@49037.4 package.scala 96:25:@49038.4]
  wire [31:0] x1155_x597_sum_D16_number; // @[package.scala 96:25:@49071.4 package.scala 96:25:@49072.4]
  wire [31:0] x1160_x1054_D7_number; // @[package.scala 96:25:@49141.4 package.scala 96:25:@49142.4]
  wire [31:0] x1161_x609_sum_D6_number; // @[package.scala 96:25:@49150.4 package.scala 96:25:@49151.4]
  wire [31:0] x1162_x618_sum_D6_number; // @[package.scala 96:25:@49185.4 package.scala 96:25:@49186.4]
  wire [31:0] x1165_x626_sum_D6_number; // @[package.scala 96:25:@49238.4 package.scala 96:25:@49239.4]
  wire [31:0] x1166_x634_sum_D6_number; // @[package.scala 96:25:@49273.4 package.scala 96:25:@49274.4]
  wire [31:0] x1168_x645_sum_D6_number; // @[package.scala 96:25:@49317.4 package.scala 96:25:@49318.4]
  wire [31:0] x1171_x669_sum_D6_number; // @[package.scala 96:25:@49370.4 package.scala 96:25:@49371.4]
  wire [31:0] x1172_x1056_D8_number; // @[package.scala 96:25:@49379.4 package.scala 96:25:@49380.4]
  wire [31:0] x1173_x677_sum_D6_number; // @[package.scala 96:25:@49414.4 package.scala 96:25:@49415.4]
  wire [31:0] x1176_x684_sum_D6_number; // @[package.scala 96:25:@49467.4 package.scala 96:25:@49468.4]
  wire [31:0] x1178_x691_sum_D7_number; // @[package.scala 96:25:@49511.4 package.scala 96:25:@49512.4]
  wire [31:0] x1179_x698_sum_D6_number; // @[package.scala 96:25:@49546.4 package.scala 96:25:@49547.4]
  wire [31:0] x1182_x1058_D7_number; // @[package.scala 96:25:@49599.4 package.scala 96:25:@49600.4]
  wire [31:0] x1183_x717_sum_D6_number; // @[package.scala 96:25:@49608.4 package.scala 96:25:@49609.4]
  wire [31:0] x1185_x725_sum_D6_number; // @[package.scala 96:25:@49652.4 package.scala 96:25:@49653.4]
  wire [31:0] x1186_x732_sum_D6_number; // @[package.scala 96:25:@49687.4 package.scala 96:25:@49688.4]
  wire [31:0] x1189_x739_sum_D6_number; // @[package.scala 96:25:@49740.4 package.scala 96:25:@49741.4]
  wire [31:0] x1190_x746_sum_D6_number; // @[package.scala 96:25:@49775.4 package.scala 96:25:@49776.4]
  _ _ ( // @[Math.scala 709:24:@44929.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@44941.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x524_lb_0 x524_lb_0 ( // @[m_x524_lb_0.scala 57:17:@44951.4]
    .clock(x524_lb_0_clock),
    .reset(x524_lb_0_reset),
    .io_rPort_23_banks_0(x524_lb_0_io_rPort_23_banks_0),
    .io_rPort_23_ofs_0(x524_lb_0_io_rPort_23_ofs_0),
    .io_rPort_23_en_0(x524_lb_0_io_rPort_23_en_0),
    .io_rPort_23_backpressure(x524_lb_0_io_rPort_23_backpressure),
    .io_rPort_23_output_0(x524_lb_0_io_rPort_23_output_0),
    .io_rPort_22_banks_0(x524_lb_0_io_rPort_22_banks_0),
    .io_rPort_22_ofs_0(x524_lb_0_io_rPort_22_ofs_0),
    .io_rPort_22_en_0(x524_lb_0_io_rPort_22_en_0),
    .io_rPort_22_backpressure(x524_lb_0_io_rPort_22_backpressure),
    .io_rPort_22_output_0(x524_lb_0_io_rPort_22_output_0),
    .io_rPort_21_banks_0(x524_lb_0_io_rPort_21_banks_0),
    .io_rPort_21_ofs_0(x524_lb_0_io_rPort_21_ofs_0),
    .io_rPort_21_en_0(x524_lb_0_io_rPort_21_en_0),
    .io_rPort_21_backpressure(x524_lb_0_io_rPort_21_backpressure),
    .io_rPort_21_output_0(x524_lb_0_io_rPort_21_output_0),
    .io_rPort_20_banks_0(x524_lb_0_io_rPort_20_banks_0),
    .io_rPort_20_ofs_0(x524_lb_0_io_rPort_20_ofs_0),
    .io_rPort_20_en_0(x524_lb_0_io_rPort_20_en_0),
    .io_rPort_20_backpressure(x524_lb_0_io_rPort_20_backpressure),
    .io_rPort_20_output_0(x524_lb_0_io_rPort_20_output_0),
    .io_rPort_19_banks_0(x524_lb_0_io_rPort_19_banks_0),
    .io_rPort_19_ofs_0(x524_lb_0_io_rPort_19_ofs_0),
    .io_rPort_19_en_0(x524_lb_0_io_rPort_19_en_0),
    .io_rPort_19_backpressure(x524_lb_0_io_rPort_19_backpressure),
    .io_rPort_19_output_0(x524_lb_0_io_rPort_19_output_0),
    .io_rPort_18_banks_0(x524_lb_0_io_rPort_18_banks_0),
    .io_rPort_18_ofs_0(x524_lb_0_io_rPort_18_ofs_0),
    .io_rPort_18_en_0(x524_lb_0_io_rPort_18_en_0),
    .io_rPort_18_backpressure(x524_lb_0_io_rPort_18_backpressure),
    .io_rPort_18_output_0(x524_lb_0_io_rPort_18_output_0),
    .io_rPort_17_banks_0(x524_lb_0_io_rPort_17_banks_0),
    .io_rPort_17_ofs_0(x524_lb_0_io_rPort_17_ofs_0),
    .io_rPort_17_en_0(x524_lb_0_io_rPort_17_en_0),
    .io_rPort_17_backpressure(x524_lb_0_io_rPort_17_backpressure),
    .io_rPort_17_output_0(x524_lb_0_io_rPort_17_output_0),
    .io_rPort_16_banks_0(x524_lb_0_io_rPort_16_banks_0),
    .io_rPort_16_ofs_0(x524_lb_0_io_rPort_16_ofs_0),
    .io_rPort_16_en_0(x524_lb_0_io_rPort_16_en_0),
    .io_rPort_16_backpressure(x524_lb_0_io_rPort_16_backpressure),
    .io_rPort_16_output_0(x524_lb_0_io_rPort_16_output_0),
    .io_rPort_15_banks_0(x524_lb_0_io_rPort_15_banks_0),
    .io_rPort_15_ofs_0(x524_lb_0_io_rPort_15_ofs_0),
    .io_rPort_15_en_0(x524_lb_0_io_rPort_15_en_0),
    .io_rPort_15_backpressure(x524_lb_0_io_rPort_15_backpressure),
    .io_rPort_15_output_0(x524_lb_0_io_rPort_15_output_0),
    .io_rPort_14_banks_0(x524_lb_0_io_rPort_14_banks_0),
    .io_rPort_14_ofs_0(x524_lb_0_io_rPort_14_ofs_0),
    .io_rPort_14_en_0(x524_lb_0_io_rPort_14_en_0),
    .io_rPort_14_backpressure(x524_lb_0_io_rPort_14_backpressure),
    .io_rPort_14_output_0(x524_lb_0_io_rPort_14_output_0),
    .io_rPort_13_banks_0(x524_lb_0_io_rPort_13_banks_0),
    .io_rPort_13_ofs_0(x524_lb_0_io_rPort_13_ofs_0),
    .io_rPort_13_en_0(x524_lb_0_io_rPort_13_en_0),
    .io_rPort_13_backpressure(x524_lb_0_io_rPort_13_backpressure),
    .io_rPort_13_output_0(x524_lb_0_io_rPort_13_output_0),
    .io_rPort_12_banks_0(x524_lb_0_io_rPort_12_banks_0),
    .io_rPort_12_ofs_0(x524_lb_0_io_rPort_12_ofs_0),
    .io_rPort_12_en_0(x524_lb_0_io_rPort_12_en_0),
    .io_rPort_12_backpressure(x524_lb_0_io_rPort_12_backpressure),
    .io_rPort_12_output_0(x524_lb_0_io_rPort_12_output_0),
    .io_rPort_11_banks_0(x524_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x524_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x524_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x524_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x524_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_0(x524_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x524_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x524_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x524_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x524_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_0(x524_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x524_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x524_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x524_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x524_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_0(x524_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x524_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x524_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x524_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x524_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_0(x524_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x524_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x524_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x524_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x524_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_0(x524_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x524_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x524_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x524_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x524_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_0(x524_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x524_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x524_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x524_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x524_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_0(x524_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x524_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x524_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x524_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x524_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_0(x524_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x524_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x524_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x524_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x524_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_0(x524_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x524_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x524_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x524_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x524_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_0(x524_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x524_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x524_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x524_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x524_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_0(x524_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x524_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x524_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x524_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x524_lb_0_io_rPort_0_output_0),
    .io_wPort_7_banks_0(x524_lb_0_io_wPort_7_banks_0),
    .io_wPort_7_ofs_0(x524_lb_0_io_wPort_7_ofs_0),
    .io_wPort_7_data_0(x524_lb_0_io_wPort_7_data_0),
    .io_wPort_7_en_0(x524_lb_0_io_wPort_7_en_0),
    .io_wPort_6_banks_0(x524_lb_0_io_wPort_6_banks_0),
    .io_wPort_6_ofs_0(x524_lb_0_io_wPort_6_ofs_0),
    .io_wPort_6_data_0(x524_lb_0_io_wPort_6_data_0),
    .io_wPort_6_en_0(x524_lb_0_io_wPort_6_en_0),
    .io_wPort_5_banks_0(x524_lb_0_io_wPort_5_banks_0),
    .io_wPort_5_ofs_0(x524_lb_0_io_wPort_5_ofs_0),
    .io_wPort_5_data_0(x524_lb_0_io_wPort_5_data_0),
    .io_wPort_5_en_0(x524_lb_0_io_wPort_5_en_0),
    .io_wPort_4_banks_0(x524_lb_0_io_wPort_4_banks_0),
    .io_wPort_4_ofs_0(x524_lb_0_io_wPort_4_ofs_0),
    .io_wPort_4_data_0(x524_lb_0_io_wPort_4_data_0),
    .io_wPort_4_en_0(x524_lb_0_io_wPort_4_en_0),
    .io_wPort_3_banks_0(x524_lb_0_io_wPort_3_banks_0),
    .io_wPort_3_ofs_0(x524_lb_0_io_wPort_3_ofs_0),
    .io_wPort_3_data_0(x524_lb_0_io_wPort_3_data_0),
    .io_wPort_3_en_0(x524_lb_0_io_wPort_3_en_0),
    .io_wPort_2_banks_0(x524_lb_0_io_wPort_2_banks_0),
    .io_wPort_2_ofs_0(x524_lb_0_io_wPort_2_ofs_0),
    .io_wPort_2_data_0(x524_lb_0_io_wPort_2_data_0),
    .io_wPort_2_en_0(x524_lb_0_io_wPort_2_en_0),
    .io_wPort_1_banks_0(x524_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x524_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x524_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x524_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_0(x524_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x524_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x524_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x524_lb_0_io_wPort_0_en_0)
  );
  x525_lb2_0 x525_lb2_0 ( // @[m_x525_lb2_0.scala 48:17:@45164.4]
    .clock(x525_lb2_0_clock),
    .reset(x525_lb2_0_reset),
    .io_rPort_14_banks_0(x525_lb2_0_io_rPort_14_banks_0),
    .io_rPort_14_ofs_0(x525_lb2_0_io_rPort_14_ofs_0),
    .io_rPort_14_en_0(x525_lb2_0_io_rPort_14_en_0),
    .io_rPort_14_backpressure(x525_lb2_0_io_rPort_14_backpressure),
    .io_rPort_14_output_0(x525_lb2_0_io_rPort_14_output_0),
    .io_rPort_13_banks_0(x525_lb2_0_io_rPort_13_banks_0),
    .io_rPort_13_ofs_0(x525_lb2_0_io_rPort_13_ofs_0),
    .io_rPort_13_en_0(x525_lb2_0_io_rPort_13_en_0),
    .io_rPort_13_backpressure(x525_lb2_0_io_rPort_13_backpressure),
    .io_rPort_13_output_0(x525_lb2_0_io_rPort_13_output_0),
    .io_rPort_12_banks_0(x525_lb2_0_io_rPort_12_banks_0),
    .io_rPort_12_ofs_0(x525_lb2_0_io_rPort_12_ofs_0),
    .io_rPort_12_en_0(x525_lb2_0_io_rPort_12_en_0),
    .io_rPort_12_backpressure(x525_lb2_0_io_rPort_12_backpressure),
    .io_rPort_12_output_0(x525_lb2_0_io_rPort_12_output_0),
    .io_rPort_11_banks_0(x525_lb2_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x525_lb2_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x525_lb2_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x525_lb2_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x525_lb2_0_io_rPort_11_output_0),
    .io_rPort_10_banks_0(x525_lb2_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x525_lb2_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x525_lb2_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x525_lb2_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x525_lb2_0_io_rPort_10_output_0),
    .io_rPort_9_banks_0(x525_lb2_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x525_lb2_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x525_lb2_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x525_lb2_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x525_lb2_0_io_rPort_9_output_0),
    .io_rPort_8_banks_0(x525_lb2_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x525_lb2_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x525_lb2_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x525_lb2_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x525_lb2_0_io_rPort_8_output_0),
    .io_rPort_7_banks_0(x525_lb2_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x525_lb2_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x525_lb2_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x525_lb2_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x525_lb2_0_io_rPort_7_output_0),
    .io_rPort_6_banks_0(x525_lb2_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x525_lb2_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x525_lb2_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x525_lb2_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x525_lb2_0_io_rPort_6_output_0),
    .io_rPort_5_banks_0(x525_lb2_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x525_lb2_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x525_lb2_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x525_lb2_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x525_lb2_0_io_rPort_5_output_0),
    .io_rPort_4_banks_0(x525_lb2_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x525_lb2_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x525_lb2_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x525_lb2_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x525_lb2_0_io_rPort_4_output_0),
    .io_rPort_3_banks_0(x525_lb2_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x525_lb2_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x525_lb2_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x525_lb2_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x525_lb2_0_io_rPort_3_output_0),
    .io_rPort_2_banks_0(x525_lb2_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x525_lb2_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x525_lb2_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x525_lb2_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x525_lb2_0_io_rPort_2_output_0),
    .io_rPort_1_banks_0(x525_lb2_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x525_lb2_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x525_lb2_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x525_lb2_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x525_lb2_0_io_rPort_1_output_0),
    .io_rPort_0_banks_0(x525_lb2_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x525_lb2_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x525_lb2_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x525_lb2_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x525_lb2_0_io_rPort_0_output_0),
    .io_wPort_7_banks_0(x525_lb2_0_io_wPort_7_banks_0),
    .io_wPort_7_ofs_0(x525_lb2_0_io_wPort_7_ofs_0),
    .io_wPort_7_data_0(x525_lb2_0_io_wPort_7_data_0),
    .io_wPort_7_en_0(x525_lb2_0_io_wPort_7_en_0),
    .io_wPort_6_banks_0(x525_lb2_0_io_wPort_6_banks_0),
    .io_wPort_6_ofs_0(x525_lb2_0_io_wPort_6_ofs_0),
    .io_wPort_6_data_0(x525_lb2_0_io_wPort_6_data_0),
    .io_wPort_6_en_0(x525_lb2_0_io_wPort_6_en_0),
    .io_wPort_5_banks_0(x525_lb2_0_io_wPort_5_banks_0),
    .io_wPort_5_ofs_0(x525_lb2_0_io_wPort_5_ofs_0),
    .io_wPort_5_data_0(x525_lb2_0_io_wPort_5_data_0),
    .io_wPort_5_en_0(x525_lb2_0_io_wPort_5_en_0),
    .io_wPort_4_banks_0(x525_lb2_0_io_wPort_4_banks_0),
    .io_wPort_4_ofs_0(x525_lb2_0_io_wPort_4_ofs_0),
    .io_wPort_4_data_0(x525_lb2_0_io_wPort_4_data_0),
    .io_wPort_4_en_0(x525_lb2_0_io_wPort_4_en_0),
    .io_wPort_3_banks_0(x525_lb2_0_io_wPort_3_banks_0),
    .io_wPort_3_ofs_0(x525_lb2_0_io_wPort_3_ofs_0),
    .io_wPort_3_data_0(x525_lb2_0_io_wPort_3_data_0),
    .io_wPort_3_en_0(x525_lb2_0_io_wPort_3_en_0),
    .io_wPort_2_banks_0(x525_lb2_0_io_wPort_2_banks_0),
    .io_wPort_2_ofs_0(x525_lb2_0_io_wPort_2_ofs_0),
    .io_wPort_2_data_0(x525_lb2_0_io_wPort_2_data_0),
    .io_wPort_2_en_0(x525_lb2_0_io_wPort_2_en_0),
    .io_wPort_1_banks_0(x525_lb2_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x525_lb2_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x525_lb2_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x525_lb2_0_io_wPort_1_en_0),
    .io_wPort_0_banks_0(x525_lb2_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x525_lb2_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x525_lb2_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x525_lb2_0_io_wPort_0_en_0)
  );
  RetimeWrapper_240 RetimeWrapper ( // @[package.scala 93:22:@45336.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x539_sum x539_sum_1 ( // @[Math.scala 150:24:@45444.4]
    .clock(x539_sum_1_clock),
    .reset(x539_sum_1_reset),
    .io_a(x539_sum_1_io_a),
    .io_b(x539_sum_1_io_b),
    .io_flow(x539_sum_1_io_flow),
    .io_result(x539_sum_1_io_result)
  );
  RetimeWrapper_242 RetimeWrapper_1 ( // @[package.scala 93:22:@45454.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_2 ( // @[package.scala 93:22:@45463.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_244 RetimeWrapper_3 ( // @[package.scala 93:22:@45472.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_242 RetimeWrapper_4 ( // @[package.scala 93:22:@45481.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_5 ( // @[package.scala 93:22:@45490.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_242 RetimeWrapper_6 ( // @[package.scala 93:22:@45503.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x539_sum x545_rdcol_1 ( // @[Math.scala 150:24:@45526.4]
    .clock(x545_rdcol_1_clock),
    .reset(x545_rdcol_1_reset),
    .io_a(x545_rdcol_1_io_a),
    .io_b(x545_rdcol_1_io_b),
    .io_flow(x545_rdcol_1_io_flow),
    .io_result(x545_rdcol_1_io_result)
  );
  RetimeWrapper_241 RetimeWrapper_7 ( // @[package.scala 93:22:@45547.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  x539_sum x549_sum_1 ( // @[Math.scala 150:24:@45556.4]
    .clock(x549_sum_1_clock),
    .reset(x549_sum_1_reset),
    .io_a(x549_sum_1_io_a),
    .io_b(x549_sum_1_io_b),
    .io_flow(x549_sum_1_io_flow),
    .io_result(x549_sum_1_io_result)
  );
  RetimeWrapper_244 RetimeWrapper_8 ( // @[package.scala 93:22:@45566.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_9 ( // @[package.scala 93:22:@45575.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_242 RetimeWrapper_10 ( // @[package.scala 93:22:@45588.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  x539_sum x554_rdcol_1 ( // @[Math.scala 150:24:@45611.4]
    .clock(x554_rdcol_1_clock),
    .reset(x554_rdcol_1_reset),
    .io_a(x554_rdcol_1_io_a),
    .io_b(x554_rdcol_1_io_b),
    .io_flow(x554_rdcol_1_io_flow),
    .io_result(x554_rdcol_1_io_result)
  );
  x539_sum x558_sum_1 ( // @[Math.scala 150:24:@45632.4]
    .clock(x558_sum_1_clock),
    .reset(x558_sum_1_reset),
    .io_a(x558_sum_1_io_a),
    .io_b(x558_sum_1_io_b),
    .io_flow(x558_sum_1_io_flow),
    .io_result(x558_sum_1_io_result)
  );
  RetimeWrapper_244 RetimeWrapper_11 ( // @[package.scala 93:22:@45642.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_12 ( // @[package.scala 93:22:@45651.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_242 RetimeWrapper_13 ( // @[package.scala 93:22:@45664.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  x539_sum x563_rdcol_1 ( // @[Math.scala 150:24:@45687.4]
    .clock(x563_rdcol_1_clock),
    .reset(x563_rdcol_1_reset),
    .io_a(x563_rdcol_1_io_a),
    .io_b(x563_rdcol_1_io_b),
    .io_flow(x563_rdcol_1_io_flow),
    .io_result(x563_rdcol_1_io_result)
  );
  x539_sum x567_sum_1 ( // @[Math.scala 150:24:@45708.4]
    .clock(x567_sum_1_clock),
    .reset(x567_sum_1_reset),
    .io_a(x567_sum_1_io_a),
    .io_b(x567_sum_1_io_b),
    .io_flow(x567_sum_1_io_flow),
    .io_result(x567_sum_1_io_result)
  );
  RetimeWrapper_252 RetimeWrapper_14 ( // @[package.scala 93:22:@45718.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_244 RetimeWrapper_15 ( // @[package.scala 93:22:@45727.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_242 RetimeWrapper_16 ( // @[package.scala 93:22:@45740.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  x539_sum x572_rdrow_1 ( // @[Math.scala 150:24:@45763.4]
    .clock(x572_rdrow_1_clock),
    .reset(x572_rdrow_1_reset),
    .io_a(x572_rdrow_1_io_a),
    .io_b(x572_rdrow_1_io_b),
    .io_flow(x572_rdrow_1_io_flow),
    .io_result(x572_rdrow_1_io_result)
  );
  RetimeWrapper_241 RetimeWrapper_17 ( // @[package.scala 93:22:@45844.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  x539_sum x581_sum_1 ( // @[Math.scala 150:24:@45853.4]
    .clock(x581_sum_1_clock),
    .reset(x581_sum_1_reset),
    .io_a(x581_sum_1_io_a),
    .io_b(x581_sum_1_io_b),
    .io_flow(x581_sum_1_io_flow),
    .io_result(x581_sum_1_io_result)
  );
  RetimeWrapper_244 RetimeWrapper_18 ( // @[package.scala 93:22:@45863.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_19 ( // @[package.scala 93:22:@45872.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_20 ( // @[package.scala 93:22:@45881.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_242 RetimeWrapper_21 ( // @[package.scala 93:22:@45894.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  x539_sum x587_sum_1 ( // @[Math.scala 150:24:@45917.4]
    .clock(x587_sum_1_clock),
    .reset(x587_sum_1_reset),
    .io_a(x587_sum_1_io_a),
    .io_b(x587_sum_1_io_b),
    .io_flow(x587_sum_1_io_flow),
    .io_result(x587_sum_1_io_result)
  );
  RetimeWrapper_252 RetimeWrapper_22 ( // @[package.scala 93:22:@45927.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_244 RetimeWrapper_23 ( // @[package.scala 93:22:@45936.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_242 RetimeWrapper_24 ( // @[package.scala 93:22:@45949.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  x539_sum x592_sum_1 ( // @[Math.scala 150:24:@45972.4]
    .clock(x592_sum_1_clock),
    .reset(x592_sum_1_reset),
    .io_a(x592_sum_1_io_a),
    .io_b(x592_sum_1_io_b),
    .io_flow(x592_sum_1_io_flow),
    .io_result(x592_sum_1_io_result)
  );
  RetimeWrapper_244 RetimeWrapper_25 ( // @[package.scala 93:22:@45982.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_26 ( // @[package.scala 93:22:@45991.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_242 RetimeWrapper_27 ( // @[package.scala 93:22:@46004.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x539_sum x597_sum_1 ( // @[Math.scala 150:24:@46027.4]
    .clock(x597_sum_1_clock),
    .reset(x597_sum_1_reset),
    .io_a(x597_sum_1_io_a),
    .io_b(x597_sum_1_io_b),
    .io_flow(x597_sum_1_io_flow),
    .io_result(x597_sum_1_io_result)
  );
  RetimeWrapper_252 RetimeWrapper_28 ( // @[package.scala 93:22:@46037.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_244 RetimeWrapper_29 ( // @[package.scala 93:22:@46046.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_242 RetimeWrapper_30 ( // @[package.scala 93:22:@46059.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_283 RetimeWrapper_31 ( // @[package.scala 93:22:@46080.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_283 RetimeWrapper_32 ( // @[package.scala 93:22:@46107.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_283 RetimeWrapper_33 ( // @[package.scala 93:22:@46149.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  x539_sum x609_sum_1 ( // @[Math.scala 150:24:@46158.4]
    .clock(x609_sum_1_clock),
    .reset(x609_sum_1_reset),
    .io_a(x609_sum_1_io_a),
    .io_b(x609_sum_1_io_b),
    .io_flow(x609_sum_1_io_flow),
    .io_result(x609_sum_1_io_result)
  );
  RetimeWrapper_287 RetimeWrapper_34 ( // @[package.scala 93:22:@46168.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper RetimeWrapper_35 ( // @[package.scala 93:22:@46177.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_36 ( // @[package.scala 93:22:@46186.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_241 RetimeWrapper_37 ( // @[package.scala 93:22:@46195.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_38 ( // @[package.scala 93:22:@46209.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_283 RetimeWrapper_39 ( // @[package.scala 93:22:@46230.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_283 RetimeWrapper_40 ( // @[package.scala 93:22:@46252.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  x539_sum x618_sum_1 ( // @[Math.scala 150:24:@46261.4]
    .clock(x618_sum_1_clock),
    .reset(x618_sum_1_reset),
    .io_a(x618_sum_1_io_a),
    .io_b(x618_sum_1_io_b),
    .io_flow(x618_sum_1_io_flow),
    .io_result(x618_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_41 ( // @[package.scala 93:22:@46271.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_42 ( // @[package.scala 93:22:@46285.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_283 RetimeWrapper_43 ( // @[package.scala 93:22:@46306.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_283 RetimeWrapper_44 ( // @[package.scala 93:22:@46330.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  x539_sum x626_sum_1 ( // @[Math.scala 150:24:@46339.4]
    .clock(x626_sum_1_clock),
    .reset(x626_sum_1_reset),
    .io_a(x626_sum_1_io_a),
    .io_b(x626_sum_1_io_b),
    .io_flow(x626_sum_1_io_flow),
    .io_result(x626_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_45 ( // @[package.scala 93:22:@46349.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_46 ( // @[package.scala 93:22:@46363.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_283 RetimeWrapper_47 ( // @[package.scala 93:22:@46384.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper RetimeWrapper_48 ( // @[package.scala 93:22:@46400.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_304 RetimeWrapper_49 ( // @[package.scala 93:22:@46415.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  x539_sum x634_sum_1 ( // @[Math.scala 150:24:@46424.4]
    .clock(x634_sum_1_clock),
    .reset(x634_sum_1_reset),
    .io_a(x634_sum_1_io_a),
    .io_b(x634_sum_1_io_b),
    .io_flow(x634_sum_1_io_flow),
    .io_result(x634_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_50 ( // @[package.scala 93:22:@46434.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_51 ( // @[package.scala 93:22:@46448.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  x539_sum x639_rdcol_1 ( // @[Math.scala 150:24:@46471.4]
    .clock(x639_rdcol_1_clock),
    .reset(x639_rdcol_1_reset),
    .io_a(x639_rdcol_1_io_a),
    .io_b(x639_rdcol_1_io_b),
    .io_flow(x639_rdcol_1_io_flow),
    .io_result(x639_rdcol_1_io_result)
  );
  x539_sum x645_sum_1 ( // @[Math.scala 150:24:@46503.4]
    .clock(x645_sum_1_clock),
    .reset(x645_sum_1_reset),
    .io_a(x645_sum_1_io_a),
    .io_b(x645_sum_1_io_b),
    .io_flow(x645_sum_1_io_flow),
    .io_result(x645_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_52 ( // @[package.scala 93:22:@46513.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_53 ( // @[package.scala 93:22:@46527.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  x539_sum x651_rdcol_1 ( // @[Math.scala 150:24:@46550.4]
    .clock(x651_rdcol_1_clock),
    .reset(x651_rdcol_1_reset),
    .io_a(x651_rdcol_1_io_a),
    .io_b(x651_rdcol_1_io_b),
    .io_flow(x651_rdcol_1_io_flow),
    .io_result(x651_rdcol_1_io_result)
  );
  x539_sum x657_sum_1 ( // @[Math.scala 150:24:@46582.4]
    .clock(x657_sum_1_clock),
    .reset(x657_sum_1_reset),
    .io_a(x657_sum_1_io_a),
    .io_b(x657_sum_1_io_b),
    .io_flow(x657_sum_1_io_flow),
    .io_result(x657_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_54 ( // @[package.scala 93:22:@46592.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_55 ( // @[package.scala 93:22:@46606.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_283 RetimeWrapper_56 ( // @[package.scala 93:22:@46627.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper RetimeWrapper_57 ( // @[package.scala 93:22:@46654.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_241 RetimeWrapper_58 ( // @[package.scala 93:22:@46689.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  x539_sum x669_sum_1 ( // @[Math.scala 150:24:@46700.4]
    .clock(x669_sum_1_clock),
    .reset(x669_sum_1_reset),
    .io_a(x669_sum_1_io_a),
    .io_b(x669_sum_1_io_b),
    .io_flow(x669_sum_1_io_flow),
    .io_result(x669_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_59 ( // @[package.scala 93:22:@46710.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_60 ( // @[package.scala 93:22:@46719.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_61 ( // @[package.scala 93:22:@46733.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x539_sum x677_sum_1 ( // @[Math.scala 150:24:@46760.4]
    .clock(x677_sum_1_clock),
    .reset(x677_sum_1_reset),
    .io_a(x677_sum_1_io_a),
    .io_b(x677_sum_1_io_b),
    .io_flow(x677_sum_1_io_flow),
    .io_result(x677_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_62 ( // @[package.scala 93:22:@46770.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_63 ( // @[package.scala 93:22:@46784.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  x539_sum x684_sum_1 ( // @[Math.scala 150:24:@46811.4]
    .clock(x684_sum_1_clock),
    .reset(x684_sum_1_reset),
    .io_a(x684_sum_1_io_a),
    .io_b(x684_sum_1_io_b),
    .io_flow(x684_sum_1_io_flow),
    .io_result(x684_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_64 ( // @[package.scala 93:22:@46821.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_65 ( // @[package.scala 93:22:@46835.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_283 RetimeWrapper_66 ( // @[package.scala 93:22:@46862.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  x539_sum x691_sum_1 ( // @[Math.scala 150:24:@46871.4]
    .clock(x691_sum_1_clock),
    .reset(x691_sum_1_reset),
    .io_a(x691_sum_1_io_a),
    .io_b(x691_sum_1_io_b),
    .io_flow(x691_sum_1_io_flow),
    .io_result(x691_sum_1_io_result)
  );
  RetimeWrapper_52 RetimeWrapper_67 ( // @[package.scala 93:22:@46881.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_241 RetimeWrapper_68 ( // @[package.scala 93:22:@46890.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_69 ( // @[package.scala 93:22:@46904.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  x539_sum x698_sum_1 ( // @[Math.scala 150:24:@46931.4]
    .clock(x698_sum_1_clock),
    .reset(x698_sum_1_reset),
    .io_a(x698_sum_1_io_a),
    .io_b(x698_sum_1_io_b),
    .io_flow(x698_sum_1_io_flow),
    .io_result(x698_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_70 ( // @[package.scala 93:22:@46941.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_71 ( // @[package.scala 93:22:@46955.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  x539_sum x705_sum_1 ( // @[Math.scala 150:24:@46982.4]
    .clock(x705_sum_1_clock),
    .reset(x705_sum_1_reset),
    .io_a(x705_sum_1_io_a),
    .io_b(x705_sum_1_io_b),
    .io_flow(x705_sum_1_io_flow),
    .io_result(x705_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_72 ( // @[package.scala 93:22:@46992.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_73 ( // @[package.scala 93:22:@47006.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  x539_sum x710_rdrow_1 ( // @[Math.scala 150:24:@47029.4]
    .clock(x710_rdrow_1_clock),
    .reset(x710_rdrow_1_reset),
    .io_a(x710_rdrow_1_io_a),
    .io_b(x710_rdrow_1_io_b),
    .io_flow(x710_rdrow_1_io_flow),
    .io_result(x710_rdrow_1_io_result)
  );
  x539_sum x717_sum_1 ( // @[Math.scala 150:24:@47083.4]
    .clock(x717_sum_1_clock),
    .reset(x717_sum_1_reset),
    .io_a(x717_sum_1_io_a),
    .io_b(x717_sum_1_io_b),
    .io_flow(x717_sum_1_io_flow),
    .io_result(x717_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_74 ( // @[package.scala 93:22:@47093.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_241 RetimeWrapper_75 ( // @[package.scala 93:22:@47102.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_76 ( // @[package.scala 93:22:@47116.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  x539_sum x725_sum_1 ( // @[Math.scala 150:24:@47145.4]
    .clock(x725_sum_1_clock),
    .reset(x725_sum_1_reset),
    .io_a(x725_sum_1_io_a),
    .io_b(x725_sum_1_io_b),
    .io_flow(x725_sum_1_io_flow),
    .io_result(x725_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_77 ( // @[package.scala 93:22:@47155.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_78 ( // @[package.scala 93:22:@47169.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  x539_sum x732_sum_1 ( // @[Math.scala 150:24:@47196.4]
    .clock(x732_sum_1_clock),
    .reset(x732_sum_1_reset),
    .io_a(x732_sum_1_io_a),
    .io_b(x732_sum_1_io_b),
    .io_flow(x732_sum_1_io_flow),
    .io_result(x732_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_79 ( // @[package.scala 93:22:@47206.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_80 ( // @[package.scala 93:22:@47220.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  x539_sum x739_sum_1 ( // @[Math.scala 150:24:@47247.4]
    .clock(x739_sum_1_clock),
    .reset(x739_sum_1_reset),
    .io_a(x739_sum_1_io_a),
    .io_b(x739_sum_1_io_b),
    .io_flow(x739_sum_1_io_flow),
    .io_result(x739_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_81 ( // @[package.scala 93:22:@47257.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_82 ( // @[package.scala 93:22:@47271.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  x539_sum x746_sum_1 ( // @[Math.scala 150:24:@47298.4]
    .clock(x746_sum_1_clock),
    .reset(x746_sum_1_reset),
    .io_a(x746_sum_1_io_a),
    .io_b(x746_sum_1_io_b),
    .io_flow(x746_sum_1_io_flow),
    .io_result(x746_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_83 ( // @[package.scala 93:22:@47308.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_84 ( // @[package.scala 93:22:@47322.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  x539_sum x753_sum_1 ( // @[Math.scala 150:24:@47349.4]
    .clock(x753_sum_1_clock),
    .reset(x753_sum_1_reset),
    .io_a(x753_sum_1_io_a),
    .io_b(x753_sum_1_io_b),
    .io_flow(x753_sum_1_io_flow),
    .io_result(x753_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_85 ( // @[package.scala 93:22:@47359.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_86 ( // @[package.scala 93:22:@47373.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  x539_sum x758_rdrow_1 ( // @[Math.scala 150:24:@47396.4]
    .clock(x758_rdrow_1_clock),
    .reset(x758_rdrow_1_reset),
    .io_a(x758_rdrow_1_io_a),
    .io_b(x758_rdrow_1_io_b),
    .io_flow(x758_rdrow_1_io_flow),
    .io_result(x758_rdrow_1_io_result)
  );
  x539_sum x765_sum_1 ( // @[Math.scala 150:24:@47450.4]
    .clock(x765_sum_1_clock),
    .reset(x765_sum_1_reset),
    .io_a(x765_sum_1_io_a),
    .io_b(x765_sum_1_io_b),
    .io_flow(x765_sum_1_io_flow),
    .io_result(x765_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_87 ( // @[package.scala 93:22:@47460.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_241 RetimeWrapper_88 ( // @[package.scala 93:22:@47469.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_89 ( // @[package.scala 93:22:@47483.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  x539_sum x773_sum_1 ( // @[Math.scala 150:24:@47510.4]
    .clock(x773_sum_1_clock),
    .reset(x773_sum_1_reset),
    .io_a(x773_sum_1_io_a),
    .io_b(x773_sum_1_io_b),
    .io_flow(x773_sum_1_io_flow),
    .io_result(x773_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_90 ( // @[package.scala 93:22:@47520.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_91 ( // @[package.scala 93:22:@47534.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  x539_sum x780_sum_1 ( // @[Math.scala 150:24:@47563.4]
    .clock(x780_sum_1_clock),
    .reset(x780_sum_1_reset),
    .io_a(x780_sum_1_io_a),
    .io_b(x780_sum_1_io_b),
    .io_flow(x780_sum_1_io_flow),
    .io_result(x780_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_92 ( // @[package.scala 93:22:@47573.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_93 ( // @[package.scala 93:22:@47587.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  x539_sum x787_sum_1 ( // @[Math.scala 150:24:@47614.4]
    .clock(x787_sum_1_clock),
    .reset(x787_sum_1_reset),
    .io_a(x787_sum_1_io_a),
    .io_b(x787_sum_1_io_b),
    .io_flow(x787_sum_1_io_flow),
    .io_result(x787_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_94 ( // @[package.scala 93:22:@47624.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_95 ( // @[package.scala 93:22:@47638.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  x539_sum x794_sum_1 ( // @[Math.scala 150:24:@47665.4]
    .clock(x794_sum_1_clock),
    .reset(x794_sum_1_reset),
    .io_a(x794_sum_1_io_a),
    .io_b(x794_sum_1_io_b),
    .io_flow(x794_sum_1_io_flow),
    .io_result(x794_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_96 ( // @[package.scala 93:22:@47675.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_97 ( // @[package.scala 93:22:@47689.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  x539_sum x801_sum_1 ( // @[Math.scala 150:24:@47716.4]
    .clock(x801_sum_1_clock),
    .reset(x801_sum_1_reset),
    .io_a(x801_sum_1_io_a),
    .io_b(x801_sum_1_io_b),
    .io_flow(x801_sum_1_io_flow),
    .io_result(x801_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_98 ( // @[package.scala 93:22:@47726.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_287 RetimeWrapper_99 ( // @[package.scala 93:22:@47740.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  x811_x23 x811_x23_1 ( // @[Math.scala 150:24:@47786.4]
    .clock(x811_x23_1_clock),
    .reset(x811_x23_1_reset),
    .io_a(x811_x23_1_io_a),
    .io_b(x811_x23_1_io_b),
    .io_flow(x811_x23_1_io_flow),
    .io_result(x811_x23_1_io_result)
  );
  x811_x23 x812_x24_1 ( // @[Math.scala 150:24:@47796.4]
    .clock(x812_x24_1_clock),
    .reset(x812_x24_1_reset),
    .io_a(x812_x24_1_io_a),
    .io_b(x812_x24_1_io_b),
    .io_flow(x812_x24_1_io_flow),
    .io_result(x812_x24_1_io_result)
  );
  x811_x23 x813_x23_1 ( // @[Math.scala 150:24:@47806.4]
    .clock(x813_x23_1_clock),
    .reset(x813_x23_1_reset),
    .io_a(x813_x23_1_io_a),
    .io_b(x813_x23_1_io_b),
    .io_flow(x813_x23_1_io_flow),
    .io_result(x813_x23_1_io_result)
  );
  x811_x23 x814_x24_1 ( // @[Math.scala 150:24:@47816.4]
    .clock(x814_x24_1_clock),
    .reset(x814_x24_1_reset),
    .io_a(x814_x24_1_io_a),
    .io_b(x814_x24_1_io_b),
    .io_flow(x814_x24_1_io_flow),
    .io_result(x814_x24_1_io_result)
  );
  x815_x23 x815_x23_1 ( // @[Math.scala 150:24:@47826.4]
    .io_a(x815_x23_1_io_a),
    .io_b(x815_x23_1_io_b),
    .io_result(x815_x23_1_io_result)
  );
  x815_x23 x816_x24_1 ( // @[Math.scala 150:24:@47836.4]
    .io_a(x816_x24_1_io_a),
    .io_b(x816_x24_1_io_b),
    .io_result(x816_x24_1_io_result)
  );
  x815_x23 x817_x23_1 ( // @[Math.scala 150:24:@47846.4]
    .io_a(x817_x23_1_io_a),
    .io_b(x817_x23_1_io_b),
    .io_result(x817_x23_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_100 ( // @[package.scala 93:22:@47856.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  x815_x23 x818_sum_1 ( // @[Math.scala 150:24:@47865.4]
    .io_a(x818_sum_1_io_a),
    .io_b(x818_sum_1_io_b),
    .io_result(x818_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_101 ( // @[package.scala 93:22:@47879.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  x811_x23 x825_x23_1 ( // @[Math.scala 150:24:@47914.4]
    .clock(x825_x23_1_clock),
    .reset(x825_x23_1_reset),
    .io_a(x825_x23_1_io_a),
    .io_b(x825_x23_1_io_b),
    .io_flow(x825_x23_1_io_flow),
    .io_result(x825_x23_1_io_result)
  );
  x811_x23 x826_x24_1 ( // @[Math.scala 150:24:@47924.4]
    .clock(x826_x24_1_clock),
    .reset(x826_x24_1_reset),
    .io_a(x826_x24_1_io_a),
    .io_b(x826_x24_1_io_b),
    .io_flow(x826_x24_1_io_flow),
    .io_result(x826_x24_1_io_result)
  );
  x811_x23 x827_x23_1 ( // @[Math.scala 150:24:@47934.4]
    .clock(x827_x23_1_clock),
    .reset(x827_x23_1_reset),
    .io_a(x827_x23_1_io_a),
    .io_b(x827_x23_1_io_b),
    .io_flow(x827_x23_1_io_flow),
    .io_result(x827_x23_1_io_result)
  );
  x811_x23 x828_x24_1 ( // @[Math.scala 150:24:@47944.4]
    .clock(x828_x24_1_clock),
    .reset(x828_x24_1_reset),
    .io_a(x828_x24_1_io_a),
    .io_b(x828_x24_1_io_b),
    .io_flow(x828_x24_1_io_flow),
    .io_result(x828_x24_1_io_result)
  );
  x815_x23 x829_x23_1 ( // @[Math.scala 150:24:@47954.4]
    .io_a(x829_x23_1_io_a),
    .io_b(x829_x23_1_io_b),
    .io_result(x829_x23_1_io_result)
  );
  x815_x23 x830_x24_1 ( // @[Math.scala 150:24:@47964.4]
    .io_a(x830_x24_1_io_a),
    .io_b(x830_x24_1_io_b),
    .io_result(x830_x24_1_io_result)
  );
  x815_x23 x831_x23_1 ( // @[Math.scala 150:24:@47976.4]
    .io_a(x831_x23_1_io_a),
    .io_b(x831_x23_1_io_b),
    .io_result(x831_x23_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_102 ( // @[package.scala 93:22:@47986.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  x815_x23 x832_sum_1 ( // @[Math.scala 150:24:@47995.4]
    .io_a(x832_sum_1_io_a),
    .io_b(x832_sum_1_io_b),
    .io_result(x832_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_103 ( // @[package.scala 93:22:@48009.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  x811_x23 x838_x23_1 ( // @[Math.scala 150:24:@48039.4]
    .clock(x838_x23_1_clock),
    .reset(x838_x23_1_reset),
    .io_a(x838_x23_1_io_a),
    .io_b(x838_x23_1_io_b),
    .io_flow(x838_x23_1_io_flow),
    .io_result(x838_x23_1_io_result)
  );
  x811_x23 x839_x24_1 ( // @[Math.scala 150:24:@48049.4]
    .clock(x839_x24_1_clock),
    .reset(x839_x24_1_reset),
    .io_a(x839_x24_1_io_a),
    .io_b(x839_x24_1_io_b),
    .io_flow(x839_x24_1_io_flow),
    .io_result(x839_x24_1_io_result)
  );
  x811_x23 x840_x23_1 ( // @[Math.scala 150:24:@48059.4]
    .clock(x840_x23_1_clock),
    .reset(x840_x23_1_reset),
    .io_a(x840_x23_1_io_a),
    .io_b(x840_x23_1_io_b),
    .io_flow(x840_x23_1_io_flow),
    .io_result(x840_x23_1_io_result)
  );
  x811_x23 x841_x24_1 ( // @[Math.scala 150:24:@48069.4]
    .clock(x841_x24_1_clock),
    .reset(x841_x24_1_reset),
    .io_a(x841_x24_1_io_a),
    .io_b(x841_x24_1_io_b),
    .io_flow(x841_x24_1_io_flow),
    .io_result(x841_x24_1_io_result)
  );
  x815_x23 x842_x23_1 ( // @[Math.scala 150:24:@48079.4]
    .io_a(x842_x23_1_io_a),
    .io_b(x842_x23_1_io_b),
    .io_result(x842_x23_1_io_result)
  );
  x815_x23 x843_x24_1 ( // @[Math.scala 150:24:@48089.4]
    .io_a(x843_x24_1_io_a),
    .io_b(x843_x24_1_io_b),
    .io_result(x843_x24_1_io_result)
  );
  x815_x23 x844_x23_1 ( // @[Math.scala 150:24:@48099.4]
    .io_a(x844_x23_1_io_a),
    .io_b(x844_x23_1_io_b),
    .io_result(x844_x23_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_104 ( // @[package.scala 93:22:@48109.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  x815_x23 x845_sum_1 ( // @[Math.scala 150:24:@48118.4]
    .io_a(x845_sum_1_io_a),
    .io_b(x845_sum_1_io_b),
    .io_result(x845_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_105 ( // @[package.scala 93:22:@48132.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  x811_x23 x851_x23_1 ( // @[Math.scala 150:24:@48162.4]
    .clock(x851_x23_1_clock),
    .reset(x851_x23_1_reset),
    .io_a(x851_x23_1_io_a),
    .io_b(x851_x23_1_io_b),
    .io_flow(x851_x23_1_io_flow),
    .io_result(x851_x23_1_io_result)
  );
  x811_x23 x852_x24_1 ( // @[Math.scala 150:24:@48172.4]
    .clock(x852_x24_1_clock),
    .reset(x852_x24_1_reset),
    .io_a(x852_x24_1_io_a),
    .io_b(x852_x24_1_io_b),
    .io_flow(x852_x24_1_io_flow),
    .io_result(x852_x24_1_io_result)
  );
  x811_x23 x853_x23_1 ( // @[Math.scala 150:24:@48182.4]
    .clock(x853_x23_1_clock),
    .reset(x853_x23_1_reset),
    .io_a(x853_x23_1_io_a),
    .io_b(x853_x23_1_io_b),
    .io_flow(x853_x23_1_io_flow),
    .io_result(x853_x23_1_io_result)
  );
  x811_x23 x854_x24_1 ( // @[Math.scala 150:24:@48192.4]
    .clock(x854_x24_1_clock),
    .reset(x854_x24_1_reset),
    .io_a(x854_x24_1_io_a),
    .io_b(x854_x24_1_io_b),
    .io_flow(x854_x24_1_io_flow),
    .io_result(x854_x24_1_io_result)
  );
  x815_x23 x855_x23_1 ( // @[Math.scala 150:24:@48202.4]
    .io_a(x855_x23_1_io_a),
    .io_b(x855_x23_1_io_b),
    .io_result(x855_x23_1_io_result)
  );
  x815_x23 x856_x24_1 ( // @[Math.scala 150:24:@48212.4]
    .io_a(x856_x24_1_io_a),
    .io_b(x856_x24_1_io_b),
    .io_result(x856_x24_1_io_result)
  );
  x815_x23 x857_x23_1 ( // @[Math.scala 150:24:@48222.4]
    .io_a(x857_x23_1_io_a),
    .io_b(x857_x23_1_io_b),
    .io_result(x857_x23_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_106 ( // @[package.scala 93:22:@48232.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  x815_x23 x858_sum_1 ( // @[Math.scala 150:24:@48241.4]
    .io_a(x858_sum_1_io_a),
    .io_b(x858_sum_1_io_b),
    .io_result(x858_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_107 ( // @[package.scala 93:22:@48255.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  x811_x23 x863_x23_1 ( // @[Math.scala 150:24:@48280.4]
    .clock(x863_x23_1_clock),
    .reset(x863_x23_1_reset),
    .io_a(x863_x23_1_io_a),
    .io_b(x863_x23_1_io_b),
    .io_flow(x863_x23_1_io_flow),
    .io_result(x863_x23_1_io_result)
  );
  x811_x23 x864_x24_1 ( // @[Math.scala 150:24:@48290.4]
    .clock(x864_x24_1_clock),
    .reset(x864_x24_1_reset),
    .io_a(x864_x24_1_io_a),
    .io_b(x864_x24_1_io_b),
    .io_flow(x864_x24_1_io_flow),
    .io_result(x864_x24_1_io_result)
  );
  x811_x23 x865_x23_1 ( // @[Math.scala 150:24:@48300.4]
    .clock(x865_x23_1_clock),
    .reset(x865_x23_1_reset),
    .io_a(x865_x23_1_io_a),
    .io_b(x865_x23_1_io_b),
    .io_flow(x865_x23_1_io_flow),
    .io_result(x865_x23_1_io_result)
  );
  x811_x23 x866_x24_1 ( // @[Math.scala 150:24:@48310.4]
    .clock(x866_x24_1_clock),
    .reset(x866_x24_1_reset),
    .io_a(x866_x24_1_io_a),
    .io_b(x866_x24_1_io_b),
    .io_flow(x866_x24_1_io_flow),
    .io_result(x866_x24_1_io_result)
  );
  x815_x23 x867_x23_1 ( // @[Math.scala 150:24:@48320.4]
    .io_a(x867_x23_1_io_a),
    .io_b(x867_x23_1_io_b),
    .io_result(x867_x23_1_io_result)
  );
  x815_x23 x868_x24_1 ( // @[Math.scala 150:24:@48330.4]
    .io_a(x868_x24_1_io_a),
    .io_b(x868_x24_1_io_b),
    .io_result(x868_x24_1_io_result)
  );
  x815_x23 x869_x23_1 ( // @[Math.scala 150:24:@48340.4]
    .io_a(x869_x23_1_io_a),
    .io_b(x869_x23_1_io_b),
    .io_result(x869_x23_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_108 ( // @[package.scala 93:22:@48350.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  x815_x23 x870_sum_1 ( // @[Math.scala 150:24:@48359.4]
    .io_a(x870_sum_1_io_a),
    .io_b(x870_sum_1_io_b),
    .io_result(x870_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_109 ( // @[package.scala 93:22:@48373.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  x811_x23 x874_x23_1 ( // @[Math.scala 150:24:@48393.4]
    .clock(x874_x23_1_clock),
    .reset(x874_x23_1_reset),
    .io_a(x874_x23_1_io_a),
    .io_b(x874_x23_1_io_b),
    .io_flow(x874_x23_1_io_flow),
    .io_result(x874_x23_1_io_result)
  );
  x811_x23 x875_x24_1 ( // @[Math.scala 150:24:@48403.4]
    .clock(x875_x24_1_clock),
    .reset(x875_x24_1_reset),
    .io_a(x875_x24_1_io_a),
    .io_b(x875_x24_1_io_b),
    .io_flow(x875_x24_1_io_flow),
    .io_result(x875_x24_1_io_result)
  );
  x811_x23 x876_x23_1 ( // @[Math.scala 150:24:@48415.4]
    .clock(x876_x23_1_clock),
    .reset(x876_x23_1_reset),
    .io_a(x876_x23_1_io_a),
    .io_b(x876_x23_1_io_b),
    .io_flow(x876_x23_1_io_flow),
    .io_result(x876_x23_1_io_result)
  );
  x811_x23 x877_x24_1 ( // @[Math.scala 150:24:@48425.4]
    .clock(x877_x24_1_clock),
    .reset(x877_x24_1_reset),
    .io_a(x877_x24_1_io_a),
    .io_b(x877_x24_1_io_b),
    .io_flow(x877_x24_1_io_flow),
    .io_result(x877_x24_1_io_result)
  );
  x815_x23 x878_x23_1 ( // @[Math.scala 150:24:@48435.4]
    .io_a(x878_x23_1_io_a),
    .io_b(x878_x23_1_io_b),
    .io_result(x878_x23_1_io_result)
  );
  x815_x23 x879_x24_1 ( // @[Math.scala 150:24:@48445.4]
    .io_a(x879_x24_1_io_a),
    .io_b(x879_x24_1_io_b),
    .io_result(x879_x24_1_io_result)
  );
  x815_x23 x880_x23_1 ( // @[Math.scala 150:24:@48455.4]
    .io_a(x880_x23_1_io_a),
    .io_b(x880_x23_1_io_b),
    .io_result(x880_x23_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_110 ( // @[package.scala 93:22:@48465.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  x815_x23 x881_sum_1 ( // @[Math.scala 150:24:@48474.4]
    .io_a(x881_sum_1_io_a),
    .io_b(x881_sum_1_io_b),
    .io_result(x881_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_111 ( // @[package.scala 93:22:@48488.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  x811_x23 x885_x23_1 ( // @[Math.scala 150:24:@48508.4]
    .clock(x885_x23_1_clock),
    .reset(x885_x23_1_reset),
    .io_a(x885_x23_1_io_a),
    .io_b(x885_x23_1_io_b),
    .io_flow(x885_x23_1_io_flow),
    .io_result(x885_x23_1_io_result)
  );
  x811_x23 x886_x24_1 ( // @[Math.scala 150:24:@48518.4]
    .clock(x886_x24_1_clock),
    .reset(x886_x24_1_reset),
    .io_a(x886_x24_1_io_a),
    .io_b(x886_x24_1_io_b),
    .io_flow(x886_x24_1_io_flow),
    .io_result(x886_x24_1_io_result)
  );
  x811_x23 x887_x23_1 ( // @[Math.scala 150:24:@48528.4]
    .clock(x887_x23_1_clock),
    .reset(x887_x23_1_reset),
    .io_a(x887_x23_1_io_a),
    .io_b(x887_x23_1_io_b),
    .io_flow(x887_x23_1_io_flow),
    .io_result(x887_x23_1_io_result)
  );
  x811_x23 x888_x24_1 ( // @[Math.scala 150:24:@48538.4]
    .clock(x888_x24_1_clock),
    .reset(x888_x24_1_reset),
    .io_a(x888_x24_1_io_a),
    .io_b(x888_x24_1_io_b),
    .io_flow(x888_x24_1_io_flow),
    .io_result(x888_x24_1_io_result)
  );
  x815_x23 x889_x23_1 ( // @[Math.scala 150:24:@48548.4]
    .io_a(x889_x23_1_io_a),
    .io_b(x889_x23_1_io_b),
    .io_result(x889_x23_1_io_result)
  );
  x815_x23 x890_x24_1 ( // @[Math.scala 150:24:@48558.4]
    .io_a(x890_x24_1_io_a),
    .io_b(x890_x24_1_io_b),
    .io_result(x890_x24_1_io_result)
  );
  x815_x23 x891_x23_1 ( // @[Math.scala 150:24:@48568.4]
    .io_a(x891_x23_1_io_a),
    .io_b(x891_x23_1_io_b),
    .io_result(x891_x23_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_112 ( // @[package.scala 93:22:@48578.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  x815_x23 x892_sum_1 ( // @[Math.scala 150:24:@48587.4]
    .io_a(x892_sum_1_io_a),
    .io_b(x892_sum_1_io_b),
    .io_result(x892_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_113 ( // @[package.scala 93:22:@48601.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  x811_x23 x897_x23_1 ( // @[Math.scala 150:24:@48626.4]
    .clock(x897_x23_1_clock),
    .reset(x897_x23_1_reset),
    .io_a(x897_x23_1_io_a),
    .io_b(x897_x23_1_io_b),
    .io_flow(x897_x23_1_io_flow),
    .io_result(x897_x23_1_io_result)
  );
  x811_x23 x898_x24_1 ( // @[Math.scala 150:24:@48636.4]
    .clock(x898_x24_1_clock),
    .reset(x898_x24_1_reset),
    .io_a(x898_x24_1_io_a),
    .io_b(x898_x24_1_io_b),
    .io_flow(x898_x24_1_io_flow),
    .io_result(x898_x24_1_io_result)
  );
  x811_x23 x899_x23_1 ( // @[Math.scala 150:24:@48646.4]
    .clock(x899_x23_1_clock),
    .reset(x899_x23_1_reset),
    .io_a(x899_x23_1_io_a),
    .io_b(x899_x23_1_io_b),
    .io_flow(x899_x23_1_io_flow),
    .io_result(x899_x23_1_io_result)
  );
  x811_x23 x900_x24_1 ( // @[Math.scala 150:24:@48656.4]
    .clock(x900_x24_1_clock),
    .reset(x900_x24_1_reset),
    .io_a(x900_x24_1_io_a),
    .io_b(x900_x24_1_io_b),
    .io_flow(x900_x24_1_io_flow),
    .io_result(x900_x24_1_io_result)
  );
  x815_x23 x901_x23_1 ( // @[Math.scala 150:24:@48666.4]
    .io_a(x901_x23_1_io_a),
    .io_b(x901_x23_1_io_b),
    .io_result(x901_x23_1_io_result)
  );
  x815_x23 x902_x24_1 ( // @[Math.scala 150:24:@48676.4]
    .io_a(x902_x24_1_io_a),
    .io_b(x902_x24_1_io_b),
    .io_result(x902_x24_1_io_result)
  );
  x815_x23 x903_x23_1 ( // @[Math.scala 150:24:@48686.4]
    .io_a(x903_x23_1_io_a),
    .io_b(x903_x23_1_io_b),
    .io_result(x903_x23_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_114 ( // @[package.scala 93:22:@48696.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  x815_x23 x904_sum_1 ( // @[Math.scala 150:24:@48705.4]
    .io_a(x904_sum_1_io_a),
    .io_b(x904_sum_1_io_b),
    .io_result(x904_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_115 ( // @[package.scala 93:22:@48719.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_428 RetimeWrapper_116 ( // @[package.scala 93:22:@48729.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  RetimeWrapper_429 RetimeWrapper_117 ( // @[package.scala 93:22:@48738.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_118 ( // @[package.scala 93:22:@48747.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  RetimeWrapper_428 RetimeWrapper_119 ( // @[package.scala 93:22:@48756.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  RetimeWrapper_432 RetimeWrapper_120 ( // @[package.scala 93:22:@48765.4]
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  RetimeWrapper_428 RetimeWrapper_121 ( // @[package.scala 93:22:@48778.4]
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_122 ( // @[package.scala 93:22:@48799.4]
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  RetimeWrapper_435 RetimeWrapper_123 ( // @[package.scala 93:22:@48808.4]
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  RetimeWrapper_428 RetimeWrapper_124 ( // @[package.scala 93:22:@48821.4]
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  RetimeWrapper_435 RetimeWrapper_125 ( // @[package.scala 93:22:@48842.4]
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_126 ( // @[package.scala 93:22:@48851.4]
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  RetimeWrapper_428 RetimeWrapper_127 ( // @[package.scala 93:22:@48864.4]
    .clock(RetimeWrapper_127_clock),
    .reset(RetimeWrapper_127_reset),
    .io_flow(RetimeWrapper_127_io_flow),
    .io_in(RetimeWrapper_127_io_in),
    .io_out(RetimeWrapper_127_io_out)
  );
  RetimeWrapper_435 RetimeWrapper_128 ( // @[package.scala 93:22:@48885.4]
    .clock(RetimeWrapper_128_clock),
    .reset(RetimeWrapper_128_reset),
    .io_flow(RetimeWrapper_128_io_flow),
    .io_in(RetimeWrapper_128_io_in),
    .io_out(RetimeWrapper_128_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_129 ( // @[package.scala 93:22:@48894.4]
    .clock(RetimeWrapper_129_clock),
    .reset(RetimeWrapper_129_reset),
    .io_flow(RetimeWrapper_129_io_flow),
    .io_in(RetimeWrapper_129_io_in),
    .io_out(RetimeWrapper_129_io_out)
  );
  RetimeWrapper_428 RetimeWrapper_130 ( // @[package.scala 93:22:@48907.4]
    .clock(RetimeWrapper_130_clock),
    .reset(RetimeWrapper_130_reset),
    .io_flow(RetimeWrapper_130_io_flow),
    .io_in(RetimeWrapper_130_io_in),
    .io_out(RetimeWrapper_130_io_out)
  );
  RetimeWrapper_432 RetimeWrapper_131 ( // @[package.scala 93:22:@48928.4]
    .clock(RetimeWrapper_131_clock),
    .reset(RetimeWrapper_131_reset),
    .io_flow(RetimeWrapper_131_io_flow),
    .io_in(RetimeWrapper_131_io_in),
    .io_out(RetimeWrapper_131_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_132 ( // @[package.scala 93:22:@48937.4]
    .clock(RetimeWrapper_132_clock),
    .reset(RetimeWrapper_132_reset),
    .io_flow(RetimeWrapper_132_io_flow),
    .io_in(RetimeWrapper_132_io_in),
    .io_out(RetimeWrapper_132_io_out)
  );
  RetimeWrapper_435 RetimeWrapper_133 ( // @[package.scala 93:22:@48946.4]
    .clock(RetimeWrapper_133_clock),
    .reset(RetimeWrapper_133_reset),
    .io_flow(RetimeWrapper_133_io_flow),
    .io_in(RetimeWrapper_133_io_in),
    .io_out(RetimeWrapper_133_io_out)
  );
  RetimeWrapper_428 RetimeWrapper_134 ( // @[package.scala 93:22:@48959.4]
    .clock(RetimeWrapper_134_clock),
    .reset(RetimeWrapper_134_reset),
    .io_flow(RetimeWrapper_134_io_flow),
    .io_in(RetimeWrapper_134_io_in),
    .io_out(RetimeWrapper_134_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_135 ( // @[package.scala 93:22:@48980.4]
    .clock(RetimeWrapper_135_clock),
    .reset(RetimeWrapper_135_reset),
    .io_flow(RetimeWrapper_135_io_flow),
    .io_in(RetimeWrapper_135_io_in),
    .io_out(RetimeWrapper_135_io_out)
  );
  RetimeWrapper_435 RetimeWrapper_136 ( // @[package.scala 93:22:@48989.4]
    .clock(RetimeWrapper_136_clock),
    .reset(RetimeWrapper_136_reset),
    .io_flow(RetimeWrapper_136_io_flow),
    .io_in(RetimeWrapper_136_io_in),
    .io_out(RetimeWrapper_136_io_out)
  );
  RetimeWrapper_428 RetimeWrapper_137 ( // @[package.scala 93:22:@49002.4]
    .clock(RetimeWrapper_137_clock),
    .reset(RetimeWrapper_137_reset),
    .io_flow(RetimeWrapper_137_io_flow),
    .io_in(RetimeWrapper_137_io_in),
    .io_out(RetimeWrapper_137_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_138 ( // @[package.scala 93:22:@49023.4]
    .clock(RetimeWrapper_138_clock),
    .reset(RetimeWrapper_138_reset),
    .io_flow(RetimeWrapper_138_io_flow),
    .io_in(RetimeWrapper_138_io_in),
    .io_out(RetimeWrapper_138_io_out)
  );
  RetimeWrapper_435 RetimeWrapper_139 ( // @[package.scala 93:22:@49032.4]
    .clock(RetimeWrapper_139_clock),
    .reset(RetimeWrapper_139_reset),
    .io_flow(RetimeWrapper_139_io_flow),
    .io_in(RetimeWrapper_139_io_in),
    .io_out(RetimeWrapper_139_io_out)
  );
  RetimeWrapper_428 RetimeWrapper_140 ( // @[package.scala 93:22:@49045.4]
    .clock(RetimeWrapper_140_clock),
    .reset(RetimeWrapper_140_reset),
    .io_flow(RetimeWrapper_140_io_flow),
    .io_in(RetimeWrapper_140_io_in),
    .io_out(RetimeWrapper_140_io_out)
  );
  RetimeWrapper_435 RetimeWrapper_141 ( // @[package.scala 93:22:@49066.4]
    .clock(RetimeWrapper_141_clock),
    .reset(RetimeWrapper_141_reset),
    .io_flow(RetimeWrapper_141_io_flow),
    .io_in(RetimeWrapper_141_io_in),
    .io_out(RetimeWrapper_141_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_142 ( // @[package.scala 93:22:@49075.4]
    .clock(RetimeWrapper_142_clock),
    .reset(RetimeWrapper_142_reset),
    .io_flow(RetimeWrapper_142_io_flow),
    .io_in(RetimeWrapper_142_io_in),
    .io_out(RetimeWrapper_142_io_out)
  );
  RetimeWrapper_428 RetimeWrapper_143 ( // @[package.scala 93:22:@49088.4]
    .clock(RetimeWrapper_143_clock),
    .reset(RetimeWrapper_143_reset),
    .io_flow(RetimeWrapper_143_io_flow),
    .io_in(RetimeWrapper_143_io_in),
    .io_out(RetimeWrapper_143_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_144 ( // @[package.scala 93:22:@49109.4]
    .clock(RetimeWrapper_144_clock),
    .reset(RetimeWrapper_144_reset),
    .io_flow(RetimeWrapper_144_io_flow),
    .io_in(RetimeWrapper_144_io_in),
    .io_out(RetimeWrapper_144_io_out)
  );
  RetimeWrapper_457 RetimeWrapper_145 ( // @[package.scala 93:22:@49118.4]
    .clock(RetimeWrapper_145_clock),
    .reset(RetimeWrapper_145_reset),
    .io_flow(RetimeWrapper_145_io_flow),
    .io_in(RetimeWrapper_145_io_in),
    .io_out(RetimeWrapper_145_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_146 ( // @[package.scala 93:22:@49127.4]
    .clock(RetimeWrapper_146_clock),
    .reset(RetimeWrapper_146_reset),
    .io_flow(RetimeWrapper_146_io_flow),
    .io_in(RetimeWrapper_146_io_in),
    .io_out(RetimeWrapper_146_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_147 ( // @[package.scala 93:22:@49136.4]
    .clock(RetimeWrapper_147_clock),
    .reset(RetimeWrapper_147_reset),
    .io_flow(RetimeWrapper_147_io_flow),
    .io_in(RetimeWrapper_147_io_in),
    .io_out(RetimeWrapper_147_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_148 ( // @[package.scala 93:22:@49145.4]
    .clock(RetimeWrapper_148_clock),
    .reset(RetimeWrapper_148_reset),
    .io_flow(RetimeWrapper_148_io_flow),
    .io_in(RetimeWrapper_148_io_in),
    .io_out(RetimeWrapper_148_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_149 ( // @[package.scala 93:22:@49159.4]
    .clock(RetimeWrapper_149_clock),
    .reset(RetimeWrapper_149_reset),
    .io_flow(RetimeWrapper_149_io_flow),
    .io_in(RetimeWrapper_149_io_in),
    .io_out(RetimeWrapper_149_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_150 ( // @[package.scala 93:22:@49180.4]
    .clock(RetimeWrapper_150_clock),
    .reset(RetimeWrapper_150_reset),
    .io_flow(RetimeWrapper_150_io_flow),
    .io_in(RetimeWrapper_150_io_in),
    .io_out(RetimeWrapper_150_io_out)
  );
  RetimeWrapper_457 RetimeWrapper_151 ( // @[package.scala 93:22:@49189.4]
    .clock(RetimeWrapper_151_clock),
    .reset(RetimeWrapper_151_reset),
    .io_flow(RetimeWrapper_151_io_flow),
    .io_in(RetimeWrapper_151_io_in),
    .io_out(RetimeWrapper_151_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_152 ( // @[package.scala 93:22:@49203.4]
    .clock(RetimeWrapper_152_clock),
    .reset(RetimeWrapper_152_reset),
    .io_flow(RetimeWrapper_152_io_flow),
    .io_in(RetimeWrapper_152_io_in),
    .io_out(RetimeWrapper_152_io_out)
  );
  RetimeWrapper_457 RetimeWrapper_153 ( // @[package.scala 93:22:@49224.4]
    .clock(RetimeWrapper_153_clock),
    .reset(RetimeWrapper_153_reset),
    .io_flow(RetimeWrapper_153_io_flow),
    .io_in(RetimeWrapper_153_io_in),
    .io_out(RetimeWrapper_153_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_154 ( // @[package.scala 93:22:@49233.4]
    .clock(RetimeWrapper_154_clock),
    .reset(RetimeWrapper_154_reset),
    .io_flow(RetimeWrapper_154_io_flow),
    .io_in(RetimeWrapper_154_io_in),
    .io_out(RetimeWrapper_154_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_155 ( // @[package.scala 93:22:@49247.4]
    .clock(RetimeWrapper_155_clock),
    .reset(RetimeWrapper_155_reset),
    .io_flow(RetimeWrapper_155_io_flow),
    .io_in(RetimeWrapper_155_io_in),
    .io_out(RetimeWrapper_155_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_156 ( // @[package.scala 93:22:@49268.4]
    .clock(RetimeWrapper_156_clock),
    .reset(RetimeWrapper_156_reset),
    .io_flow(RetimeWrapper_156_io_flow),
    .io_in(RetimeWrapper_156_io_in),
    .io_out(RetimeWrapper_156_io_out)
  );
  RetimeWrapper_457 RetimeWrapper_157 ( // @[package.scala 93:22:@49277.4]
    .clock(RetimeWrapper_157_clock),
    .reset(RetimeWrapper_157_reset),
    .io_flow(RetimeWrapper_157_io_flow),
    .io_in(RetimeWrapper_157_io_in),
    .io_out(RetimeWrapper_157_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_158 ( // @[package.scala 93:22:@49291.4]
    .clock(RetimeWrapper_158_clock),
    .reset(RetimeWrapper_158_reset),
    .io_flow(RetimeWrapper_158_io_flow),
    .io_in(RetimeWrapper_158_io_in),
    .io_out(RetimeWrapper_158_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_159 ( // @[package.scala 93:22:@49312.4]
    .clock(RetimeWrapper_159_clock),
    .reset(RetimeWrapper_159_reset),
    .io_flow(RetimeWrapper_159_io_flow),
    .io_in(RetimeWrapper_159_io_in),
    .io_out(RetimeWrapper_159_io_out)
  );
  RetimeWrapper_457 RetimeWrapper_160 ( // @[package.scala 93:22:@49321.4]
    .clock(RetimeWrapper_160_clock),
    .reset(RetimeWrapper_160_reset),
    .io_flow(RetimeWrapper_160_io_flow),
    .io_in(RetimeWrapper_160_io_in),
    .io_out(RetimeWrapper_160_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_161 ( // @[package.scala 93:22:@49335.4]
    .clock(RetimeWrapper_161_clock),
    .reset(RetimeWrapper_161_reset),
    .io_flow(RetimeWrapper_161_io_flow),
    .io_in(RetimeWrapper_161_io_in),
    .io_out(RetimeWrapper_161_io_out)
  );
  RetimeWrapper_457 RetimeWrapper_162 ( // @[package.scala 93:22:@49356.4]
    .clock(RetimeWrapper_162_clock),
    .reset(RetimeWrapper_162_reset),
    .io_flow(RetimeWrapper_162_io_flow),
    .io_in(RetimeWrapper_162_io_in),
    .io_out(RetimeWrapper_162_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_163 ( // @[package.scala 93:22:@49365.4]
    .clock(RetimeWrapper_163_clock),
    .reset(RetimeWrapper_163_reset),
    .io_flow(RetimeWrapper_163_io_flow),
    .io_in(RetimeWrapper_163_io_in),
    .io_out(RetimeWrapper_163_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_164 ( // @[package.scala 93:22:@49374.4]
    .clock(RetimeWrapper_164_clock),
    .reset(RetimeWrapper_164_reset),
    .io_flow(RetimeWrapper_164_io_flow),
    .io_in(RetimeWrapper_164_io_in),
    .io_out(RetimeWrapper_164_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_165 ( // @[package.scala 93:22:@49388.4]
    .clock(RetimeWrapper_165_clock),
    .reset(RetimeWrapper_165_reset),
    .io_flow(RetimeWrapper_165_io_flow),
    .io_in(RetimeWrapper_165_io_in),
    .io_out(RetimeWrapper_165_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_166 ( // @[package.scala 93:22:@49409.4]
    .clock(RetimeWrapper_166_clock),
    .reset(RetimeWrapper_166_reset),
    .io_flow(RetimeWrapper_166_io_flow),
    .io_in(RetimeWrapper_166_io_in),
    .io_out(RetimeWrapper_166_io_out)
  );
  RetimeWrapper_457 RetimeWrapper_167 ( // @[package.scala 93:22:@49418.4]
    .clock(RetimeWrapper_167_clock),
    .reset(RetimeWrapper_167_reset),
    .io_flow(RetimeWrapper_167_io_flow),
    .io_in(RetimeWrapper_167_io_in),
    .io_out(RetimeWrapper_167_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_168 ( // @[package.scala 93:22:@49432.4]
    .clock(RetimeWrapper_168_clock),
    .reset(RetimeWrapper_168_reset),
    .io_flow(RetimeWrapper_168_io_flow),
    .io_in(RetimeWrapper_168_io_in),
    .io_out(RetimeWrapper_168_io_out)
  );
  RetimeWrapper_457 RetimeWrapper_169 ( // @[package.scala 93:22:@49453.4]
    .clock(RetimeWrapper_169_clock),
    .reset(RetimeWrapper_169_reset),
    .io_flow(RetimeWrapper_169_io_flow),
    .io_in(RetimeWrapper_169_io_in),
    .io_out(RetimeWrapper_169_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_170 ( // @[package.scala 93:22:@49462.4]
    .clock(RetimeWrapper_170_clock),
    .reset(RetimeWrapper_170_reset),
    .io_flow(RetimeWrapper_170_io_flow),
    .io_in(RetimeWrapper_170_io_in),
    .io_out(RetimeWrapper_170_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_171 ( // @[package.scala 93:22:@49476.4]
    .clock(RetimeWrapper_171_clock),
    .reset(RetimeWrapper_171_reset),
    .io_flow(RetimeWrapper_171_io_flow),
    .io_in(RetimeWrapper_171_io_in),
    .io_out(RetimeWrapper_171_io_out)
  );
  RetimeWrapper_242 RetimeWrapper_172 ( // @[package.scala 93:22:@49497.4]
    .clock(RetimeWrapper_172_clock),
    .reset(RetimeWrapper_172_reset),
    .io_flow(RetimeWrapper_172_io_flow),
    .io_in(RetimeWrapper_172_io_in),
    .io_out(RetimeWrapper_172_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_173 ( // @[package.scala 93:22:@49506.4]
    .clock(RetimeWrapper_173_clock),
    .reset(RetimeWrapper_173_reset),
    .io_flow(RetimeWrapper_173_io_flow),
    .io_in(RetimeWrapper_173_io_in),
    .io_out(RetimeWrapper_173_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_174 ( // @[package.scala 93:22:@49520.4]
    .clock(RetimeWrapper_174_clock),
    .reset(RetimeWrapper_174_reset),
    .io_flow(RetimeWrapper_174_io_flow),
    .io_in(RetimeWrapper_174_io_in),
    .io_out(RetimeWrapper_174_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_175 ( // @[package.scala 93:22:@49541.4]
    .clock(RetimeWrapper_175_clock),
    .reset(RetimeWrapper_175_reset),
    .io_flow(RetimeWrapper_175_io_flow),
    .io_in(RetimeWrapper_175_io_in),
    .io_out(RetimeWrapper_175_io_out)
  );
  RetimeWrapper_457 RetimeWrapper_176 ( // @[package.scala 93:22:@49550.4]
    .clock(RetimeWrapper_176_clock),
    .reset(RetimeWrapper_176_reset),
    .io_flow(RetimeWrapper_176_io_flow),
    .io_in(RetimeWrapper_176_io_in),
    .io_out(RetimeWrapper_176_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_177 ( // @[package.scala 93:22:@49564.4]
    .clock(RetimeWrapper_177_clock),
    .reset(RetimeWrapper_177_reset),
    .io_flow(RetimeWrapper_177_io_flow),
    .io_in(RetimeWrapper_177_io_in),
    .io_out(RetimeWrapper_177_io_out)
  );
  RetimeWrapper_457 RetimeWrapper_178 ( // @[package.scala 93:22:@49585.4]
    .clock(RetimeWrapper_178_clock),
    .reset(RetimeWrapper_178_reset),
    .io_flow(RetimeWrapper_178_io_flow),
    .io_in(RetimeWrapper_178_io_in),
    .io_out(RetimeWrapper_178_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_179 ( // @[package.scala 93:22:@49594.4]
    .clock(RetimeWrapper_179_clock),
    .reset(RetimeWrapper_179_reset),
    .io_flow(RetimeWrapper_179_io_flow),
    .io_in(RetimeWrapper_179_io_in),
    .io_out(RetimeWrapper_179_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_180 ( // @[package.scala 93:22:@49603.4]
    .clock(RetimeWrapper_180_clock),
    .reset(RetimeWrapper_180_reset),
    .io_flow(RetimeWrapper_180_io_flow),
    .io_in(RetimeWrapper_180_io_in),
    .io_out(RetimeWrapper_180_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_181 ( // @[package.scala 93:22:@49617.4]
    .clock(RetimeWrapper_181_clock),
    .reset(RetimeWrapper_181_reset),
    .io_flow(RetimeWrapper_181_io_flow),
    .io_in(RetimeWrapper_181_io_in),
    .io_out(RetimeWrapper_181_io_out)
  );
  RetimeWrapper_457 RetimeWrapper_182 ( // @[package.scala 93:22:@49638.4]
    .clock(RetimeWrapper_182_clock),
    .reset(RetimeWrapper_182_reset),
    .io_flow(RetimeWrapper_182_io_flow),
    .io_in(RetimeWrapper_182_io_in),
    .io_out(RetimeWrapper_182_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_183 ( // @[package.scala 93:22:@49647.4]
    .clock(RetimeWrapper_183_clock),
    .reset(RetimeWrapper_183_reset),
    .io_flow(RetimeWrapper_183_io_flow),
    .io_in(RetimeWrapper_183_io_in),
    .io_out(RetimeWrapper_183_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_184 ( // @[package.scala 93:22:@49661.4]
    .clock(RetimeWrapper_184_clock),
    .reset(RetimeWrapper_184_reset),
    .io_flow(RetimeWrapper_184_io_flow),
    .io_in(RetimeWrapper_184_io_in),
    .io_out(RetimeWrapper_184_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_185 ( // @[package.scala 93:22:@49682.4]
    .clock(RetimeWrapper_185_clock),
    .reset(RetimeWrapper_185_reset),
    .io_flow(RetimeWrapper_185_io_flow),
    .io_in(RetimeWrapper_185_io_in),
    .io_out(RetimeWrapper_185_io_out)
  );
  RetimeWrapper_457 RetimeWrapper_186 ( // @[package.scala 93:22:@49691.4]
    .clock(RetimeWrapper_186_clock),
    .reset(RetimeWrapper_186_reset),
    .io_flow(RetimeWrapper_186_io_flow),
    .io_in(RetimeWrapper_186_io_in),
    .io_out(RetimeWrapper_186_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_187 ( // @[package.scala 93:22:@49705.4]
    .clock(RetimeWrapper_187_clock),
    .reset(RetimeWrapper_187_reset),
    .io_flow(RetimeWrapper_187_io_flow),
    .io_in(RetimeWrapper_187_io_in),
    .io_out(RetimeWrapper_187_io_out)
  );
  RetimeWrapper_457 RetimeWrapper_188 ( // @[package.scala 93:22:@49726.4]
    .clock(RetimeWrapper_188_clock),
    .reset(RetimeWrapper_188_reset),
    .io_flow(RetimeWrapper_188_io_flow),
    .io_in(RetimeWrapper_188_io_in),
    .io_out(RetimeWrapper_188_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_189 ( // @[package.scala 93:22:@49735.4]
    .clock(RetimeWrapper_189_clock),
    .reset(RetimeWrapper_189_reset),
    .io_flow(RetimeWrapper_189_io_flow),
    .io_in(RetimeWrapper_189_io_in),
    .io_out(RetimeWrapper_189_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_190 ( // @[package.scala 93:22:@49749.4]
    .clock(RetimeWrapper_190_clock),
    .reset(RetimeWrapper_190_reset),
    .io_flow(RetimeWrapper_190_io_flow),
    .io_in(RetimeWrapper_190_io_in),
    .io_out(RetimeWrapper_190_io_out)
  );
  RetimeWrapper_252 RetimeWrapper_191 ( // @[package.scala 93:22:@49770.4]
    .clock(RetimeWrapper_191_clock),
    .reset(RetimeWrapper_191_reset),
    .io_flow(RetimeWrapper_191_io_flow),
    .io_in(RetimeWrapper_191_io_in),
    .io_out(RetimeWrapper_191_io_out)
  );
  RetimeWrapper_457 RetimeWrapper_192 ( // @[package.scala 93:22:@49779.4]
    .clock(RetimeWrapper_192_clock),
    .reset(RetimeWrapper_192_reset),
    .io_flow(RetimeWrapper_192_io_flow),
    .io_in(RetimeWrapper_192_io_in),
    .io_out(RetimeWrapper_192_io_out)
  );
  RetimeWrapper_456 RetimeWrapper_193 ( // @[package.scala 93:22:@49793.4]
    .clock(RetimeWrapper_193_clock),
    .reset(RetimeWrapper_193_reset),
    .io_flow(RetimeWrapper_193_io_flow),
    .io_in(RetimeWrapper_193_io_in),
    .io_out(RetimeWrapper_193_io_out)
  );
  x815_x23 x948_x25_1 ( // @[Math.scala 150:24:@49826.4]
    .io_a(x948_x25_1_io_a),
    .io_b(x948_x25_1_io_b),
    .io_result(x948_x25_1_io_result)
  );
  x815_x23 x949_x26_1 ( // @[Math.scala 150:24:@49836.4]
    .io_a(x949_x26_1_io_a),
    .io_b(x949_x26_1_io_b),
    .io_result(x949_x26_1_io_result)
  );
  x815_x23 x950_sum_1 ( // @[Math.scala 150:24:@49846.4]
    .io_a(x950_sum_1_io_a),
    .io_b(x950_sum_1_io_b),
    .io_result(x950_sum_1_io_result)
  );
  x951_div x951_div_1 ( // @[Math.scala 327:24:@49858.4]
    .clock(x951_div_1_clock),
    .reset(x951_div_1_reset),
    .io_a(x951_div_1_io_a),
    .io_flow(x951_div_1_io_flow),
    .io_result(x951_div_1_io_result)
  );
  x815_x23 x954_x25_1 ( // @[Math.scala 150:24:@49878.4]
    .io_a(x954_x25_1_io_a),
    .io_b(x954_x25_1_io_b),
    .io_result(x954_x25_1_io_result)
  );
  x815_x23 x955_x26_1 ( // @[Math.scala 150:24:@49888.4]
    .io_a(x955_x26_1_io_a),
    .io_b(x955_x26_1_io_b),
    .io_result(x955_x26_1_io_result)
  );
  x815_x23 x956_sum_1 ( // @[Math.scala 150:24:@49898.4]
    .io_a(x956_sum_1_io_a),
    .io_b(x956_sum_1_io_b),
    .io_result(x956_sum_1_io_result)
  );
  x951_div x957_div_1 ( // @[Math.scala 327:24:@49910.4]
    .clock(x957_div_1_clock),
    .reset(x957_div_1_reset),
    .io_a(x957_div_1_io_a),
    .io_flow(x957_div_1_io_flow),
    .io_result(x957_div_1_io_result)
  );
  x815_x23 x960_x25_1 ( // @[Math.scala 150:24:@49930.4]
    .io_a(x960_x25_1_io_a),
    .io_b(x960_x25_1_io_b),
    .io_result(x960_x25_1_io_result)
  );
  x815_x23 x961_x26_1 ( // @[Math.scala 150:24:@49940.4]
    .io_a(x961_x26_1_io_a),
    .io_b(x961_x26_1_io_b),
    .io_result(x961_x26_1_io_result)
  );
  x815_x23 x962_sum_1 ( // @[Math.scala 150:24:@49950.4]
    .io_a(x962_sum_1_io_a),
    .io_b(x962_sum_1_io_b),
    .io_result(x962_sum_1_io_result)
  );
  x951_div x963_div_1 ( // @[Math.scala 327:24:@49962.4]
    .clock(x963_div_1_clock),
    .reset(x963_div_1_reset),
    .io_a(x963_div_1_io_a),
    .io_flow(x963_div_1_io_flow),
    .io_result(x963_div_1_io_result)
  );
  x815_x23 x966_x25_1 ( // @[Math.scala 150:24:@49984.4]
    .io_a(x966_x25_1_io_a),
    .io_b(x966_x25_1_io_b),
    .io_result(x966_x25_1_io_result)
  );
  x815_x23 x967_x26_1 ( // @[Math.scala 150:24:@49994.4]
    .io_a(x967_x26_1_io_a),
    .io_b(x967_x26_1_io_b),
    .io_result(x967_x26_1_io_result)
  );
  x815_x23 x968_sum_1 ( // @[Math.scala 150:24:@50004.4]
    .io_a(x968_sum_1_io_a),
    .io_b(x968_sum_1_io_b),
    .io_result(x968_sum_1_io_result)
  );
  x951_div x969_div_1 ( // @[Math.scala 327:24:@50016.4]
    .clock(x969_div_1_clock),
    .reset(x969_div_1_reset),
    .io_a(x969_div_1_io_a),
    .io_flow(x969_div_1_io_flow),
    .io_result(x969_div_1_io_result)
  );
  x815_x23 x971_x25_1 ( // @[Math.scala 150:24:@50031.4]
    .io_a(x971_x25_1_io_a),
    .io_b(x971_x25_1_io_b),
    .io_result(x971_x25_1_io_result)
  );
  x815_x23 x972_x26_1 ( // @[Math.scala 150:24:@50041.4]
    .io_a(x972_x26_1_io_a),
    .io_b(x972_x26_1_io_b),
    .io_result(x972_x26_1_io_result)
  );
  x815_x23 x973_sum_1 ( // @[Math.scala 150:24:@50051.4]
    .io_a(x973_sum_1_io_a),
    .io_b(x973_sum_1_io_b),
    .io_result(x973_sum_1_io_result)
  );
  x951_div x974_div_1 ( // @[Math.scala 327:24:@50063.4]
    .clock(x974_div_1_clock),
    .reset(x974_div_1_reset),
    .io_a(x974_div_1_io_a),
    .io_flow(x974_div_1_io_flow),
    .io_result(x974_div_1_io_result)
  );
  x815_x23 x976_x25_1 ( // @[Math.scala 150:24:@50078.4]
    .io_a(x976_x25_1_io_a),
    .io_b(x976_x25_1_io_b),
    .io_result(x976_x25_1_io_result)
  );
  x815_x23 x977_x26_1 ( // @[Math.scala 150:24:@50088.4]
    .io_a(x977_x26_1_io_a),
    .io_b(x977_x26_1_io_b),
    .io_result(x977_x26_1_io_result)
  );
  x815_x23 x978_sum_1 ( // @[Math.scala 150:24:@50098.4]
    .io_a(x978_sum_1_io_a),
    .io_b(x978_sum_1_io_b),
    .io_result(x978_sum_1_io_result)
  );
  x951_div x979_div_1 ( // @[Math.scala 327:24:@50110.4]
    .clock(x979_div_1_clock),
    .reset(x979_div_1_reset),
    .io_a(x979_div_1_io_a),
    .io_flow(x979_div_1_io_flow),
    .io_result(x979_div_1_io_result)
  );
  x815_x23 x981_x25_1 ( // @[Math.scala 150:24:@50125.4]
    .io_a(x981_x25_1_io_a),
    .io_b(x981_x25_1_io_b),
    .io_result(x981_x25_1_io_result)
  );
  x815_x23 x982_x26_1 ( // @[Math.scala 150:24:@50135.4]
    .io_a(x982_x26_1_io_a),
    .io_b(x982_x26_1_io_b),
    .io_result(x982_x26_1_io_result)
  );
  x815_x23 x983_sum_1 ( // @[Math.scala 150:24:@50145.4]
    .io_a(x983_sum_1_io_a),
    .io_b(x983_sum_1_io_b),
    .io_result(x983_sum_1_io_result)
  );
  x951_div x984_div_1 ( // @[Math.scala 327:24:@50157.4]
    .clock(x984_div_1_clock),
    .reset(x984_div_1_reset),
    .io_a(x984_div_1_io_a),
    .io_flow(x984_div_1_io_flow),
    .io_result(x984_div_1_io_result)
  );
  x815_x23 x987_x25_1 ( // @[Math.scala 150:24:@50177.4]
    .io_a(x987_x25_1_io_a),
    .io_b(x987_x25_1_io_b),
    .io_result(x987_x25_1_io_result)
  );
  x815_x23 x988_x26_1 ( // @[Math.scala 150:24:@50187.4]
    .io_a(x988_x26_1_io_a),
    .io_b(x988_x26_1_io_b),
    .io_result(x988_x26_1_io_result)
  );
  x815_x23 x989_sum_1 ( // @[Math.scala 150:24:@50197.4]
    .io_a(x989_sum_1_io_a),
    .io_b(x989_sum_1_io_b),
    .io_result(x989_sum_1_io_result)
  );
  x951_div x990_div_1 ( // @[Math.scala 327:24:@50209.4]
    .clock(x990_div_1_clock),
    .reset(x990_div_1_reset),
    .io_a(x990_div_1_io_a),
    .io_flow(x990_div_1_io_flow),
    .io_result(x990_div_1_io_result)
  );
  RetimeWrapper_514 RetimeWrapper_194 ( // @[package.scala 93:22:@50237.4]
    .clock(RetimeWrapper_194_clock),
    .reset(RetimeWrapper_194_reset),
    .io_flow(RetimeWrapper_194_io_flow),
    .io_in(RetimeWrapper_194_io_in),
    .io_out(RetimeWrapper_194_io_out)
  );
  RetimeWrapper_515 RetimeWrapper_195 ( // @[package.scala 93:22:@50246.4]
    .clock(RetimeWrapper_195_clock),
    .reset(RetimeWrapper_195_reset),
    .io_flow(RetimeWrapper_195_io_flow),
    .io_in(RetimeWrapper_195_io_in),
    .io_out(RetimeWrapper_195_io_out)
  );
  RetimeWrapper_515 RetimeWrapper_196 ( // @[package.scala 93:22:@50255.4]
    .clock(RetimeWrapper_196_clock),
    .reset(RetimeWrapper_196_reset),
    .io_flow(RetimeWrapper_196_io_flow),
    .io_in(RetimeWrapper_196_io_in),
    .io_out(RetimeWrapper_196_io_out)
  );
  RetimeWrapper_515 RetimeWrapper_197 ( // @[package.scala 93:22:@50264.4]
    .clock(RetimeWrapper_197_clock),
    .reset(RetimeWrapper_197_reset),
    .io_flow(RetimeWrapper_197_io_flow),
    .io_in(RetimeWrapper_197_io_in),
    .io_out(RetimeWrapper_197_io_out)
  );
  assign b522 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 62:18:@44949.4]
  assign b523 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 63:18:@44950.4]
  assign _T_207 = b522 & b523; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 69:30:@45324.4]
  assign _T_208 = _T_207 & io_sigsIn_datapathEn; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 69:37:@45325.4]
  assign _T_212 = io_in_x511_TID == 8'h0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 71:76:@45330.4]
  assign _T_213 = _T_208 & _T_212; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 71:62:@45331.4]
  assign _T_215 = io_in_x511_TDEST == 8'h0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 71:101:@45332.4]
  assign x1061_x526_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@45341.4 package.scala 96:25:@45342.4]
  assign b520_number = __io_result; // @[Math.scala 712:22:@44934.4 Math.scala 713:14:@44935.4]
  assign _T_255 = $signed(b520_number); // @[Math.scala 499:52:@45369.4]
  assign x530 = $signed(32'sh1) == $signed(_T_255); // @[Math.scala 499:44:@45377.4]
  assign x531 = $signed(32'sh2) == $signed(_T_255); // @[Math.scala 499:44:@45384.4]
  assign x532 = $signed(32'sh3) == $signed(_T_255); // @[Math.scala 499:44:@45391.4]
  assign _T_302 = x530 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@45403.4]
  assign _T_304 = x531 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@45404.4]
  assign _T_306 = x532 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@45405.4]
  assign _T_308 = _T_302 | _T_304; // @[Mux.scala 19:72:@45407.4]
  assign x533_number = _T_308 | _T_306; // @[Mux.scala 19:72:@45408.4]
  assign _T_320 = $signed(x533_number); // @[Math.scala 406:49:@45418.4]
  assign _T_322 = $signed(_T_320) & $signed(32'sh3); // @[Math.scala 406:56:@45420.4]
  assign _T_323 = $signed(_T_322); // @[Math.scala 406:56:@45421.4]
  assign _T_328 = x533_number[31]; // @[FixedPoint.scala 50:25:@45427.4]
  assign _T_332 = _T_328 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@45429.4]
  assign _T_333 = x533_number[31:2]; // @[FixedPoint.scala 18:52:@45430.4]
  assign b521_number = __1_io_result; // @[Math.scala 712:22:@44946.4 Math.scala 713:14:@44947.4]
  assign _T_338 = b521_number[31]; // @[FixedPoint.scala 50:25:@45436.4]
  assign _T_342 = _T_338 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@45438.4]
  assign _T_343 = b521_number[31:2]; // @[FixedPoint.scala 18:52:@45439.4]
  assign _T_368 = ~ io_sigsIn_break; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 114:101:@45500.4]
  assign _T_372 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@45508.4 package.scala 96:25:@45509.4]
  assign _T_374 = io_rr ? _T_372 : 1'h0; // @[implicits.scala 55:10:@45510.4]
  assign _T_375 = _T_368 & _T_374; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 114:118:@45511.4]
  assign _T_377 = _T_375 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 114:205:@45513.4]
  assign _T_378 = _T_377 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 114:224:@45514.4]
  assign x1065_b522_D8 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@45486.4 package.scala 96:25:@45487.4]
  assign _T_379 = _T_378 & x1065_b522_D8; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 114:250:@45515.4]
  assign x1062_b523_D8 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@45459.4 package.scala 96:25:@45460.4]
  assign x545_rdcol_number = x545_rdcol_1_io_result; // @[Math.scala 154:22:@45532.4 Math.scala 155:14:@45533.4]
  assign _T_392 = x545_rdcol_number[31]; // @[FixedPoint.scala 50:25:@45539.4]
  assign _T_396 = _T_392 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@45541.4]
  assign _T_397 = x545_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@45542.4]
  assign _T_420 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@45593.4 package.scala 96:25:@45594.4]
  assign _T_422 = io_rr ? _T_420 : 1'h0; // @[implicits.scala 55:10:@45595.4]
  assign _T_423 = _T_368 & _T_422; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 133:118:@45596.4]
  assign _T_425 = _T_423 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 133:205:@45598.4]
  assign _T_426 = _T_425 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 133:224:@45599.4]
  assign _T_427 = _T_426 & x1065_b522_D8; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 133:250:@45600.4]
  assign x554_rdcol_number = x554_rdcol_1_io_result; // @[Math.scala 154:22:@45617.4 Math.scala 155:14:@45618.4]
  assign _T_440 = x554_rdcol_number[31]; // @[FixedPoint.scala 50:25:@45624.4]
  assign _T_444 = _T_440 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@45626.4]
  assign _T_445 = x554_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@45627.4]
  assign _T_465 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@45669.4 package.scala 96:25:@45670.4]
  assign _T_467 = io_rr ? _T_465 : 1'h0; // @[implicits.scala 55:10:@45671.4]
  assign _T_468 = _T_368 & _T_467; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 150:118:@45672.4]
  assign _T_470 = _T_468 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 150:205:@45674.4]
  assign _T_471 = _T_470 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 150:224:@45675.4]
  assign _T_472 = _T_471 & x1065_b522_D8; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 150:250:@45676.4]
  assign x563_rdcol_number = x563_rdcol_1_io_result; // @[Math.scala 154:22:@45693.4 Math.scala 155:14:@45694.4]
  assign _T_485 = x563_rdcol_number[31]; // @[FixedPoint.scala 50:25:@45700.4]
  assign _T_489 = _T_485 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@45702.4]
  assign _T_490 = x563_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@45703.4]
  assign _T_510 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@45745.4 package.scala 96:25:@45746.4]
  assign _T_512 = io_rr ? _T_510 : 1'h0; // @[implicits.scala 55:10:@45747.4]
  assign _T_513 = _T_368 & _T_512; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 167:118:@45748.4]
  assign _T_515 = _T_513 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 167:205:@45750.4]
  assign _T_516 = _T_515 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 167:224:@45751.4]
  assign _T_517 = _T_516 & x1065_b522_D8; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 167:250:@45752.4]
  assign x572_rdrow_number = x572_rdrow_1_io_result; // @[Math.scala 154:22:@45769.4 Math.scala 155:14:@45770.4]
  assign _T_532 = $signed(x572_rdrow_number); // @[Math.scala 499:52:@45776.4]
  assign x574 = $signed(32'sh1) == $signed(_T_532); // @[Math.scala 499:44:@45784.4]
  assign x575 = $signed(32'sh2) == $signed(_T_532); // @[Math.scala 499:44:@45791.4]
  assign x576 = $signed(32'sh3) == $signed(_T_532); // @[Math.scala 499:44:@45798.4]
  assign _T_579 = x574 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@45810.4]
  assign _T_581 = x575 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@45811.4]
  assign _T_583 = x576 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@45812.4]
  assign _T_585 = _T_579 | _T_581; // @[Mux.scala 19:72:@45814.4]
  assign x577_number = _T_585 | _T_583; // @[Mux.scala 19:72:@45815.4]
  assign _T_599 = $signed(x577_number); // @[Math.scala 406:49:@45827.4]
  assign _T_601 = $signed(_T_599) & $signed(32'sh3); // @[Math.scala 406:56:@45829.4]
  assign _T_602 = $signed(_T_601); // @[Math.scala 406:56:@45830.4]
  assign _T_607 = x577_number[31]; // @[FixedPoint.scala 50:25:@45836.4]
  assign _T_611 = _T_607 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@45838.4]
  assign _T_612 = x577_number[31:2]; // @[FixedPoint.scala 18:52:@45839.4]
  assign _T_638 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@45899.4 package.scala 96:25:@45900.4]
  assign _T_640 = io_rr ? _T_638 : 1'h0; // @[implicits.scala 55:10:@45901.4]
  assign _T_641 = _T_368 & _T_640; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 208:166:@45902.4]
  assign _T_643 = _T_641 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 208:253:@45904.4]
  assign _T_644 = _T_643 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 208:272:@45905.4]
  assign _T_645 = _T_644 & x1065_b522_D8; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 208:298:@45906.4]
  assign _T_666 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@45954.4 package.scala 96:25:@45955.4]
  assign _T_668 = io_rr ? _T_666 : 1'h0; // @[implicits.scala 55:10:@45956.4]
  assign _T_669 = _T_368 & _T_668; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 221:166:@45957.4]
  assign _T_671 = _T_669 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 221:253:@45959.4]
  assign _T_672 = _T_671 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 221:272:@45960.4]
  assign _T_673 = _T_672 & x1065_b522_D8; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 221:298:@45961.4]
  assign _T_694 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@46009.4 package.scala 96:25:@46010.4]
  assign _T_696 = io_rr ? _T_694 : 1'h0; // @[implicits.scala 55:10:@46011.4]
  assign _T_697 = _T_368 & _T_696; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 234:166:@46012.4]
  assign _T_699 = _T_697 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 234:253:@46014.4]
  assign _T_700 = _T_699 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 234:272:@46015.4]
  assign _T_701 = _T_700 & x1065_b522_D8; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 234:298:@46016.4]
  assign _T_722 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@46064.4 package.scala 96:25:@46065.4]
  assign _T_724 = io_rr ? _T_722 : 1'h0; // @[implicits.scala 55:10:@46066.4]
  assign _T_725 = _T_368 & _T_724; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 247:166:@46067.4]
  assign _T_727 = _T_725 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 247:253:@46069.4]
  assign _T_728 = _T_727 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 247:272:@46070.4]
  assign _T_729 = _T_728 & x1065_b522_D8; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 247:298:@46071.4]
  assign x1084_x572_rdrow_D11_number = RetimeWrapper_31_io_out; // @[package.scala 96:25:@46085.4 package.scala 96:25:@46086.4]
  assign _T_741 = $signed(x1084_x572_rdrow_D11_number); // @[Math.scala 406:49:@46092.4]
  assign _T_743 = $signed(_T_741) & $signed(32'sh3); // @[Math.scala 406:56:@46094.4]
  assign _T_744 = $signed(_T_743); // @[Math.scala 406:56:@46095.4]
  assign x1053_number = $unsigned(_T_744); // @[implicits.scala 133:21:@46096.4]
  assign x603 = $signed(_T_741) < $signed(32'sh0); // @[Math.scala 465:44:@46104.4]
  assign x1085_x563_rdcol_D11_number = RetimeWrapper_32_io_out; // @[package.scala 96:25:@46112.4 package.scala 96:25:@46113.4]
  assign _T_762 = $signed(x1085_x563_rdcol_D11_number); // @[Math.scala 465:37:@46118.4]
  assign x604 = $signed(_T_762) < $signed(32'sh0); // @[Math.scala 465:44:@46120.4]
  assign x605 = x603 | x604; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 260:24:@46123.4]
  assign _T_776 = $signed(x1053_number); // @[Math.scala 406:49:@46132.4]
  assign _T_778 = $signed(_T_776) & $signed(32'sh3); // @[Math.scala 406:56:@46134.4]
  assign _T_779 = $signed(_T_778); // @[Math.scala 406:56:@46135.4]
  assign _T_784 = x1053_number[31]; // @[FixedPoint.scala 50:25:@46141.4]
  assign _T_788 = _T_784 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@46143.4]
  assign _T_789 = x1053_number[31:2]; // @[FixedPoint.scala 18:52:@46144.4]
  assign _T_824 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@46214.4 package.scala 96:25:@46215.4]
  assign _T_826 = io_rr ? _T_824 : 1'h0; // @[implicits.scala 55:10:@46216.4]
  assign _T_827 = _T_368 & _T_826; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 283:194:@46217.4]
  assign x1088_x606_D1 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@46182.4 package.scala 96:25:@46183.4]
  assign _T_828 = _T_827 & x1088_x606_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 283:282:@46218.4]
  assign x1089_b522_D13 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@46191.4 package.scala 96:25:@46192.4]
  assign _T_829 = _T_828 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 283:291:@46219.4]
  assign x1087_b523_D13 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@46173.4 package.scala 96:25:@46174.4]
  assign x1091_x554_rdcol_D11_number = RetimeWrapper_39_io_out; // @[package.scala 96:25:@46235.4 package.scala 96:25:@46236.4]
  assign _T_840 = $signed(x1091_x554_rdcol_D11_number); // @[Math.scala 465:37:@46241.4]
  assign x615 = $signed(_T_840) < $signed(32'sh0); // @[Math.scala 465:44:@46243.4]
  assign x616 = x603 | x615; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 291:24:@46246.4]
  assign _T_871 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@46290.4 package.scala 96:25:@46291.4]
  assign _T_873 = io_rr ? _T_871 : 1'h0; // @[implicits.scala 55:10:@46292.4]
  assign _T_874 = _T_368 & _T_873; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 310:194:@46293.4]
  assign x1093_x617_D1 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@46276.4 package.scala 96:25:@46277.4]
  assign _T_875 = _T_874 & x1093_x617_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 310:282:@46294.4]
  assign _T_876 = _T_875 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 310:291:@46295.4]
  assign x1094_x545_rdcol_D11_number = RetimeWrapper_43_io_out; // @[package.scala 96:25:@46311.4 package.scala 96:25:@46312.4]
  assign _T_889 = $signed(x1094_x545_rdcol_D11_number); // @[Math.scala 465:37:@46319.4]
  assign x623 = $signed(_T_889) < $signed(32'sh0); // @[Math.scala 465:44:@46321.4]
  assign x624 = x603 | x623; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 320:59:@46324.4]
  assign _T_920 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@46368.4 package.scala 96:25:@46369.4]
  assign _T_922 = io_rr ? _T_920 : 1'h0; // @[implicits.scala 55:10:@46370.4]
  assign _T_923 = _T_368 & _T_922; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 333:194:@46371.4]
  assign x1096_x625_D1 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@46354.4 package.scala 96:25:@46355.4]
  assign _T_924 = _T_923 & x1096_x625_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 333:282:@46372.4]
  assign _T_925 = _T_924 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 333:291:@46373.4]
  assign x1097_b521_D11_number = RetimeWrapper_47_io_out; // @[package.scala 96:25:@46389.4 package.scala 96:25:@46390.4]
  assign _T_936 = $signed(x1097_b521_D11_number); // @[Math.scala 465:37:@46395.4]
  assign x631 = $signed(_T_936) < $signed(32'sh0); // @[Math.scala 465:44:@46397.4]
  assign x1098_x631_D1 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@46405.4 package.scala 96:25:@46406.4]
  assign x632 = x603 | x1098_x631_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 343:59:@46409.4]
  assign _T_970 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@46453.4 package.scala 96:25:@46454.4]
  assign _T_972 = io_rr ? _T_970 : 1'h0; // @[implicits.scala 55:10:@46455.4]
  assign _T_973 = _T_368 & _T_972; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 356:194:@46456.4]
  assign x1100_x633_D1 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@46439.4 package.scala 96:25:@46440.4]
  assign _T_974 = _T_973 & x1100_x633_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 356:282:@46457.4]
  assign _T_975 = _T_974 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 356:291:@46458.4]
  assign x639_rdcol_number = x639_rdcol_1_io_result; // @[Math.scala 154:22:@46477.4 Math.scala 155:14:@46478.4]
  assign _T_990 = $signed(x639_rdcol_number); // @[Math.scala 465:37:@46483.4]
  assign x640 = $signed(_T_990) < $signed(32'sh0); // @[Math.scala 465:44:@46485.4]
  assign x641 = x603 | x640; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 364:59:@46488.4]
  assign _T_1000 = x639_rdcol_number[31]; // @[FixedPoint.scala 50:25:@46495.4]
  assign _T_1004 = _T_1000 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@46497.4]
  assign _T_1005 = x639_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@46498.4]
  assign _T_1028 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@46532.4 package.scala 96:25:@46533.4]
  assign _T_1030 = io_rr ? _T_1028 : 1'h0; // @[implicits.scala 55:10:@46534.4]
  assign _T_1031 = _T_368 & _T_1030; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 377:194:@46535.4]
  assign x1101_x642_D1 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@46518.4 package.scala 96:25:@46519.4]
  assign _T_1032 = _T_1031 & x1101_x642_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 377:282:@46536.4]
  assign _T_1033 = _T_1032 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 377:291:@46537.4]
  assign x651_rdcol_number = x651_rdcol_1_io_result; // @[Math.scala 154:22:@46556.4 Math.scala 155:14:@46557.4]
  assign _T_1048 = $signed(x651_rdcol_number); // @[Math.scala 465:37:@46562.4]
  assign x652 = $signed(_T_1048) < $signed(32'sh0); // @[Math.scala 465:44:@46564.4]
  assign x653 = x603 | x652; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 385:59:@46567.4]
  assign _T_1058 = x651_rdcol_number[31]; // @[FixedPoint.scala 50:25:@46574.4]
  assign _T_1062 = _T_1058 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@46576.4]
  assign _T_1063 = x651_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@46577.4]
  assign _T_1086 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@46611.4 package.scala 96:25:@46612.4]
  assign _T_1088 = io_rr ? _T_1086 : 1'h0; // @[implicits.scala 55:10:@46613.4]
  assign _T_1089 = _T_368 & _T_1088; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 398:194:@46614.4]
  assign x1102_x654_D1 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@46597.4 package.scala 96:25:@46598.4]
  assign _T_1090 = _T_1089 & x1102_x654_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 398:282:@46615.4]
  assign _T_1091 = _T_1090 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 398:291:@46616.4]
  assign x1103_b520_D11_number = RetimeWrapper_56_io_out; // @[package.scala 96:25:@46632.4 package.scala 96:25:@46633.4]
  assign _T_1104 = $signed(x1103_b520_D11_number); // @[Math.scala 406:49:@46639.4]
  assign _T_1106 = $signed(_T_1104) & $signed(32'sh3); // @[Math.scala 406:56:@46641.4]
  assign _T_1107 = $signed(_T_1106); // @[Math.scala 406:56:@46642.4]
  assign x1055_number = $unsigned(_T_1107); // @[implicits.scala 133:21:@46643.4]
  assign x664 = $signed(_T_1104) < $signed(32'sh0); // @[Math.scala 465:44:@46651.4]
  assign x1104_x664_D1 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@46659.4 package.scala 96:25:@46660.4]
  assign x665 = x1104_x664_D1 | x604; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 410:25:@46663.4]
  assign _T_1131 = $signed(x1055_number); // @[Math.scala 406:49:@46672.4]
  assign _T_1133 = $signed(_T_1131) & $signed(32'sh3); // @[Math.scala 406:56:@46674.4]
  assign _T_1134 = $signed(_T_1133); // @[Math.scala 406:56:@46675.4]
  assign _T_1139 = x1055_number[31]; // @[FixedPoint.scala 50:25:@46681.4]
  assign _T_1143 = _T_1139 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@46683.4]
  assign _T_1144 = x1055_number[31:2]; // @[FixedPoint.scala 18:52:@46684.4]
  assign _T_1175 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@46738.4 package.scala 96:25:@46739.4]
  assign _T_1177 = io_rr ? _T_1175 : 1'h0; // @[implicits.scala 55:10:@46740.4]
  assign _T_1178 = _T_368 & _T_1177; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 437:194:@46741.4]
  assign x1106_x666_D1 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@46715.4 package.scala 96:25:@46716.4]
  assign _T_1179 = _T_1178 & x1106_x666_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 437:282:@46742.4]
  assign _T_1180 = _T_1179 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 437:291:@46743.4]
  assign x675 = x1104_x664_D1 | x615; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 441:60:@46754.4]
  assign _T_1208 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@46789.4 package.scala 96:25:@46790.4]
  assign _T_1210 = io_rr ? _T_1208 : 1'h0; // @[implicits.scala 55:10:@46791.4]
  assign _T_1211 = _T_368 & _T_1210; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 452:194:@46792.4]
  assign x1108_x676_D1 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@46775.4 package.scala 96:25:@46776.4]
  assign _T_1212 = _T_1211 & x1108_x676_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 452:282:@46793.4]
  assign _T_1213 = _T_1212 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 452:291:@46794.4]
  assign x682 = x1104_x664_D1 | x623; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 456:60:@46805.4]
  assign _T_1241 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@46840.4 package.scala 96:25:@46841.4]
  assign _T_1243 = io_rr ? _T_1241 : 1'h0; // @[implicits.scala 55:10:@46842.4]
  assign _T_1244 = _T_368 & _T_1243; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 467:194:@46843.4]
  assign x1109_x683_D1 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@46826.4 package.scala 96:25:@46827.4]
  assign _T_1245 = _T_1244 & x1109_x683_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 467:282:@46844.4]
  assign _T_1246 = _T_1245 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 467:291:@46845.4]
  assign x689 = x664 | x631; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 471:59:@46856.4]
  assign _T_1280 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@46909.4 package.scala 96:25:@46910.4]
  assign _T_1282 = io_rr ? _T_1280 : 1'h0; // @[implicits.scala 55:10:@46911.4]
  assign _T_1283 = _T_368 & _T_1282; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 486:194:@46912.4]
  assign x1111_x690_D2 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@46886.4 package.scala 96:25:@46887.4]
  assign _T_1284 = _T_1283 & x1111_x690_D2; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 486:282:@46913.4]
  assign _T_1285 = _T_1284 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 486:291:@46914.4]
  assign x696 = x1104_x664_D1 | x640; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 490:60:@46925.4]
  assign _T_1313 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@46960.4 package.scala 96:25:@46961.4]
  assign _T_1315 = io_rr ? _T_1313 : 1'h0; // @[implicits.scala 55:10:@46962.4]
  assign _T_1316 = _T_368 & _T_1315; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 501:194:@46963.4]
  assign x1113_x697_D1 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@46946.4 package.scala 96:25:@46947.4]
  assign _T_1317 = _T_1316 & x1113_x697_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 501:282:@46964.4]
  assign _T_1318 = _T_1317 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 501:291:@46965.4]
  assign x703 = x1104_x664_D1 | x652; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 505:60:@46976.4]
  assign _T_1346 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@47011.4 package.scala 96:25:@47012.4]
  assign _T_1348 = io_rr ? _T_1346 : 1'h0; // @[implicits.scala 55:10:@47013.4]
  assign _T_1349 = _T_368 & _T_1348; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 516:194:@47014.4]
  assign x1114_x704_D1 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@46997.4 package.scala 96:25:@46998.4]
  assign _T_1350 = _T_1349 & x1114_x704_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 516:282:@47015.4]
  assign _T_1351 = _T_1350 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 516:291:@47016.4]
  assign x710_rdrow_number = x710_rdrow_1_io_result; // @[Math.scala 154:22:@47035.4 Math.scala 155:14:@47036.4]
  assign _T_1368 = $signed(x710_rdrow_number); // @[Math.scala 406:49:@47042.4]
  assign _T_1370 = $signed(_T_1368) & $signed(32'sh3); // @[Math.scala 406:56:@47044.4]
  assign _T_1371 = $signed(_T_1370); // @[Math.scala 406:56:@47045.4]
  assign x1057_number = $unsigned(_T_1371); // @[implicits.scala 133:21:@47046.4]
  assign x712 = $signed(_T_1368) < $signed(32'sh0); // @[Math.scala 465:44:@47054.4]
  assign x713 = x712 | x604; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 526:24:@47057.4]
  assign _T_1392 = $signed(x1057_number); // @[Math.scala 406:49:@47066.4]
  assign _T_1394 = $signed(_T_1392) & $signed(32'sh3); // @[Math.scala 406:56:@47068.4]
  assign _T_1395 = $signed(_T_1394); // @[Math.scala 406:56:@47069.4]
  assign _T_1400 = x1057_number[31]; // @[FixedPoint.scala 50:25:@47075.4]
  assign _T_1404 = _T_1400 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@47077.4]
  assign _T_1405 = x1057_number[31:2]; // @[FixedPoint.scala 18:52:@47078.4]
  assign _T_1431 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@47121.4 package.scala 96:25:@47122.4]
  assign _T_1433 = io_rr ? _T_1431 : 1'h0; // @[implicits.scala 55:10:@47123.4]
  assign _T_1434 = _T_368 & _T_1433; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 543:194:@47124.4]
  assign x1115_x714_D1 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@47098.4 package.scala 96:25:@47099.4]
  assign _T_1435 = _T_1434 & x1115_x714_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 543:282:@47125.4]
  assign _T_1436 = _T_1435 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 543:291:@47126.4]
  assign x723 = x712 | x615; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 553:59:@47137.4]
  assign _T_1466 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@47174.4 package.scala 96:25:@47175.4]
  assign _T_1468 = io_rr ? _T_1466 : 1'h0; // @[implicits.scala 55:10:@47176.4]
  assign _T_1469 = _T_368 & _T_1468; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 566:194:@47177.4]
  assign x1117_x724_D1 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@47160.4 package.scala 96:25:@47161.4]
  assign _T_1470 = _T_1469 & x1117_x724_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 566:282:@47178.4]
  assign _T_1471 = _T_1470 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 566:291:@47179.4]
  assign x730 = x712 | x623; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 570:59:@47190.4]
  assign _T_1499 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@47225.4 package.scala 96:25:@47226.4]
  assign _T_1501 = io_rr ? _T_1499 : 1'h0; // @[implicits.scala 55:10:@47227.4]
  assign _T_1502 = _T_368 & _T_1501; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 581:194:@47228.4]
  assign x1118_x731_D1 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@47211.4 package.scala 96:25:@47212.4]
  assign _T_1503 = _T_1502 & x1118_x731_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 581:282:@47229.4]
  assign _T_1504 = _T_1503 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 581:291:@47230.4]
  assign x737 = x712 | x1098_x631_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 585:59:@47241.4]
  assign _T_1532 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@47276.4 package.scala 96:25:@47277.4]
  assign _T_1534 = io_rr ? _T_1532 : 1'h0; // @[implicits.scala 55:10:@47278.4]
  assign _T_1535 = _T_368 & _T_1534; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 596:194:@47279.4]
  assign x1119_x738_D1 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@47262.4 package.scala 96:25:@47263.4]
  assign _T_1536 = _T_1535 & x1119_x738_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 596:282:@47280.4]
  assign _T_1537 = _T_1536 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 596:291:@47281.4]
  assign x744 = x712 | x640; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 600:59:@47292.4]
  assign _T_1565 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@47327.4 package.scala 96:25:@47328.4]
  assign _T_1567 = io_rr ? _T_1565 : 1'h0; // @[implicits.scala 55:10:@47329.4]
  assign _T_1568 = _T_368 & _T_1567; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 611:194:@47330.4]
  assign x1120_x745_D1 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@47313.4 package.scala 96:25:@47314.4]
  assign _T_1569 = _T_1568 & x1120_x745_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 611:282:@47331.4]
  assign _T_1570 = _T_1569 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 611:291:@47332.4]
  assign x751 = x712 | x652; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 615:59:@47343.4]
  assign _T_1598 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@47378.4 package.scala 96:25:@47379.4]
  assign _T_1600 = io_rr ? _T_1598 : 1'h0; // @[implicits.scala 55:10:@47380.4]
  assign _T_1601 = _T_368 & _T_1600; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 626:194:@47381.4]
  assign x1121_x752_D1 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@47364.4 package.scala 96:25:@47365.4]
  assign _T_1602 = _T_1601 & x1121_x752_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 626:282:@47382.4]
  assign _T_1603 = _T_1602 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 626:291:@47383.4]
  assign x758_rdrow_number = x758_rdrow_1_io_result; // @[Math.scala 154:22:@47402.4 Math.scala 155:14:@47403.4]
  assign _T_1620 = $signed(x758_rdrow_number); // @[Math.scala 406:49:@47409.4]
  assign _T_1622 = $signed(_T_1620) & $signed(32'sh3); // @[Math.scala 406:56:@47411.4]
  assign _T_1623 = $signed(_T_1622); // @[Math.scala 406:56:@47412.4]
  assign x1059_number = $unsigned(_T_1623); // @[implicits.scala 133:21:@47413.4]
  assign x760 = $signed(_T_1620) < $signed(32'sh0); // @[Math.scala 465:44:@47421.4]
  assign x761 = x760 | x604; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 636:24:@47424.4]
  assign _T_1644 = $signed(x1059_number); // @[Math.scala 406:49:@47433.4]
  assign _T_1646 = $signed(_T_1644) & $signed(32'sh3); // @[Math.scala 406:56:@47435.4]
  assign _T_1647 = $signed(_T_1646); // @[Math.scala 406:56:@47436.4]
  assign _T_1652 = x1059_number[31]; // @[FixedPoint.scala 50:25:@47442.4]
  assign _T_1656 = _T_1652 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@47444.4]
  assign _T_1657 = x1059_number[31:2]; // @[FixedPoint.scala 18:52:@47445.4]
  assign _T_1683 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@47488.4 package.scala 96:25:@47489.4]
  assign _T_1685 = io_rr ? _T_1683 : 1'h0; // @[implicits.scala 55:10:@47490.4]
  assign _T_1686 = _T_368 & _T_1685; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 653:194:@47491.4]
  assign x1122_x762_D1 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@47465.4 package.scala 96:25:@47466.4]
  assign _T_1687 = _T_1686 & x1122_x762_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 653:282:@47492.4]
  assign _T_1688 = _T_1687 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 653:291:@47493.4]
  assign x771 = x760 | x615; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 657:24:@47504.4]
  assign _T_1716 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@47539.4 package.scala 96:25:@47540.4]
  assign _T_1718 = io_rr ? _T_1716 : 1'h0; // @[implicits.scala 55:10:@47541.4]
  assign _T_1719 = _T_368 & _T_1718; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 668:194:@47542.4]
  assign x1124_x772_D1 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@47525.4 package.scala 96:25:@47526.4]
  assign _T_1720 = _T_1719 & x1124_x772_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 668:282:@47543.4]
  assign _T_1721 = _T_1720 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 668:291:@47544.4]
  assign x778 = x760 | x623; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 672:24:@47555.4]
  assign _T_1751 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@47592.4 package.scala 96:25:@47593.4]
  assign _T_1753 = io_rr ? _T_1751 : 1'h0; // @[implicits.scala 55:10:@47594.4]
  assign _T_1754 = _T_368 & _T_1753; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 691:194:@47595.4]
  assign x1125_x779_D1 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@47578.4 package.scala 96:25:@47579.4]
  assign _T_1755 = _T_1754 & x1125_x779_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 691:282:@47596.4]
  assign _T_1756 = _T_1755 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 691:291:@47597.4]
  assign x785 = x760 | x1098_x631_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 695:59:@47608.4]
  assign _T_1784 = RetimeWrapper_95_io_out; // @[package.scala 96:25:@47643.4 package.scala 96:25:@47644.4]
  assign _T_1786 = io_rr ? _T_1784 : 1'h0; // @[implicits.scala 55:10:@47645.4]
  assign _T_1787 = _T_368 & _T_1786; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 706:194:@47646.4]
  assign x1126_x786_D1 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@47629.4 package.scala 96:25:@47630.4]
  assign _T_1788 = _T_1787 & x1126_x786_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 706:282:@47647.4]
  assign _T_1789 = _T_1788 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 706:291:@47648.4]
  assign x792 = x760 | x640; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 710:59:@47659.4]
  assign _T_1817 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@47694.4 package.scala 96:25:@47695.4]
  assign _T_1819 = io_rr ? _T_1817 : 1'h0; // @[implicits.scala 55:10:@47696.4]
  assign _T_1820 = _T_368 & _T_1819; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 721:194:@47697.4]
  assign x1127_x793_D1 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@47680.4 package.scala 96:25:@47681.4]
  assign _T_1821 = _T_1820 & x1127_x793_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 721:282:@47698.4]
  assign _T_1822 = _T_1821 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 721:291:@47699.4]
  assign x799 = x760 | x652; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 725:59:@47710.4]
  assign _T_1850 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@47745.4 package.scala 96:25:@47746.4]
  assign _T_1852 = io_rr ? _T_1850 : 1'h0; // @[implicits.scala 55:10:@47747.4]
  assign _T_1853 = _T_368 & _T_1852; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 736:194:@47748.4]
  assign x1128_x800_D1 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@47731.4 package.scala 96:25:@47732.4]
  assign _T_1854 = _T_1853 & x1128_x800_D1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 736:282:@47749.4]
  assign _T_1855 = _T_1854 & x1089_b522_D13; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 736:291:@47750.4]
  assign x621_rd_0_number = x524_lb_0_io_rPort_13_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 306:29:@46279.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 310:410:@46302.4]
  assign _GEN_0 = {{1'd0}, x621_rd_0_number}; // @[Math.scala 450:32:@47762.4]
  assign _T_1861 = _GEN_0 << 1; // @[Math.scala 450:32:@47762.4]
  assign x673_rd_0_number = x524_lb_0_io_rPort_18_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 433:29:@46727.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 437:410:@46750.4]
  assign _GEN_1 = {{1'd0}, x673_rd_0_number}; // @[Math.scala 450:32:@47767.4]
  assign _T_1865 = _GEN_1 << 1; // @[Math.scala 450:32:@47767.4]
  assign x680_rd_0_number = x524_lb_0_io_rPort_15_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 448:29:@46778.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 452:410:@46801.4]
  assign _GEN_2 = {{2'd0}, x680_rd_0_number}; // @[Math.scala 450:32:@47772.4]
  assign _T_1869 = _GEN_2 << 2; // @[Math.scala 450:32:@47772.4]
  assign x687_rd_0_number = x524_lb_0_io_rPort_3_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 463:29:@46829.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 467:410:@46852.4]
  assign _GEN_3 = {{1'd0}, x687_rd_0_number}; // @[Math.scala 450:32:@47777.4]
  assign _T_1873 = _GEN_3 << 1; // @[Math.scala 450:32:@47777.4]
  assign x728_rd_0_number = x524_lb_0_io_rPort_22_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 562:29:@47163.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 566:410:@47186.4]
  assign _GEN_4 = {{1'd0}, x728_rd_0_number}; // @[Math.scala 450:32:@47782.4]
  assign _T_1877 = _GEN_4 << 1; // @[Math.scala 450:32:@47782.4]
  assign x818_sum_number = x818_sum_1_io_result; // @[Math.scala 154:22:@47871.4 Math.scala 155:14:@47872.4]
  assign _T_1913 = x818_sum_number[7:4]; // @[FixedPoint.scala 18:52:@47877.4]
  assign x629_rd_0_number = x524_lb_0_io_rPort_0_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 329:29:@46357.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 333:410:@46380.4]
  assign _GEN_5 = {{1'd0}, x629_rd_0_number}; // @[Math.scala 450:32:@47890.4]
  assign _T_1920 = _GEN_5 << 1; // @[Math.scala 450:32:@47890.4]
  assign _GEN_6 = {{1'd0}, x680_rd_0_number}; // @[Math.scala 450:32:@47895.4]
  assign _T_1924 = _GEN_6 << 1; // @[Math.scala 450:32:@47895.4]
  assign _GEN_7 = {{2'd0}, x687_rd_0_number}; // @[Math.scala 450:32:@47900.4]
  assign _T_1928 = _GEN_7 << 2; // @[Math.scala 450:32:@47900.4]
  assign x694_rd_0_number = x524_lb_0_io_rPort_10_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 482:29:@46898.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 486:410:@46921.4]
  assign _GEN_8 = {{1'd0}, x694_rd_0_number}; // @[Math.scala 450:32:@47905.4]
  assign _T_1932 = _GEN_8 << 1; // @[Math.scala 450:32:@47905.4]
  assign x735_rd_0_number = x524_lb_0_io_rPort_21_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 577:29:@47214.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 581:410:@47237.4]
  assign _GEN_9 = {{1'd0}, x735_rd_0_number}; // @[Math.scala 450:32:@47910.4]
  assign _T_1936 = _GEN_9 << 1; // @[Math.scala 450:32:@47910.4]
  assign x832_sum_number = x832_sum_1_io_result; // @[Math.scala 154:22:@48001.4 Math.scala 155:14:@48002.4]
  assign _T_1974 = x832_sum_number[7:4]; // @[FixedPoint.scala 18:52:@48007.4]
  assign x637_rd_0_number = x524_lb_0_io_rPort_7_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 352:29:@46442.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 356:410:@46465.4]
  assign _GEN_10 = {{1'd0}, x637_rd_0_number}; // @[Math.scala 450:32:@48020.4]
  assign _T_1981 = _GEN_10 << 1; // @[Math.scala 450:32:@48020.4]
  assign _GEN_11 = {{2'd0}, x694_rd_0_number}; // @[Math.scala 450:32:@48025.4]
  assign _T_1985 = _GEN_11 << 2; // @[Math.scala 450:32:@48025.4]
  assign x701_rd_0_number = x524_lb_0_io_rPort_8_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 497:29:@46949.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 501:410:@46972.4]
  assign _GEN_12 = {{1'd0}, x701_rd_0_number}; // @[Math.scala 450:32:@48030.4]
  assign _T_1989 = _GEN_12 << 1; // @[Math.scala 450:32:@48030.4]
  assign x742_rd_0_number = x524_lb_0_io_rPort_5_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 592:29:@47265.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 596:410:@47288.4]
  assign _GEN_13 = {{1'd0}, x742_rd_0_number}; // @[Math.scala 450:32:@48035.4]
  assign _T_1993 = _GEN_13 << 1; // @[Math.scala 450:32:@48035.4]
  assign x845_sum_number = x845_sum_1_io_result; // @[Math.scala 154:22:@48124.4 Math.scala 155:14:@48125.4]
  assign _T_2029 = x845_sum_number[7:4]; // @[FixedPoint.scala 18:52:@48130.4]
  assign x649_rd_0_number = x524_lb_0_io_rPort_12_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 373:29:@46521.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 377:410:@46544.4]
  assign _GEN_14 = {{1'd0}, x649_rd_0_number}; // @[Math.scala 450:32:@48143.4]
  assign _T_2036 = _GEN_14 << 1; // @[Math.scala 450:32:@48143.4]
  assign _GEN_15 = {{2'd0}, x701_rd_0_number}; // @[Math.scala 450:32:@48148.4]
  assign _T_2040 = _GEN_15 << 2; // @[Math.scala 450:32:@48148.4]
  assign x708_rd_0_number = x524_lb_0_io_rPort_23_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 512:29:@47000.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 516:410:@47023.4]
  assign _GEN_16 = {{1'd0}, x708_rd_0_number}; // @[Math.scala 450:32:@48153.4]
  assign _T_2044 = _GEN_16 << 1; // @[Math.scala 450:32:@48153.4]
  assign x749_rd_0_number = x524_lb_0_io_rPort_16_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 607:29:@47316.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 611:410:@47339.4]
  assign _GEN_17 = {{1'd0}, x749_rd_0_number}; // @[Math.scala 450:32:@48158.4]
  assign _T_2048 = _GEN_17 << 1; // @[Math.scala 450:32:@48158.4]
  assign x858_sum_number = x858_sum_1_io_result; // @[Math.scala 154:22:@48247.4 Math.scala 155:14:@48248.4]
  assign _T_2084 = x858_sum_number[7:4]; // @[FixedPoint.scala 18:52:@48253.4]
  assign x721_rd_0_number = x524_lb_0_io_rPort_9_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 539:29:@47110.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 543:410:@47133.4]
  assign _GEN_18 = {{1'd0}, x721_rd_0_number}; // @[Math.scala 450:32:@48266.4]
  assign _T_2091 = _GEN_18 << 1; // @[Math.scala 450:32:@48266.4]
  assign _GEN_19 = {{2'd0}, x728_rd_0_number}; // @[Math.scala 450:32:@48271.4]
  assign _T_2095 = _GEN_19 << 2; // @[Math.scala 450:32:@48271.4]
  assign x776_rd_0_number = x524_lb_0_io_rPort_17_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 664:29:@47528.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 668:410:@47551.4]
  assign _GEN_20 = {{1'd0}, x776_rd_0_number}; // @[Math.scala 450:32:@48276.4]
  assign _T_2099 = _GEN_20 << 1; // @[Math.scala 450:32:@48276.4]
  assign x870_sum_number = x870_sum_1_io_result; // @[Math.scala 154:22:@48365.4 Math.scala 155:14:@48366.4]
  assign _T_2135 = x870_sum_number[7:4]; // @[FixedPoint.scala 18:52:@48371.4]
  assign _GEN_21 = {{2'd0}, x735_rd_0_number}; // @[Math.scala 450:32:@48384.4]
  assign _T_2142 = _GEN_21 << 2; // @[Math.scala 450:32:@48384.4]
  assign x783_rd_0_number = x524_lb_0_io_rPort_6_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 687:29:@47581.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 691:410:@47604.4]
  assign _GEN_22 = {{1'd0}, x783_rd_0_number}; // @[Math.scala 450:32:@48389.4]
  assign _T_2146 = _GEN_22 << 1; // @[Math.scala 450:32:@48389.4]
  assign x881_sum_number = x881_sum_1_io_result; // @[Math.scala 154:22:@48480.4 Math.scala 155:14:@48481.4]
  assign _T_2184 = x881_sum_number[7:4]; // @[FixedPoint.scala 18:52:@48486.4]
  assign _GEN_23 = {{2'd0}, x742_rd_0_number}; // @[Math.scala 450:32:@48499.4]
  assign _T_2191 = _GEN_23 << 2; // @[Math.scala 450:32:@48499.4]
  assign x790_rd_0_number = x524_lb_0_io_rPort_20_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 702:29:@47632.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 706:410:@47655.4]
  assign _GEN_24 = {{1'd0}, x790_rd_0_number}; // @[Math.scala 450:32:@48504.4]
  assign _T_2195 = _GEN_24 << 1; // @[Math.scala 450:32:@48504.4]
  assign x892_sum_number = x892_sum_1_io_result; // @[Math.scala 154:22:@48593.4 Math.scala 155:14:@48594.4]
  assign _T_2231 = x892_sum_number[7:4]; // @[FixedPoint.scala 18:52:@48599.4]
  assign _GEN_25 = {{2'd0}, x749_rd_0_number}; // @[Math.scala 450:32:@48612.4]
  assign _T_2238 = _GEN_25 << 2; // @[Math.scala 450:32:@48612.4]
  assign x756_rd_0_number = x524_lb_0_io_rPort_2_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 622:29:@47367.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 626:410:@47390.4]
  assign _GEN_26 = {{1'd0}, x756_rd_0_number}; // @[Math.scala 450:32:@48617.4]
  assign _T_2242 = _GEN_26 << 1; // @[Math.scala 450:32:@48617.4]
  assign x797_rd_0_number = x524_lb_0_io_rPort_1_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 717:29:@47683.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 721:410:@47706.4]
  assign _GEN_27 = {{1'd0}, x797_rd_0_number}; // @[Math.scala 450:32:@48622.4]
  assign _T_2246 = _GEN_27 << 1; // @[Math.scala 450:32:@48622.4]
  assign x904_sum_number = x904_sum_1_io_result; // @[Math.scala 154:22:@48711.4 Math.scala 155:14:@48712.4]
  assign _T_2282 = x904_sum_number[7:4]; // @[FixedPoint.scala 18:52:@48717.4]
  assign _T_2310 = RetimeWrapper_121_io_out; // @[package.scala 96:25:@48783.4 package.scala 96:25:@48784.4]
  assign _T_2312 = io_rr ? _T_2310 : 1'h0; // @[implicits.scala 55:10:@48785.4]
  assign _T_2313 = _T_368 & _T_2312; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 986:167:@48786.4]
  assign _T_2315 = _T_2313 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 986:255:@48788.4]
  assign _T_2316 = _T_2315 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 986:274:@48789.4]
  assign x1140_b522_D18 = RetimeWrapper_119_io_out; // @[package.scala 96:25:@48761.4 package.scala 96:25:@48762.4]
  assign _T_2317 = _T_2316 & x1140_b522_D18; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 986:300:@48790.4]
  assign x1137_b523_D18 = RetimeWrapper_116_io_out; // @[package.scala 96:25:@48734.4 package.scala 96:25:@48735.4]
  assign _T_2334 = RetimeWrapper_124_io_out; // @[package.scala 96:25:@48826.4 package.scala 96:25:@48827.4]
  assign _T_2336 = io_rr ? _T_2334 : 1'h0; // @[implicits.scala 55:10:@48828.4]
  assign _T_2337 = _T_368 & _T_2336; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 995:167:@48829.4]
  assign _T_2339 = _T_2337 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 995:255:@48831.4]
  assign _T_2340 = _T_2339 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 995:274:@48832.4]
  assign _T_2341 = _T_2340 & x1140_b522_D18; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 995:300:@48833.4]
  assign _T_2358 = RetimeWrapper_127_io_out; // @[package.scala 96:25:@48869.4 package.scala 96:25:@48870.4]
  assign _T_2360 = io_rr ? _T_2358 : 1'h0; // @[implicits.scala 55:10:@48871.4]
  assign _T_2361 = _T_368 & _T_2360; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1004:167:@48872.4]
  assign _T_2363 = _T_2361 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1004:255:@48874.4]
  assign _T_2364 = _T_2363 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1004:274:@48875.4]
  assign _T_2365 = _T_2364 & x1140_b522_D18; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1004:300:@48876.4]
  assign _T_2382 = RetimeWrapper_130_io_out; // @[package.scala 96:25:@48912.4 package.scala 96:25:@48913.4]
  assign _T_2384 = io_rr ? _T_2382 : 1'h0; // @[implicits.scala 55:10:@48914.4]
  assign _T_2385 = _T_368 & _T_2384; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1013:167:@48915.4]
  assign _T_2387 = _T_2385 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1013:255:@48917.4]
  assign _T_2388 = _T_2387 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1013:274:@48918.4]
  assign _T_2389 = _T_2388 & x1140_b522_D18; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1013:300:@48919.4]
  assign _T_2409 = RetimeWrapper_134_io_out; // @[package.scala 96:25:@48964.4 package.scala 96:25:@48965.4]
  assign _T_2411 = io_rr ? _T_2409 : 1'h0; // @[implicits.scala 55:10:@48966.4]
  assign _T_2412 = _T_368 & _T_2411; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1030:167:@48967.4]
  assign _T_2414 = _T_2412 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1030:255:@48969.4]
  assign _T_2415 = _T_2414 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1030:274:@48970.4]
  assign _T_2416 = _T_2415 & x1140_b522_D18; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1030:300:@48971.4]
  assign _T_2433 = RetimeWrapper_137_io_out; // @[package.scala 96:25:@49007.4 package.scala 96:25:@49008.4]
  assign _T_2435 = io_rr ? _T_2433 : 1'h0; // @[implicits.scala 55:10:@49009.4]
  assign _T_2436 = _T_368 & _T_2435; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1039:167:@49010.4]
  assign _T_2438 = _T_2436 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1039:255:@49012.4]
  assign _T_2439 = _T_2438 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1039:274:@49013.4]
  assign _T_2440 = _T_2439 & x1140_b522_D18; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1039:300:@49014.4]
  assign _T_2457 = RetimeWrapper_140_io_out; // @[package.scala 96:25:@49050.4 package.scala 96:25:@49051.4]
  assign _T_2459 = io_rr ? _T_2457 : 1'h0; // @[implicits.scala 55:10:@49052.4]
  assign _T_2460 = _T_368 & _T_2459; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1048:167:@49053.4]
  assign _T_2462 = _T_2460 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1048:255:@49055.4]
  assign _T_2463 = _T_2462 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1048:274:@49056.4]
  assign _T_2464 = _T_2463 & x1140_b522_D18; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1048:300:@49057.4]
  assign _T_2481 = RetimeWrapper_143_io_out; // @[package.scala 96:25:@49093.4 package.scala 96:25:@49094.4]
  assign _T_2483 = io_rr ? _T_2481 : 1'h0; // @[implicits.scala 55:10:@49095.4]
  assign _T_2484 = _T_368 & _T_2483; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1057:167:@49096.4]
  assign _T_2486 = _T_2484 & _T_368; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1057:255:@49098.4]
  assign _T_2487 = _T_2486 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1057:274:@49099.4]
  assign _T_2488 = _T_2487 & x1140_b522_D18; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1057:300:@49100.4]
  assign _T_2520 = RetimeWrapper_149_io_out; // @[package.scala 96:25:@49164.4 package.scala 96:25:@49165.4]
  assign _T_2522 = io_rr ? _T_2520 : 1'h0; // @[implicits.scala 55:10:@49166.4]
  assign _T_2523 = _T_368 & _T_2522; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1073:195:@49167.4]
  assign x1158_x606_D7 = RetimeWrapper_145_io_out; // @[package.scala 96:25:@49123.4 package.scala 96:25:@49124.4]
  assign _T_2524 = _T_2523 & x1158_x606_D7; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1073:283:@49168.4]
  assign x1159_b522_D19 = RetimeWrapper_146_io_out; // @[package.scala 96:25:@49132.4 package.scala 96:25:@49133.4]
  assign _T_2525 = _T_2524 & x1159_b522_D19; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1073:292:@49169.4]
  assign x1157_b523_D19 = RetimeWrapper_144_io_out; // @[package.scala 96:25:@49114.4 package.scala 96:25:@49115.4]
  assign _T_2549 = RetimeWrapper_152_io_out; // @[package.scala 96:25:@49208.4 package.scala 96:25:@49209.4]
  assign _T_2551 = io_rr ? _T_2549 : 1'h0; // @[implicits.scala 55:10:@49210.4]
  assign _T_2552 = _T_368 & _T_2551; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1084:195:@49211.4]
  assign x1163_x617_D7 = RetimeWrapper_151_io_out; // @[package.scala 96:25:@49194.4 package.scala 96:25:@49195.4]
  assign _T_2553 = _T_2552 & x1163_x617_D7; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1084:283:@49212.4]
  assign _T_2554 = _T_2553 & x1159_b522_D19; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1084:292:@49213.4]
  assign _T_2578 = RetimeWrapper_155_io_out; // @[package.scala 96:25:@49252.4 package.scala 96:25:@49253.4]
  assign _T_2580 = io_rr ? _T_2578 : 1'h0; // @[implicits.scala 55:10:@49254.4]
  assign _T_2581 = _T_368 & _T_2580; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1095:195:@49255.4]
  assign x1164_x625_D7 = RetimeWrapper_153_io_out; // @[package.scala 96:25:@49229.4 package.scala 96:25:@49230.4]
  assign _T_2582 = _T_2581 & x1164_x625_D7; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1095:283:@49256.4]
  assign _T_2583 = _T_2582 & x1159_b522_D19; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1095:292:@49257.4]
  assign _T_2607 = RetimeWrapper_158_io_out; // @[package.scala 96:25:@49296.4 package.scala 96:25:@49297.4]
  assign _T_2609 = io_rr ? _T_2607 : 1'h0; // @[implicits.scala 55:10:@49298.4]
  assign _T_2610 = _T_368 & _T_2609; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1106:195:@49299.4]
  assign x1167_x633_D7 = RetimeWrapper_157_io_out; // @[package.scala 96:25:@49282.4 package.scala 96:25:@49283.4]
  assign _T_2611 = _T_2610 & x1167_x633_D7; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1106:283:@49300.4]
  assign _T_2612 = _T_2611 & x1159_b522_D19; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1106:292:@49301.4]
  assign _T_2636 = RetimeWrapper_161_io_out; // @[package.scala 96:25:@49340.4 package.scala 96:25:@49341.4]
  assign _T_2638 = io_rr ? _T_2636 : 1'h0; // @[implicits.scala 55:10:@49342.4]
  assign _T_2639 = _T_368 & _T_2638; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1117:195:@49343.4]
  assign x1169_x642_D7 = RetimeWrapper_160_io_out; // @[package.scala 96:25:@49326.4 package.scala 96:25:@49327.4]
  assign _T_2640 = _T_2639 & x1169_x642_D7; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1117:283:@49344.4]
  assign _T_2641 = _T_2640 & x1159_b522_D19; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1117:292:@49345.4]
  assign _T_2668 = RetimeWrapper_165_io_out; // @[package.scala 96:25:@49393.4 package.scala 96:25:@49394.4]
  assign _T_2670 = io_rr ? _T_2668 : 1'h0; // @[implicits.scala 55:10:@49395.4]
  assign _T_2671 = _T_368 & _T_2670; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1130:195:@49396.4]
  assign x1170_x666_D7 = RetimeWrapper_162_io_out; // @[package.scala 96:25:@49361.4 package.scala 96:25:@49362.4]
  assign _T_2672 = _T_2671 & x1170_x666_D7; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1130:283:@49397.4]
  assign _T_2673 = _T_2672 & x1159_b522_D19; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1130:292:@49398.4]
  assign _T_2697 = RetimeWrapper_168_io_out; // @[package.scala 96:25:@49437.4 package.scala 96:25:@49438.4]
  assign _T_2699 = io_rr ? _T_2697 : 1'h0; // @[implicits.scala 55:10:@49439.4]
  assign _T_2700 = _T_368 & _T_2699; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1141:195:@49440.4]
  assign x1174_x676_D7 = RetimeWrapper_167_io_out; // @[package.scala 96:25:@49423.4 package.scala 96:25:@49424.4]
  assign _T_2701 = _T_2700 & x1174_x676_D7; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1141:283:@49441.4]
  assign _T_2702 = _T_2701 & x1159_b522_D19; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1141:292:@49442.4]
  assign _T_2726 = RetimeWrapper_171_io_out; // @[package.scala 96:25:@49481.4 package.scala 96:25:@49482.4]
  assign _T_2728 = io_rr ? _T_2726 : 1'h0; // @[implicits.scala 55:10:@49483.4]
  assign _T_2729 = _T_368 & _T_2728; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1152:195:@49484.4]
  assign x1175_x683_D7 = RetimeWrapper_169_io_out; // @[package.scala 96:25:@49458.4 package.scala 96:25:@49459.4]
  assign _T_2730 = _T_2729 & x1175_x683_D7; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1152:283:@49485.4]
  assign _T_2731 = _T_2730 & x1159_b522_D19; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1152:292:@49486.4]
  assign _T_2755 = RetimeWrapper_174_io_out; // @[package.scala 96:25:@49525.4 package.scala 96:25:@49526.4]
  assign _T_2757 = io_rr ? _T_2755 : 1'h0; // @[implicits.scala 55:10:@49527.4]
  assign _T_2758 = _T_368 & _T_2757; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1169:195:@49528.4]
  assign x1177_x690_D8 = RetimeWrapper_172_io_out; // @[package.scala 96:25:@49502.4 package.scala 96:25:@49503.4]
  assign _T_2759 = _T_2758 & x1177_x690_D8; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1169:283:@49529.4]
  assign _T_2760 = _T_2759 & x1159_b522_D19; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1169:292:@49530.4]
  assign _T_2784 = RetimeWrapper_177_io_out; // @[package.scala 96:25:@49569.4 package.scala 96:25:@49570.4]
  assign _T_2786 = io_rr ? _T_2784 : 1'h0; // @[implicits.scala 55:10:@49571.4]
  assign _T_2787 = _T_368 & _T_2786; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1180:195:@49572.4]
  assign x1180_x697_D7 = RetimeWrapper_176_io_out; // @[package.scala 96:25:@49555.4 package.scala 96:25:@49556.4]
  assign _T_2788 = _T_2787 & x1180_x697_D7; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1180:283:@49573.4]
  assign _T_2789 = _T_2788 & x1159_b522_D19; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1180:292:@49574.4]
  assign _T_2816 = RetimeWrapper_181_io_out; // @[package.scala 96:25:@49622.4 package.scala 96:25:@49623.4]
  assign _T_2818 = io_rr ? _T_2816 : 1'h0; // @[implicits.scala 55:10:@49624.4]
  assign _T_2819 = _T_368 & _T_2818; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1193:195:@49625.4]
  assign x1181_x714_D7 = RetimeWrapper_178_io_out; // @[package.scala 96:25:@49590.4 package.scala 96:25:@49591.4]
  assign _T_2820 = _T_2819 & x1181_x714_D7; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1193:283:@49626.4]
  assign _T_2821 = _T_2820 & x1159_b522_D19; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1193:292:@49627.4]
  assign _T_2845 = RetimeWrapper_184_io_out; // @[package.scala 96:25:@49666.4 package.scala 96:25:@49667.4]
  assign _T_2847 = io_rr ? _T_2845 : 1'h0; // @[implicits.scala 55:10:@49668.4]
  assign _T_2848 = _T_368 & _T_2847; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1204:195:@49669.4]
  assign x1184_x724_D7 = RetimeWrapper_182_io_out; // @[package.scala 96:25:@49643.4 package.scala 96:25:@49644.4]
  assign _T_2849 = _T_2848 & x1184_x724_D7; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1204:283:@49670.4]
  assign _T_2850 = _T_2849 & x1159_b522_D19; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1204:292:@49671.4]
  assign _T_2874 = RetimeWrapper_187_io_out; // @[package.scala 96:25:@49710.4 package.scala 96:25:@49711.4]
  assign _T_2876 = io_rr ? _T_2874 : 1'h0; // @[implicits.scala 55:10:@49712.4]
  assign _T_2877 = _T_368 & _T_2876; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1215:195:@49713.4]
  assign x1187_x731_D7 = RetimeWrapper_186_io_out; // @[package.scala 96:25:@49696.4 package.scala 96:25:@49697.4]
  assign _T_2878 = _T_2877 & x1187_x731_D7; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1215:283:@49714.4]
  assign _T_2879 = _T_2878 & x1159_b522_D19; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1215:292:@49715.4]
  assign _T_2903 = RetimeWrapper_190_io_out; // @[package.scala 96:25:@49754.4 package.scala 96:25:@49755.4]
  assign _T_2905 = io_rr ? _T_2903 : 1'h0; // @[implicits.scala 55:10:@49756.4]
  assign _T_2906 = _T_368 & _T_2905; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1226:195:@49757.4]
  assign x1188_x738_D7 = RetimeWrapper_188_io_out; // @[package.scala 96:25:@49731.4 package.scala 96:25:@49732.4]
  assign _T_2907 = _T_2906 & x1188_x738_D7; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1226:283:@49758.4]
  assign _T_2908 = _T_2907 & x1159_b522_D19; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1226:292:@49759.4]
  assign _T_2932 = RetimeWrapper_193_io_out; // @[package.scala 96:25:@49798.4 package.scala 96:25:@49799.4]
  assign _T_2934 = io_rr ? _T_2932 : 1'h0; // @[implicits.scala 55:10:@49800.4]
  assign _T_2935 = _T_368 & _T_2934; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1237:195:@49801.4]
  assign x1191_x745_D7 = RetimeWrapper_192_io_out; // @[package.scala 96:25:@49784.4 package.scala 96:25:@49785.4]
  assign _T_2936 = _T_2935 & x1191_x745_D7; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1237:283:@49802.4]
  assign _T_2937 = _T_2936 & x1159_b522_D19; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1237:292:@49803.4]
  assign x918_rd_0_number = x525_lb2_0_io_rPort_12_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1080:29:@49197.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1084:341:@49220.4]
  assign _GEN_28 = {{1'd0}, x918_rd_0_number}; // @[Math.scala 450:32:@49817.4]
  assign _T_2945 = _GEN_28 << 1; // @[Math.scala 450:32:@49817.4]
  assign x926_rd_0_number = x525_lb2_0_io_rPort_7_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1126:29:@49382.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1130:341:@49405.4]
  assign _GEN_29 = {{1'd0}, x926_rd_0_number}; // @[Math.scala 450:32:@49822.4]
  assign _T_2949 = _GEN_29 << 1; // @[Math.scala 450:32:@49822.4]
  assign x920_rd_0_number = x525_lb2_0_io_rPort_3_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1091:29:@49241.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1095:341:@49264.4]
  assign _GEN_30 = {{1'd0}, x920_rd_0_number}; // @[Math.scala 450:32:@49869.4]
  assign _T_2969 = _GEN_30 << 1; // @[Math.scala 450:32:@49869.4]
  assign x928_rd_0_number = x525_lb2_0_io_rPort_13_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1137:29:@49426.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1141:341:@49449.4]
  assign _GEN_31 = {{1'd0}, x928_rd_0_number}; // @[Math.scala 450:32:@49874.4]
  assign _T_2973 = _GEN_31 << 1; // @[Math.scala 450:32:@49874.4]
  assign x922_rd_0_number = x525_lb2_0_io_rPort_10_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1102:29:@49285.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1106:341:@49308.4]
  assign _GEN_32 = {{1'd0}, x922_rd_0_number}; // @[Math.scala 450:32:@49921.4]
  assign _T_2993 = _GEN_32 << 1; // @[Math.scala 450:32:@49921.4]
  assign x930_rd_0_number = x525_lb2_0_io_rPort_0_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1148:29:@49470.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1152:341:@49493.4]
  assign _GEN_33 = {{1'd0}, x930_rd_0_number}; // @[Math.scala 450:32:@49926.4]
  assign _T_2997 = _GEN_33 << 1; // @[Math.scala 450:32:@49926.4]
  assign x924_rd_0_number = x525_lb2_0_io_rPort_2_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1113:29:@49329.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1117:341:@49352.4]
  assign _GEN_34 = {{1'd0}, x924_rd_0_number}; // @[Math.scala 450:32:@49973.4]
  assign _T_3017 = _GEN_34 << 1; // @[Math.scala 450:32:@49973.4]
  assign x932_rd_0_number = x525_lb2_0_io_rPort_9_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1165:29:@49514.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1169:411:@49537.4]
  assign _GEN_35 = {{1'd0}, x932_rd_0_number}; // @[Math.scala 450:32:@49980.4]
  assign _T_3023 = _GEN_35 << 1; // @[Math.scala 450:32:@49980.4]
  assign x936_rd_0_number = x525_lb2_0_io_rPort_8_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1189:29:@49611.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1193:411:@49634.4]
  assign _GEN_36 = {{1'd0}, x936_rd_0_number}; // @[Math.scala 450:32:@50027.4]
  assign _T_3043 = _GEN_36 << 1; // @[Math.scala 450:32:@50027.4]
  assign x938_rd_0_number = x525_lb2_0_io_rPort_6_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1200:29:@49655.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1204:411:@49678.4]
  assign _GEN_37 = {{1'd0}, x938_rd_0_number}; // @[Math.scala 450:32:@50074.4]
  assign _T_3063 = _GEN_37 << 1; // @[Math.scala 450:32:@50074.4]
  assign x940_rd_0_number = x525_lb2_0_io_rPort_14_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1211:29:@49699.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1215:411:@49722.4]
  assign _GEN_38 = {{1'd0}, x940_rd_0_number}; // @[Math.scala 450:32:@50121.4]
  assign _T_3083 = _GEN_38 << 1; // @[Math.scala 450:32:@50121.4]
  assign x934_rd_0_number = x525_lb2_0_io_rPort_1_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1176:29:@49558.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1180:411:@49581.4]
  assign _GEN_39 = {{1'd0}, x934_rd_0_number}; // @[Math.scala 450:32:@50168.4]
  assign _T_3103 = _GEN_39 << 1; // @[Math.scala 450:32:@50168.4]
  assign x942_rd_0_number = x525_lb2_0_io_rPort_4_output_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1222:29:@49743.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 1226:411:@49766.4]
  assign _GEN_40 = {{1'd0}, x942_rd_0_number}; // @[Math.scala 450:32:@50173.4]
  assign _T_3107 = _GEN_40 << 1; // @[Math.scala 450:32:@50173.4]
  assign x984_div_number = x984_div_1_io_result; // @[Math.scala 331:22:@50163.4 Math.scala 332:14:@50164.4]
  assign x990_div_number = x990_div_1_io_result; // @[Math.scala 331:22:@50215.4 Math.scala 332:14:@50216.4]
  assign x974_div_number = x974_div_1_io_result; // @[Math.scala 331:22:@50069.4 Math.scala 332:14:@50070.4]
  assign x979_div_number = x979_div_1_io_result; // @[Math.scala 331:22:@50116.4 Math.scala 332:14:@50117.4]
  assign _T_3141 = {x974_div_number,x979_div_number,x984_div_number,x990_div_number}; // @[Cat.scala 30:58:@50230.4]
  assign x963_div_number = x963_div_1_io_result; // @[Math.scala 331:22:@49968.4 Math.scala 332:14:@49969.4]
  assign x969_div_number = x969_div_1_io_result; // @[Math.scala 331:22:@50022.4 Math.scala 332:14:@50023.4]
  assign x951_div_number = x951_div_1_io_result; // @[Math.scala 331:22:@49864.4 Math.scala 332:14:@49865.4]
  assign x957_div_number = x957_div_1_io_result; // @[Math.scala 331:22:@49916.4 Math.scala 332:14:@49917.4]
  assign _T_3144 = {x951_div_number,x957_div_number,x963_div_number,x969_div_number}; // @[Cat.scala 30:58:@50233.4]
  assign _T_3157 = RetimeWrapper_197_io_out; // @[package.scala 96:25:@50269.4 package.scala 96:25:@50270.4]
  assign _T_3159 = io_rr ? _T_3157 : 1'h0; // @[implicits.scala 55:10:@50271.4]
  assign x1192_b522_D29 = RetimeWrapper_195_io_out; // @[package.scala 96:25:@50251.4 package.scala 96:25:@50252.4]
  assign _T_3160 = _T_3159 & x1192_b522_D29; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1349:116:@50272.4]
  assign x1193_b523_D29 = RetimeWrapper_196_io_out; // @[package.scala 96:25:@50260.4 package.scala 96:25:@50261.4]
  assign _T_3161 = _T_3160 & x1193_b523_D29; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1349:123:@50273.4]
  assign x1063_x1051_D8_number = RetimeWrapper_2_io_out; // @[package.scala 96:25:@45468.4 package.scala 96:25:@45469.4]
  assign x1066_x539_sum_D7_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@45495.4 package.scala 96:25:@45496.4]
  assign x1069_x549_sum_D6_number = RetimeWrapper_9_io_out; // @[package.scala 96:25:@45580.4 package.scala 96:25:@45581.4]
  assign x1071_x558_sum_D6_number = RetimeWrapper_12_io_out; // @[package.scala 96:25:@45656.4 package.scala 96:25:@45657.4]
  assign x1072_x567_sum_D6_number = RetimeWrapper_14_io_out; // @[package.scala 96:25:@45723.4 package.scala 96:25:@45724.4]
  assign x1076_x1052_D7_number = RetimeWrapper_19_io_out; // @[package.scala 96:25:@45877.4 package.scala 96:25:@45878.4]
  assign x1077_x581_sum_D6_number = RetimeWrapper_20_io_out; // @[package.scala 96:25:@45886.4 package.scala 96:25:@45887.4]
  assign x1078_x587_sum_D6_number = RetimeWrapper_22_io_out; // @[package.scala 96:25:@45932.4 package.scala 96:25:@45933.4]
  assign x1081_x592_sum_D6_number = RetimeWrapper_26_io_out; // @[package.scala 96:25:@45996.4 package.scala 96:25:@45997.4]
  assign x1082_x597_sum_D6_number = RetimeWrapper_28_io_out; // @[package.scala 96:25:@46042.4 package.scala 96:25:@46043.4]
  assign x609_sum_number = x609_sum_1_io_result; // @[Math.scala 154:22:@46164.4 Math.scala 155:14:@46165.4]
  assign x1090_x1054_D1_number = RetimeWrapper_37_io_out; // @[package.scala 96:25:@46200.4 package.scala 96:25:@46201.4]
  assign x618_sum_number = x618_sum_1_io_result; // @[Math.scala 154:22:@46267.4 Math.scala 155:14:@46268.4]
  assign x626_sum_number = x626_sum_1_io_result; // @[Math.scala 154:22:@46345.4 Math.scala 155:14:@46346.4]
  assign x634_sum_number = x634_sum_1_io_result; // @[Math.scala 154:22:@46430.4 Math.scala 155:14:@46431.4]
  assign x645_sum_number = x645_sum_1_io_result; // @[Math.scala 154:22:@46509.4 Math.scala 155:14:@46510.4]
  assign x657_sum_number = x657_sum_1_io_result; // @[Math.scala 154:22:@46588.4 Math.scala 155:14:@46589.4]
  assign x669_sum_number = x669_sum_1_io_result; // @[Math.scala 154:22:@46706.4 Math.scala 155:14:@46707.4]
  assign x1107_x1056_D2_number = RetimeWrapper_60_io_out; // @[package.scala 96:25:@46724.4 package.scala 96:25:@46725.4]
  assign x677_sum_number = x677_sum_1_io_result; // @[Math.scala 154:22:@46766.4 Math.scala 155:14:@46767.4]
  assign x684_sum_number = x684_sum_1_io_result; // @[Math.scala 154:22:@46817.4 Math.scala 155:14:@46818.4]
  assign x1112_x691_sum_D1_number = RetimeWrapper_68_io_out; // @[package.scala 96:25:@46895.4 package.scala 96:25:@46896.4]
  assign x698_sum_number = x698_sum_1_io_result; // @[Math.scala 154:22:@46937.4 Math.scala 155:14:@46938.4]
  assign x705_sum_number = x705_sum_1_io_result; // @[Math.scala 154:22:@46988.4 Math.scala 155:14:@46989.4]
  assign x717_sum_number = x717_sum_1_io_result; // @[Math.scala 154:22:@47089.4 Math.scala 155:14:@47090.4]
  assign x1116_x1058_D1_number = RetimeWrapper_75_io_out; // @[package.scala 96:25:@47107.4 package.scala 96:25:@47108.4]
  assign x725_sum_number = x725_sum_1_io_result; // @[Math.scala 154:22:@47151.4 Math.scala 155:14:@47152.4]
  assign x732_sum_number = x732_sum_1_io_result; // @[Math.scala 154:22:@47202.4 Math.scala 155:14:@47203.4]
  assign x739_sum_number = x739_sum_1_io_result; // @[Math.scala 154:22:@47253.4 Math.scala 155:14:@47254.4]
  assign x746_sum_number = x746_sum_1_io_result; // @[Math.scala 154:22:@47304.4 Math.scala 155:14:@47305.4]
  assign x753_sum_number = x753_sum_1_io_result; // @[Math.scala 154:22:@47355.4 Math.scala 155:14:@47356.4]
  assign x765_sum_number = x765_sum_1_io_result; // @[Math.scala 154:22:@47456.4 Math.scala 155:14:@47457.4]
  assign x1123_x1060_D1_number = RetimeWrapper_88_io_out; // @[package.scala 96:25:@47474.4 package.scala 96:25:@47475.4]
  assign x773_sum_number = x773_sum_1_io_result; // @[Math.scala 154:22:@47516.4 Math.scala 155:14:@47517.4]
  assign x780_sum_number = x780_sum_1_io_result; // @[Math.scala 154:22:@47569.4 Math.scala 155:14:@47570.4]
  assign x787_sum_number = x787_sum_1_io_result; // @[Math.scala 154:22:@47620.4 Math.scala 155:14:@47621.4]
  assign x794_sum_number = x794_sum_1_io_result; // @[Math.scala 154:22:@47671.4 Math.scala 155:14:@47672.4]
  assign x801_sum_number = x801_sum_1_io_result; // @[Math.scala 154:22:@47722.4 Math.scala 155:14:@47723.4]
  assign x1138_x1051_D18_number = RetimeWrapper_117_io_out; // @[package.scala 96:25:@48743.4 package.scala 96:25:@48744.4]
  assign x1141_x539_sum_D17_number = RetimeWrapper_120_io_out; // @[package.scala 96:25:@48770.4 package.scala 96:25:@48771.4]
  assign x1143_x549_sum_D16_number = RetimeWrapper_123_io_out; // @[package.scala 96:25:@48813.4 package.scala 96:25:@48814.4]
  assign x1144_x558_sum_D16_number = RetimeWrapper_125_io_out; // @[package.scala 96:25:@48847.4 package.scala 96:25:@48848.4]
  assign x1146_x567_sum_D16_number = RetimeWrapper_128_io_out; // @[package.scala 96:25:@48890.4 package.scala 96:25:@48891.4]
  assign x1148_x1052_D17_number = RetimeWrapper_131_io_out; // @[package.scala 96:25:@48933.4 package.scala 96:25:@48934.4]
  assign x1150_x581_sum_D16_number = RetimeWrapper_133_io_out; // @[package.scala 96:25:@48951.4 package.scala 96:25:@48952.4]
  assign x1152_x587_sum_D16_number = RetimeWrapper_136_io_out; // @[package.scala 96:25:@48994.4 package.scala 96:25:@48995.4]
  assign x1154_x592_sum_D16_number = RetimeWrapper_139_io_out; // @[package.scala 96:25:@49037.4 package.scala 96:25:@49038.4]
  assign x1155_x597_sum_D16_number = RetimeWrapper_141_io_out; // @[package.scala 96:25:@49071.4 package.scala 96:25:@49072.4]
  assign x1160_x1054_D7_number = RetimeWrapper_147_io_out; // @[package.scala 96:25:@49141.4 package.scala 96:25:@49142.4]
  assign x1161_x609_sum_D6_number = RetimeWrapper_148_io_out; // @[package.scala 96:25:@49150.4 package.scala 96:25:@49151.4]
  assign x1162_x618_sum_D6_number = RetimeWrapper_150_io_out; // @[package.scala 96:25:@49185.4 package.scala 96:25:@49186.4]
  assign x1165_x626_sum_D6_number = RetimeWrapper_154_io_out; // @[package.scala 96:25:@49238.4 package.scala 96:25:@49239.4]
  assign x1166_x634_sum_D6_number = RetimeWrapper_156_io_out; // @[package.scala 96:25:@49273.4 package.scala 96:25:@49274.4]
  assign x1168_x645_sum_D6_number = RetimeWrapper_159_io_out; // @[package.scala 96:25:@49317.4 package.scala 96:25:@49318.4]
  assign x1171_x669_sum_D6_number = RetimeWrapper_163_io_out; // @[package.scala 96:25:@49370.4 package.scala 96:25:@49371.4]
  assign x1172_x1056_D8_number = RetimeWrapper_164_io_out; // @[package.scala 96:25:@49379.4 package.scala 96:25:@49380.4]
  assign x1173_x677_sum_D6_number = RetimeWrapper_166_io_out; // @[package.scala 96:25:@49414.4 package.scala 96:25:@49415.4]
  assign x1176_x684_sum_D6_number = RetimeWrapper_170_io_out; // @[package.scala 96:25:@49467.4 package.scala 96:25:@49468.4]
  assign x1178_x691_sum_D7_number = RetimeWrapper_173_io_out; // @[package.scala 96:25:@49511.4 package.scala 96:25:@49512.4]
  assign x1179_x698_sum_D6_number = RetimeWrapper_175_io_out; // @[package.scala 96:25:@49546.4 package.scala 96:25:@49547.4]
  assign x1182_x1058_D7_number = RetimeWrapper_179_io_out; // @[package.scala 96:25:@49599.4 package.scala 96:25:@49600.4]
  assign x1183_x717_sum_D6_number = RetimeWrapper_180_io_out; // @[package.scala 96:25:@49608.4 package.scala 96:25:@49609.4]
  assign x1185_x725_sum_D6_number = RetimeWrapper_183_io_out; // @[package.scala 96:25:@49652.4 package.scala 96:25:@49653.4]
  assign x1186_x732_sum_D6_number = RetimeWrapper_185_io_out; // @[package.scala 96:25:@49687.4 package.scala 96:25:@49688.4]
  assign x1189_x739_sum_D6_number = RetimeWrapper_189_io_out; // @[package.scala 96:25:@49740.4 package.scala 96:25:@49741.4]
  assign x1190_x746_sum_D6_number = RetimeWrapper_191_io_out; // @[package.scala 96:25:@49775.4 package.scala 96:25:@49776.4]
  assign io_in_x511_TREADY = _T_213 & _T_215; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 69:22:@45326.4 sm_x995_inr_Foreach_SAMPLER_BOX.scala 71:22:@45334.4]
  assign io_in_x512_TVALID = _T_3161 & io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1349:22:@50275.4]
  assign io_in_x512_TDATA = {{192'd0}, RetimeWrapper_194_io_out}; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1350:24:@50276.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@44932.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@44944.4]
  assign x524_lb_0_clock = clock; // @[:@44952.4]
  assign x524_lb_0_reset = reset; // @[:@44953.4]
  assign x524_lb_0_io_rPort_23_banks_0 = x1107_x1056_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@47018.4]
  assign x524_lb_0_io_rPort_23_ofs_0 = x705_sum_number[0]; // @[MemInterfaceType.scala 107:54:@47020.4]
  assign x524_lb_0_io_rPort_23_en_0 = _T_1351 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@47022.4]
  assign x524_lb_0_io_rPort_23_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@47021.4]
  assign x524_lb_0_io_rPort_22_banks_0 = x1116_x1058_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@47181.4]
  assign x524_lb_0_io_rPort_22_ofs_0 = x725_sum_number[0]; // @[MemInterfaceType.scala 107:54:@47183.4]
  assign x524_lb_0_io_rPort_22_en_0 = _T_1471 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@47185.4]
  assign x524_lb_0_io_rPort_22_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@47184.4]
  assign x524_lb_0_io_rPort_21_banks_0 = x1116_x1058_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@47232.4]
  assign x524_lb_0_io_rPort_21_ofs_0 = x732_sum_number[0]; // @[MemInterfaceType.scala 107:54:@47234.4]
  assign x524_lb_0_io_rPort_21_en_0 = _T_1504 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@47236.4]
  assign x524_lb_0_io_rPort_21_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@47235.4]
  assign x524_lb_0_io_rPort_20_banks_0 = x1123_x1060_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@47650.4]
  assign x524_lb_0_io_rPort_20_ofs_0 = x787_sum_number[0]; // @[MemInterfaceType.scala 107:54:@47652.4]
  assign x524_lb_0_io_rPort_20_en_0 = _T_1789 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@47654.4]
  assign x524_lb_0_io_rPort_20_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@47653.4]
  assign x524_lb_0_io_rPort_19_banks_0 = x1090_x1054_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@46221.4]
  assign x524_lb_0_io_rPort_19_ofs_0 = x609_sum_number[0]; // @[MemInterfaceType.scala 107:54:@46223.4]
  assign x524_lb_0_io_rPort_19_en_0 = _T_829 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@46225.4]
  assign x524_lb_0_io_rPort_19_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46224.4]
  assign x524_lb_0_io_rPort_18_banks_0 = x1107_x1056_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@46745.4]
  assign x524_lb_0_io_rPort_18_ofs_0 = x669_sum_number[0]; // @[MemInterfaceType.scala 107:54:@46747.4]
  assign x524_lb_0_io_rPort_18_en_0 = _T_1180 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@46749.4]
  assign x524_lb_0_io_rPort_18_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46748.4]
  assign x524_lb_0_io_rPort_17_banks_0 = x1123_x1060_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@47546.4]
  assign x524_lb_0_io_rPort_17_ofs_0 = x773_sum_number[0]; // @[MemInterfaceType.scala 107:54:@47548.4]
  assign x524_lb_0_io_rPort_17_en_0 = _T_1721 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@47550.4]
  assign x524_lb_0_io_rPort_17_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@47549.4]
  assign x524_lb_0_io_rPort_16_banks_0 = x1116_x1058_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@47334.4]
  assign x524_lb_0_io_rPort_16_ofs_0 = x746_sum_number[0]; // @[MemInterfaceType.scala 107:54:@47336.4]
  assign x524_lb_0_io_rPort_16_en_0 = _T_1570 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@47338.4]
  assign x524_lb_0_io_rPort_16_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@47337.4]
  assign x524_lb_0_io_rPort_15_banks_0 = x1107_x1056_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@46796.4]
  assign x524_lb_0_io_rPort_15_ofs_0 = x677_sum_number[0]; // @[MemInterfaceType.scala 107:54:@46798.4]
  assign x524_lb_0_io_rPort_15_en_0 = _T_1213 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@46800.4]
  assign x524_lb_0_io_rPort_15_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46799.4]
  assign x524_lb_0_io_rPort_14_banks_0 = x1123_x1060_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@47495.4]
  assign x524_lb_0_io_rPort_14_ofs_0 = x765_sum_number[0]; // @[MemInterfaceType.scala 107:54:@47497.4]
  assign x524_lb_0_io_rPort_14_en_0 = _T_1688 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@47499.4]
  assign x524_lb_0_io_rPort_14_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@47498.4]
  assign x524_lb_0_io_rPort_13_banks_0 = x1090_x1054_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@46297.4]
  assign x524_lb_0_io_rPort_13_ofs_0 = x618_sum_number[0]; // @[MemInterfaceType.scala 107:54:@46299.4]
  assign x524_lb_0_io_rPort_13_en_0 = _T_876 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@46301.4]
  assign x524_lb_0_io_rPort_13_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46300.4]
  assign x524_lb_0_io_rPort_12_banks_0 = x1090_x1054_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@46539.4]
  assign x524_lb_0_io_rPort_12_ofs_0 = x645_sum_number[0]; // @[MemInterfaceType.scala 107:54:@46541.4]
  assign x524_lb_0_io_rPort_12_en_0 = _T_1033 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@46543.4]
  assign x524_lb_0_io_rPort_12_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46542.4]
  assign x524_lb_0_io_rPort_11_banks_0 = x1123_x1060_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@47752.4]
  assign x524_lb_0_io_rPort_11_ofs_0 = x801_sum_number[0]; // @[MemInterfaceType.scala 107:54:@47754.4]
  assign x524_lb_0_io_rPort_11_en_0 = _T_1855 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@47756.4]
  assign x524_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@47755.4]
  assign x524_lb_0_io_rPort_10_banks_0 = x1107_x1056_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@46916.4]
  assign x524_lb_0_io_rPort_10_ofs_0 = x1112_x691_sum_D1_number[0]; // @[MemInterfaceType.scala 107:54:@46918.4]
  assign x524_lb_0_io_rPort_10_en_0 = _T_1285 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@46920.4]
  assign x524_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46919.4]
  assign x524_lb_0_io_rPort_9_banks_0 = x1116_x1058_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@47128.4]
  assign x524_lb_0_io_rPort_9_ofs_0 = x717_sum_number[0]; // @[MemInterfaceType.scala 107:54:@47130.4]
  assign x524_lb_0_io_rPort_9_en_0 = _T_1436 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@47132.4]
  assign x524_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@47131.4]
  assign x524_lb_0_io_rPort_8_banks_0 = x1107_x1056_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@46967.4]
  assign x524_lb_0_io_rPort_8_ofs_0 = x698_sum_number[0]; // @[MemInterfaceType.scala 107:54:@46969.4]
  assign x524_lb_0_io_rPort_8_en_0 = _T_1318 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@46971.4]
  assign x524_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46970.4]
  assign x524_lb_0_io_rPort_7_banks_0 = x1090_x1054_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@46460.4]
  assign x524_lb_0_io_rPort_7_ofs_0 = x634_sum_number[0]; // @[MemInterfaceType.scala 107:54:@46462.4]
  assign x524_lb_0_io_rPort_7_en_0 = _T_975 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@46464.4]
  assign x524_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46463.4]
  assign x524_lb_0_io_rPort_6_banks_0 = x1123_x1060_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@47599.4]
  assign x524_lb_0_io_rPort_6_ofs_0 = x780_sum_number[0]; // @[MemInterfaceType.scala 107:54:@47601.4]
  assign x524_lb_0_io_rPort_6_en_0 = _T_1756 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@47603.4]
  assign x524_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@47602.4]
  assign x524_lb_0_io_rPort_5_banks_0 = x1116_x1058_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@47283.4]
  assign x524_lb_0_io_rPort_5_ofs_0 = x739_sum_number[0]; // @[MemInterfaceType.scala 107:54:@47285.4]
  assign x524_lb_0_io_rPort_5_en_0 = _T_1537 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@47287.4]
  assign x524_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@47286.4]
  assign x524_lb_0_io_rPort_4_banks_0 = x1090_x1054_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@46618.4]
  assign x524_lb_0_io_rPort_4_ofs_0 = x657_sum_number[0]; // @[MemInterfaceType.scala 107:54:@46620.4]
  assign x524_lb_0_io_rPort_4_en_0 = _T_1091 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@46622.4]
  assign x524_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46621.4]
  assign x524_lb_0_io_rPort_3_banks_0 = x1107_x1056_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@46847.4]
  assign x524_lb_0_io_rPort_3_ofs_0 = x684_sum_number[0]; // @[MemInterfaceType.scala 107:54:@46849.4]
  assign x524_lb_0_io_rPort_3_en_0 = _T_1246 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@46851.4]
  assign x524_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46850.4]
  assign x524_lb_0_io_rPort_2_banks_0 = x1116_x1058_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@47385.4]
  assign x524_lb_0_io_rPort_2_ofs_0 = x753_sum_number[0]; // @[MemInterfaceType.scala 107:54:@47387.4]
  assign x524_lb_0_io_rPort_2_en_0 = _T_1603 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@47389.4]
  assign x524_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@47388.4]
  assign x524_lb_0_io_rPort_1_banks_0 = x1123_x1060_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@47701.4]
  assign x524_lb_0_io_rPort_1_ofs_0 = x794_sum_number[0]; // @[MemInterfaceType.scala 107:54:@47703.4]
  assign x524_lb_0_io_rPort_1_en_0 = _T_1822 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@47705.4]
  assign x524_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@47704.4]
  assign x524_lb_0_io_rPort_0_banks_0 = x1090_x1054_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@46375.4]
  assign x524_lb_0_io_rPort_0_ofs_0 = x626_sum_number[0]; // @[MemInterfaceType.scala 107:54:@46377.4]
  assign x524_lb_0_io_rPort_0_en_0 = _T_925 & x1087_b523_D13; // @[MemInterfaceType.scala 110:79:@46379.4]
  assign x524_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@46378.4]
  assign x524_lb_0_io_wPort_7_banks_0 = x1076_x1052_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@46018.4]
  assign x524_lb_0_io_wPort_7_ofs_0 = x1081_x592_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@46020.4]
  assign x524_lb_0_io_wPort_7_data_0 = RetimeWrapper_25_io_out; // @[MemInterfaceType.scala 90:56:@46021.4]
  assign x524_lb_0_io_wPort_7_en_0 = _T_701 & x1062_b523_D8; // @[MemInterfaceType.scala 93:57:@46023.4]
  assign x524_lb_0_io_wPort_6_banks_0 = x1063_x1051_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@45754.4]
  assign x524_lb_0_io_wPort_6_ofs_0 = x1072_x567_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@45756.4]
  assign x524_lb_0_io_wPort_6_data_0 = RetimeWrapper_15_io_out; // @[MemInterfaceType.scala 90:56:@45757.4]
  assign x524_lb_0_io_wPort_6_en_0 = _T_517 & x1062_b523_D8; // @[MemInterfaceType.scala 93:57:@45759.4]
  assign x524_lb_0_io_wPort_5_banks_0 = x1076_x1052_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@46073.4]
  assign x524_lb_0_io_wPort_5_ofs_0 = x1082_x597_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@46075.4]
  assign x524_lb_0_io_wPort_5_data_0 = RetimeWrapper_29_io_out; // @[MemInterfaceType.scala 90:56:@46076.4]
  assign x524_lb_0_io_wPort_5_en_0 = _T_729 & x1062_b523_D8; // @[MemInterfaceType.scala 93:57:@46078.4]
  assign x524_lb_0_io_wPort_4_banks_0 = x1063_x1051_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@45517.4]
  assign x524_lb_0_io_wPort_4_ofs_0 = x1066_x539_sum_D7_number[0]; // @[MemInterfaceType.scala 89:54:@45519.4]
  assign x524_lb_0_io_wPort_4_data_0 = RetimeWrapper_3_io_out; // @[MemInterfaceType.scala 90:56:@45520.4]
  assign x524_lb_0_io_wPort_4_en_0 = _T_379 & x1062_b523_D8; // @[MemInterfaceType.scala 93:57:@45522.4]
  assign x524_lb_0_io_wPort_3_banks_0 = x1076_x1052_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@45908.4]
  assign x524_lb_0_io_wPort_3_ofs_0 = x1077_x581_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@45910.4]
  assign x524_lb_0_io_wPort_3_data_0 = RetimeWrapper_18_io_out; // @[MemInterfaceType.scala 90:56:@45911.4]
  assign x524_lb_0_io_wPort_3_en_0 = _T_645 & x1062_b523_D8; // @[MemInterfaceType.scala 93:57:@45913.4]
  assign x524_lb_0_io_wPort_2_banks_0 = x1063_x1051_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@45602.4]
  assign x524_lb_0_io_wPort_2_ofs_0 = x1069_x549_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@45604.4]
  assign x524_lb_0_io_wPort_2_data_0 = RetimeWrapper_8_io_out; // @[MemInterfaceType.scala 90:56:@45605.4]
  assign x524_lb_0_io_wPort_2_en_0 = _T_427 & x1062_b523_D8; // @[MemInterfaceType.scala 93:57:@45607.4]
  assign x524_lb_0_io_wPort_1_banks_0 = x1063_x1051_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@45678.4]
  assign x524_lb_0_io_wPort_1_ofs_0 = x1071_x558_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@45680.4]
  assign x524_lb_0_io_wPort_1_data_0 = RetimeWrapper_11_io_out; // @[MemInterfaceType.scala 90:56:@45681.4]
  assign x524_lb_0_io_wPort_1_en_0 = _T_472 & x1062_b523_D8; // @[MemInterfaceType.scala 93:57:@45683.4]
  assign x524_lb_0_io_wPort_0_banks_0 = x1076_x1052_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@45963.4]
  assign x524_lb_0_io_wPort_0_ofs_0 = x1078_x587_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@45965.4]
  assign x524_lb_0_io_wPort_0_data_0 = RetimeWrapper_23_io_out; // @[MemInterfaceType.scala 90:56:@45966.4]
  assign x524_lb_0_io_wPort_0_en_0 = _T_673 & x1062_b523_D8; // @[MemInterfaceType.scala 93:57:@45968.4]
  assign x525_lb2_0_clock = clock; // @[:@45165.4]
  assign x525_lb2_0_reset = reset; // @[:@45166.4]
  assign x525_lb2_0_io_rPort_14_banks_0 = x1182_x1058_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@49717.4]
  assign x525_lb2_0_io_rPort_14_ofs_0 = x1186_x732_sum_D6_number[0]; // @[MemInterfaceType.scala 107:54:@49719.4]
  assign x525_lb2_0_io_rPort_14_en_0 = _T_2879 & x1157_b523_D19; // @[MemInterfaceType.scala 110:79:@49721.4]
  assign x525_lb2_0_io_rPort_14_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49720.4]
  assign x525_lb2_0_io_rPort_13_banks_0 = x1172_x1056_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@49444.4]
  assign x525_lb2_0_io_rPort_13_ofs_0 = x1173_x677_sum_D6_number[0]; // @[MemInterfaceType.scala 107:54:@49446.4]
  assign x525_lb2_0_io_rPort_13_en_0 = _T_2702 & x1157_b523_D19; // @[MemInterfaceType.scala 110:79:@49448.4]
  assign x525_lb2_0_io_rPort_13_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49447.4]
  assign x525_lb2_0_io_rPort_12_banks_0 = x1160_x1054_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@49215.4]
  assign x525_lb2_0_io_rPort_12_ofs_0 = x1162_x618_sum_D6_number[0]; // @[MemInterfaceType.scala 107:54:@49217.4]
  assign x525_lb2_0_io_rPort_12_en_0 = _T_2554 & x1157_b523_D19; // @[MemInterfaceType.scala 110:79:@49219.4]
  assign x525_lb2_0_io_rPort_12_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49218.4]
  assign x525_lb2_0_io_rPort_11_banks_0 = x1182_x1058_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@49805.4]
  assign x525_lb2_0_io_rPort_11_ofs_0 = x1190_x746_sum_D6_number[0]; // @[MemInterfaceType.scala 107:54:@49807.4]
  assign x525_lb2_0_io_rPort_11_en_0 = _T_2937 & x1157_b523_D19; // @[MemInterfaceType.scala 110:79:@49809.4]
  assign x525_lb2_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49808.4]
  assign x525_lb2_0_io_rPort_10_banks_0 = x1160_x1054_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@49303.4]
  assign x525_lb2_0_io_rPort_10_ofs_0 = x1166_x634_sum_D6_number[0]; // @[MemInterfaceType.scala 107:54:@49305.4]
  assign x525_lb2_0_io_rPort_10_en_0 = _T_2612 & x1157_b523_D19; // @[MemInterfaceType.scala 110:79:@49307.4]
  assign x525_lb2_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49306.4]
  assign x525_lb2_0_io_rPort_9_banks_0 = x1172_x1056_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@49532.4]
  assign x525_lb2_0_io_rPort_9_ofs_0 = x1178_x691_sum_D7_number[0]; // @[MemInterfaceType.scala 107:54:@49534.4]
  assign x525_lb2_0_io_rPort_9_en_0 = _T_2760 & x1157_b523_D19; // @[MemInterfaceType.scala 110:79:@49536.4]
  assign x525_lb2_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49535.4]
  assign x525_lb2_0_io_rPort_8_banks_0 = x1182_x1058_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@49629.4]
  assign x525_lb2_0_io_rPort_8_ofs_0 = x1183_x717_sum_D6_number[0]; // @[MemInterfaceType.scala 107:54:@49631.4]
  assign x525_lb2_0_io_rPort_8_en_0 = _T_2821 & x1157_b523_D19; // @[MemInterfaceType.scala 110:79:@49633.4]
  assign x525_lb2_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49632.4]
  assign x525_lb2_0_io_rPort_7_banks_0 = x1172_x1056_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@49400.4]
  assign x525_lb2_0_io_rPort_7_ofs_0 = x1171_x669_sum_D6_number[0]; // @[MemInterfaceType.scala 107:54:@49402.4]
  assign x525_lb2_0_io_rPort_7_en_0 = _T_2673 & x1157_b523_D19; // @[MemInterfaceType.scala 110:79:@49404.4]
  assign x525_lb2_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49403.4]
  assign x525_lb2_0_io_rPort_6_banks_0 = x1182_x1058_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@49673.4]
  assign x525_lb2_0_io_rPort_6_ofs_0 = x1185_x725_sum_D6_number[0]; // @[MemInterfaceType.scala 107:54:@49675.4]
  assign x525_lb2_0_io_rPort_6_en_0 = _T_2850 & x1157_b523_D19; // @[MemInterfaceType.scala 110:79:@49677.4]
  assign x525_lb2_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49676.4]
  assign x525_lb2_0_io_rPort_5_banks_0 = x1160_x1054_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@49171.4]
  assign x525_lb2_0_io_rPort_5_ofs_0 = x1161_x609_sum_D6_number[0]; // @[MemInterfaceType.scala 107:54:@49173.4]
  assign x525_lb2_0_io_rPort_5_en_0 = _T_2525 & x1157_b523_D19; // @[MemInterfaceType.scala 110:79:@49175.4]
  assign x525_lb2_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49174.4]
  assign x525_lb2_0_io_rPort_4_banks_0 = x1182_x1058_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@49761.4]
  assign x525_lb2_0_io_rPort_4_ofs_0 = x1189_x739_sum_D6_number[0]; // @[MemInterfaceType.scala 107:54:@49763.4]
  assign x525_lb2_0_io_rPort_4_en_0 = _T_2908 & x1157_b523_D19; // @[MemInterfaceType.scala 110:79:@49765.4]
  assign x525_lb2_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49764.4]
  assign x525_lb2_0_io_rPort_3_banks_0 = x1160_x1054_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@49259.4]
  assign x525_lb2_0_io_rPort_3_ofs_0 = x1165_x626_sum_D6_number[0]; // @[MemInterfaceType.scala 107:54:@49261.4]
  assign x525_lb2_0_io_rPort_3_en_0 = _T_2583 & x1157_b523_D19; // @[MemInterfaceType.scala 110:79:@49263.4]
  assign x525_lb2_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49262.4]
  assign x525_lb2_0_io_rPort_2_banks_0 = x1160_x1054_D7_number[2:0]; // @[MemInterfaceType.scala 106:58:@49347.4]
  assign x525_lb2_0_io_rPort_2_ofs_0 = x1168_x645_sum_D6_number[0]; // @[MemInterfaceType.scala 107:54:@49349.4]
  assign x525_lb2_0_io_rPort_2_en_0 = _T_2641 & x1157_b523_D19; // @[MemInterfaceType.scala 110:79:@49351.4]
  assign x525_lb2_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49350.4]
  assign x525_lb2_0_io_rPort_1_banks_0 = x1172_x1056_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@49576.4]
  assign x525_lb2_0_io_rPort_1_ofs_0 = x1179_x698_sum_D6_number[0]; // @[MemInterfaceType.scala 107:54:@49578.4]
  assign x525_lb2_0_io_rPort_1_en_0 = _T_2789 & x1157_b523_D19; // @[MemInterfaceType.scala 110:79:@49580.4]
  assign x525_lb2_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49579.4]
  assign x525_lb2_0_io_rPort_0_banks_0 = x1172_x1056_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@49488.4]
  assign x525_lb2_0_io_rPort_0_ofs_0 = x1176_x684_sum_D6_number[0]; // @[MemInterfaceType.scala 107:54:@49490.4]
  assign x525_lb2_0_io_rPort_0_en_0 = _T_2731 & x1157_b523_D19; // @[MemInterfaceType.scala 110:79:@49492.4]
  assign x525_lb2_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@49491.4]
  assign x525_lb2_0_io_wPort_7_banks_0 = x1138_x1051_D18_number[2:0]; // @[MemInterfaceType.scala 88:58:@48835.4]
  assign x525_lb2_0_io_wPort_7_ofs_0 = x1143_x549_sum_D16_number[0]; // @[MemInterfaceType.scala 89:54:@48837.4]
  assign x525_lb2_0_io_wPort_7_data_0 = RetimeWrapper_122_io_out; // @[MemInterfaceType.scala 90:56:@48838.4]
  assign x525_lb2_0_io_wPort_7_en_0 = _T_2341 & x1137_b523_D18; // @[MemInterfaceType.scala 93:57:@48840.4]
  assign x525_lb2_0_io_wPort_6_banks_0 = x1148_x1052_D17_number[2:0]; // @[MemInterfaceType.scala 88:58:@49102.4]
  assign x525_lb2_0_io_wPort_6_ofs_0 = x1155_x597_sum_D16_number[0]; // @[MemInterfaceType.scala 89:54:@49104.4]
  assign x525_lb2_0_io_wPort_6_data_0 = RetimeWrapper_142_io_out; // @[MemInterfaceType.scala 90:56:@49105.4]
  assign x525_lb2_0_io_wPort_6_en_0 = _T_2488 & x1137_b523_D18; // @[MemInterfaceType.scala 93:57:@49107.4]
  assign x525_lb2_0_io_wPort_5_banks_0 = x1138_x1051_D18_number[2:0]; // @[MemInterfaceType.scala 88:58:@48792.4]
  assign x525_lb2_0_io_wPort_5_ofs_0 = x1141_x539_sum_D17_number[0]; // @[MemInterfaceType.scala 89:54:@48794.4]
  assign x525_lb2_0_io_wPort_5_data_0 = RetimeWrapper_118_io_out; // @[MemInterfaceType.scala 90:56:@48795.4]
  assign x525_lb2_0_io_wPort_5_en_0 = _T_2317 & x1137_b523_D18; // @[MemInterfaceType.scala 93:57:@48797.4]
  assign x525_lb2_0_io_wPort_4_banks_0 = x1148_x1052_D17_number[2:0]; // @[MemInterfaceType.scala 88:58:@49016.4]
  assign x525_lb2_0_io_wPort_4_ofs_0 = x1152_x587_sum_D16_number[0]; // @[MemInterfaceType.scala 89:54:@49018.4]
  assign x525_lb2_0_io_wPort_4_data_0 = RetimeWrapper_135_io_out; // @[MemInterfaceType.scala 90:56:@49019.4]
  assign x525_lb2_0_io_wPort_4_en_0 = _T_2440 & x1137_b523_D18; // @[MemInterfaceType.scala 93:57:@49021.4]
  assign x525_lb2_0_io_wPort_3_banks_0 = x1148_x1052_D17_number[2:0]; // @[MemInterfaceType.scala 88:58:@48973.4]
  assign x525_lb2_0_io_wPort_3_ofs_0 = x1150_x581_sum_D16_number[0]; // @[MemInterfaceType.scala 89:54:@48975.4]
  assign x525_lb2_0_io_wPort_3_data_0 = RetimeWrapper_132_io_out; // @[MemInterfaceType.scala 90:56:@48976.4]
  assign x525_lb2_0_io_wPort_3_en_0 = _T_2416 & x1137_b523_D18; // @[MemInterfaceType.scala 93:57:@48978.4]
  assign x525_lb2_0_io_wPort_2_banks_0 = x1138_x1051_D18_number[2:0]; // @[MemInterfaceType.scala 88:58:@48921.4]
  assign x525_lb2_0_io_wPort_2_ofs_0 = x1146_x567_sum_D16_number[0]; // @[MemInterfaceType.scala 89:54:@48923.4]
  assign x525_lb2_0_io_wPort_2_data_0 = RetimeWrapper_129_io_out; // @[MemInterfaceType.scala 90:56:@48924.4]
  assign x525_lb2_0_io_wPort_2_en_0 = _T_2389 & x1137_b523_D18; // @[MemInterfaceType.scala 93:57:@48926.4]
  assign x525_lb2_0_io_wPort_1_banks_0 = x1148_x1052_D17_number[2:0]; // @[MemInterfaceType.scala 88:58:@49059.4]
  assign x525_lb2_0_io_wPort_1_ofs_0 = x1154_x592_sum_D16_number[0]; // @[MemInterfaceType.scala 89:54:@49061.4]
  assign x525_lb2_0_io_wPort_1_data_0 = RetimeWrapper_138_io_out; // @[MemInterfaceType.scala 90:56:@49062.4]
  assign x525_lb2_0_io_wPort_1_en_0 = _T_2464 & x1137_b523_D18; // @[MemInterfaceType.scala 93:57:@49064.4]
  assign x525_lb2_0_io_wPort_0_banks_0 = x1138_x1051_D18_number[2:0]; // @[MemInterfaceType.scala 88:58:@48878.4]
  assign x525_lb2_0_io_wPort_0_ofs_0 = x1144_x558_sum_D16_number[0]; // @[MemInterfaceType.scala 89:54:@48880.4]
  assign x525_lb2_0_io_wPort_0_data_0 = RetimeWrapper_126_io_out; // @[MemInterfaceType.scala 90:56:@48881.4]
  assign x525_lb2_0_io_wPort_0_en_0 = _T_2365 & x1137_b523_D18; // @[MemInterfaceType.scala 93:57:@48883.4]
  assign RetimeWrapper_clock = clock; // @[:@45337.4]
  assign RetimeWrapper_reset = reset; // @[:@45338.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45340.4]
  assign RetimeWrapper_io_in = io_in_x511_TDATA[63:0]; // @[package.scala 94:16:@45339.4]
  assign x539_sum_1_clock = clock; // @[:@45445.4]
  assign x539_sum_1_reset = reset; // @[:@45446.4]
  assign x539_sum_1_io_a = {_T_332,_T_333}; // @[Math.scala 151:17:@45447.4]
  assign x539_sum_1_io_b = {_T_342,_T_343}; // @[Math.scala 152:17:@45448.4]
  assign x539_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@45449.4]
  assign RetimeWrapper_1_clock = clock; // @[:@45455.4]
  assign RetimeWrapper_1_reset = reset; // @[:@45456.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45458.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@45457.4]
  assign RetimeWrapper_2_clock = clock; // @[:@45464.4]
  assign RetimeWrapper_2_reset = reset; // @[:@45465.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45467.4]
  assign RetimeWrapper_2_io_in = $unsigned(_T_323); // @[package.scala 94:16:@45466.4]
  assign RetimeWrapper_3_clock = clock; // @[:@45473.4]
  assign RetimeWrapper_3_reset = reset; // @[:@45474.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45476.4]
  assign RetimeWrapper_3_io_in = x1061_x526_D1_0_number[7:0]; // @[package.scala 94:16:@45475.4]
  assign RetimeWrapper_4_clock = clock; // @[:@45482.4]
  assign RetimeWrapper_4_reset = reset; // @[:@45483.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45485.4]
  assign RetimeWrapper_4_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@45484.4]
  assign RetimeWrapper_5_clock = clock; // @[:@45491.4]
  assign RetimeWrapper_5_reset = reset; // @[:@45492.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45494.4]
  assign RetimeWrapper_5_io_in = x539_sum_1_io_result; // @[package.scala 94:16:@45493.4]
  assign RetimeWrapper_6_clock = clock; // @[:@45504.4]
  assign RetimeWrapper_6_reset = reset; // @[:@45505.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45507.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45506.4]
  assign x545_rdcol_1_clock = clock; // @[:@45527.4]
  assign x545_rdcol_1_reset = reset; // @[:@45528.4]
  assign x545_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@45529.4]
  assign x545_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@45530.4]
  assign x545_rdcol_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@45531.4]
  assign RetimeWrapper_7_clock = clock; // @[:@45548.4]
  assign RetimeWrapper_7_reset = reset; // @[:@45549.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45551.4]
  assign RetimeWrapper_7_io_in = {_T_332,_T_333}; // @[package.scala 94:16:@45550.4]
  assign x549_sum_1_clock = clock; // @[:@45557.4]
  assign x549_sum_1_reset = reset; // @[:@45558.4]
  assign x549_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@45559.4]
  assign x549_sum_1_io_b = {_T_396,_T_397}; // @[Math.scala 152:17:@45560.4]
  assign x549_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@45561.4]
  assign RetimeWrapper_8_clock = clock; // @[:@45567.4]
  assign RetimeWrapper_8_reset = reset; // @[:@45568.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45570.4]
  assign RetimeWrapper_8_io_in = x1061_x526_D1_0_number[15:8]; // @[package.scala 94:16:@45569.4]
  assign RetimeWrapper_9_clock = clock; // @[:@45576.4]
  assign RetimeWrapper_9_reset = reset; // @[:@45577.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45579.4]
  assign RetimeWrapper_9_io_in = x549_sum_1_io_result; // @[package.scala 94:16:@45578.4]
  assign RetimeWrapper_10_clock = clock; // @[:@45589.4]
  assign RetimeWrapper_10_reset = reset; // @[:@45590.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45592.4]
  assign RetimeWrapper_10_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45591.4]
  assign x554_rdcol_1_clock = clock; // @[:@45612.4]
  assign x554_rdcol_1_reset = reset; // @[:@45613.4]
  assign x554_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@45614.4]
  assign x554_rdcol_1_io_b = 32'h2; // @[Math.scala 152:17:@45615.4]
  assign x554_rdcol_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@45616.4]
  assign x558_sum_1_clock = clock; // @[:@45633.4]
  assign x558_sum_1_reset = reset; // @[:@45634.4]
  assign x558_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@45635.4]
  assign x558_sum_1_io_b = {_T_444,_T_445}; // @[Math.scala 152:17:@45636.4]
  assign x558_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@45637.4]
  assign RetimeWrapper_11_clock = clock; // @[:@45643.4]
  assign RetimeWrapper_11_reset = reset; // @[:@45644.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45646.4]
  assign RetimeWrapper_11_io_in = x1061_x526_D1_0_number[23:16]; // @[package.scala 94:16:@45645.4]
  assign RetimeWrapper_12_clock = clock; // @[:@45652.4]
  assign RetimeWrapper_12_reset = reset; // @[:@45653.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45655.4]
  assign RetimeWrapper_12_io_in = x558_sum_1_io_result; // @[package.scala 94:16:@45654.4]
  assign RetimeWrapper_13_clock = clock; // @[:@45665.4]
  assign RetimeWrapper_13_reset = reset; // @[:@45666.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45668.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45667.4]
  assign x563_rdcol_1_clock = clock; // @[:@45688.4]
  assign x563_rdcol_1_reset = reset; // @[:@45689.4]
  assign x563_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@45690.4]
  assign x563_rdcol_1_io_b = 32'h3; // @[Math.scala 152:17:@45691.4]
  assign x563_rdcol_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@45692.4]
  assign x567_sum_1_clock = clock; // @[:@45709.4]
  assign x567_sum_1_reset = reset; // @[:@45710.4]
  assign x567_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@45711.4]
  assign x567_sum_1_io_b = {_T_489,_T_490}; // @[Math.scala 152:17:@45712.4]
  assign x567_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@45713.4]
  assign RetimeWrapper_14_clock = clock; // @[:@45719.4]
  assign RetimeWrapper_14_reset = reset; // @[:@45720.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45722.4]
  assign RetimeWrapper_14_io_in = x567_sum_1_io_result; // @[package.scala 94:16:@45721.4]
  assign RetimeWrapper_15_clock = clock; // @[:@45728.4]
  assign RetimeWrapper_15_reset = reset; // @[:@45729.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45731.4]
  assign RetimeWrapper_15_io_in = x1061_x526_D1_0_number[31:24]; // @[package.scala 94:16:@45730.4]
  assign RetimeWrapper_16_clock = clock; // @[:@45741.4]
  assign RetimeWrapper_16_reset = reset; // @[:@45742.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45744.4]
  assign RetimeWrapper_16_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45743.4]
  assign x572_rdrow_1_clock = clock; // @[:@45764.4]
  assign x572_rdrow_1_reset = reset; // @[:@45765.4]
  assign x572_rdrow_1_io_a = __io_result; // @[Math.scala 151:17:@45766.4]
  assign x572_rdrow_1_io_b = 32'h1; // @[Math.scala 152:17:@45767.4]
  assign x572_rdrow_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@45768.4]
  assign RetimeWrapper_17_clock = clock; // @[:@45845.4]
  assign RetimeWrapper_17_reset = reset; // @[:@45846.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45848.4]
  assign RetimeWrapper_17_io_in = {_T_342,_T_343}; // @[package.scala 94:16:@45847.4]
  assign x581_sum_1_clock = clock; // @[:@45854.4]
  assign x581_sum_1_reset = reset; // @[:@45855.4]
  assign x581_sum_1_io_a = {_T_611,_T_612}; // @[Math.scala 151:17:@45856.4]
  assign x581_sum_1_io_b = RetimeWrapper_17_io_out; // @[Math.scala 152:17:@45857.4]
  assign x581_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@45858.4]
  assign RetimeWrapper_18_clock = clock; // @[:@45864.4]
  assign RetimeWrapper_18_reset = reset; // @[:@45865.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45867.4]
  assign RetimeWrapper_18_io_in = x1061_x526_D1_0_number[39:32]; // @[package.scala 94:16:@45866.4]
  assign RetimeWrapper_19_clock = clock; // @[:@45873.4]
  assign RetimeWrapper_19_reset = reset; // @[:@45874.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45876.4]
  assign RetimeWrapper_19_io_in = $unsigned(_T_602); // @[package.scala 94:16:@45875.4]
  assign RetimeWrapper_20_clock = clock; // @[:@45882.4]
  assign RetimeWrapper_20_reset = reset; // @[:@45883.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45885.4]
  assign RetimeWrapper_20_io_in = x581_sum_1_io_result; // @[package.scala 94:16:@45884.4]
  assign RetimeWrapper_21_clock = clock; // @[:@45895.4]
  assign RetimeWrapper_21_reset = reset; // @[:@45896.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45898.4]
  assign RetimeWrapper_21_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45897.4]
  assign x587_sum_1_clock = clock; // @[:@45918.4]
  assign x587_sum_1_reset = reset; // @[:@45919.4]
  assign x587_sum_1_io_a = {_T_611,_T_612}; // @[Math.scala 151:17:@45920.4]
  assign x587_sum_1_io_b = {_T_396,_T_397}; // @[Math.scala 152:17:@45921.4]
  assign x587_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@45922.4]
  assign RetimeWrapper_22_clock = clock; // @[:@45928.4]
  assign RetimeWrapper_22_reset = reset; // @[:@45929.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45931.4]
  assign RetimeWrapper_22_io_in = x587_sum_1_io_result; // @[package.scala 94:16:@45930.4]
  assign RetimeWrapper_23_clock = clock; // @[:@45937.4]
  assign RetimeWrapper_23_reset = reset; // @[:@45938.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45940.4]
  assign RetimeWrapper_23_io_in = x1061_x526_D1_0_number[47:40]; // @[package.scala 94:16:@45939.4]
  assign RetimeWrapper_24_clock = clock; // @[:@45950.4]
  assign RetimeWrapper_24_reset = reset; // @[:@45951.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45953.4]
  assign RetimeWrapper_24_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45952.4]
  assign x592_sum_1_clock = clock; // @[:@45973.4]
  assign x592_sum_1_reset = reset; // @[:@45974.4]
  assign x592_sum_1_io_a = {_T_611,_T_612}; // @[Math.scala 151:17:@45975.4]
  assign x592_sum_1_io_b = {_T_444,_T_445}; // @[Math.scala 152:17:@45976.4]
  assign x592_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@45977.4]
  assign RetimeWrapper_25_clock = clock; // @[:@45983.4]
  assign RetimeWrapper_25_reset = reset; // @[:@45984.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45986.4]
  assign RetimeWrapper_25_io_in = x1061_x526_D1_0_number[55:48]; // @[package.scala 94:16:@45985.4]
  assign RetimeWrapper_26_clock = clock; // @[:@45992.4]
  assign RetimeWrapper_26_reset = reset; // @[:@45993.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@45995.4]
  assign RetimeWrapper_26_io_in = x592_sum_1_io_result; // @[package.scala 94:16:@45994.4]
  assign RetimeWrapper_27_clock = clock; // @[:@46005.4]
  assign RetimeWrapper_27_reset = reset; // @[:@46006.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46008.4]
  assign RetimeWrapper_27_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46007.4]
  assign x597_sum_1_clock = clock; // @[:@46028.4]
  assign x597_sum_1_reset = reset; // @[:@46029.4]
  assign x597_sum_1_io_a = {_T_611,_T_612}; // @[Math.scala 151:17:@46030.4]
  assign x597_sum_1_io_b = {_T_489,_T_490}; // @[Math.scala 152:17:@46031.4]
  assign x597_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@46032.4]
  assign RetimeWrapper_28_clock = clock; // @[:@46038.4]
  assign RetimeWrapper_28_reset = reset; // @[:@46039.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46041.4]
  assign RetimeWrapper_28_io_in = x597_sum_1_io_result; // @[package.scala 94:16:@46040.4]
  assign RetimeWrapper_29_clock = clock; // @[:@46047.4]
  assign RetimeWrapper_29_reset = reset; // @[:@46048.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46050.4]
  assign RetimeWrapper_29_io_in = x1061_x526_D1_0_number[63:56]; // @[package.scala 94:16:@46049.4]
  assign RetimeWrapper_30_clock = clock; // @[:@46060.4]
  assign RetimeWrapper_30_reset = reset; // @[:@46061.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46063.4]
  assign RetimeWrapper_30_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46062.4]
  assign RetimeWrapper_31_clock = clock; // @[:@46081.4]
  assign RetimeWrapper_31_reset = reset; // @[:@46082.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46084.4]
  assign RetimeWrapper_31_io_in = x572_rdrow_1_io_result; // @[package.scala 94:16:@46083.4]
  assign RetimeWrapper_32_clock = clock; // @[:@46108.4]
  assign RetimeWrapper_32_reset = reset; // @[:@46109.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46111.4]
  assign RetimeWrapper_32_io_in = x563_rdcol_1_io_result; // @[package.scala 94:16:@46110.4]
  assign RetimeWrapper_33_clock = clock; // @[:@46150.4]
  assign RetimeWrapper_33_reset = reset; // @[:@46151.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46153.4]
  assign RetimeWrapper_33_io_in = {_T_489,_T_490}; // @[package.scala 94:16:@46152.4]
  assign x609_sum_1_clock = clock; // @[:@46159.4]
  assign x609_sum_1_reset = reset; // @[:@46160.4]
  assign x609_sum_1_io_a = {_T_788,_T_789}; // @[Math.scala 151:17:@46161.4]
  assign x609_sum_1_io_b = RetimeWrapper_33_io_out; // @[Math.scala 152:17:@46162.4]
  assign x609_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@46163.4]
  assign RetimeWrapper_34_clock = clock; // @[:@46169.4]
  assign RetimeWrapper_34_reset = reset; // @[:@46170.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46172.4]
  assign RetimeWrapper_34_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@46171.4]
  assign RetimeWrapper_35_clock = clock; // @[:@46178.4]
  assign RetimeWrapper_35_reset = reset; // @[:@46179.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46181.4]
  assign RetimeWrapper_35_io_in = ~ x605; // @[package.scala 94:16:@46180.4]
  assign RetimeWrapper_36_clock = clock; // @[:@46187.4]
  assign RetimeWrapper_36_reset = reset; // @[:@46188.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46190.4]
  assign RetimeWrapper_36_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@46189.4]
  assign RetimeWrapper_37_clock = clock; // @[:@46196.4]
  assign RetimeWrapper_37_reset = reset; // @[:@46197.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46199.4]
  assign RetimeWrapper_37_io_in = $unsigned(_T_779); // @[package.scala 94:16:@46198.4]
  assign RetimeWrapper_38_clock = clock; // @[:@46210.4]
  assign RetimeWrapper_38_reset = reset; // @[:@46211.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46213.4]
  assign RetimeWrapper_38_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46212.4]
  assign RetimeWrapper_39_clock = clock; // @[:@46231.4]
  assign RetimeWrapper_39_reset = reset; // @[:@46232.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46234.4]
  assign RetimeWrapper_39_io_in = x554_rdcol_1_io_result; // @[package.scala 94:16:@46233.4]
  assign RetimeWrapper_40_clock = clock; // @[:@46253.4]
  assign RetimeWrapper_40_reset = reset; // @[:@46254.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46256.4]
  assign RetimeWrapper_40_io_in = {_T_444,_T_445}; // @[package.scala 94:16:@46255.4]
  assign x618_sum_1_clock = clock; // @[:@46262.4]
  assign x618_sum_1_reset = reset; // @[:@46263.4]
  assign x618_sum_1_io_a = {_T_788,_T_789}; // @[Math.scala 151:17:@46264.4]
  assign x618_sum_1_io_b = RetimeWrapper_40_io_out; // @[Math.scala 152:17:@46265.4]
  assign x618_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@46266.4]
  assign RetimeWrapper_41_clock = clock; // @[:@46272.4]
  assign RetimeWrapper_41_reset = reset; // @[:@46273.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46275.4]
  assign RetimeWrapper_41_io_in = ~ x616; // @[package.scala 94:16:@46274.4]
  assign RetimeWrapper_42_clock = clock; // @[:@46286.4]
  assign RetimeWrapper_42_reset = reset; // @[:@46287.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46289.4]
  assign RetimeWrapper_42_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46288.4]
  assign RetimeWrapper_43_clock = clock; // @[:@46307.4]
  assign RetimeWrapper_43_reset = reset; // @[:@46308.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46310.4]
  assign RetimeWrapper_43_io_in = x545_rdcol_1_io_result; // @[package.scala 94:16:@46309.4]
  assign RetimeWrapper_44_clock = clock; // @[:@46331.4]
  assign RetimeWrapper_44_reset = reset; // @[:@46332.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46334.4]
  assign RetimeWrapper_44_io_in = {_T_396,_T_397}; // @[package.scala 94:16:@46333.4]
  assign x626_sum_1_clock = clock; // @[:@46340.4]
  assign x626_sum_1_reset = reset; // @[:@46341.4]
  assign x626_sum_1_io_a = {_T_788,_T_789}; // @[Math.scala 151:17:@46342.4]
  assign x626_sum_1_io_b = RetimeWrapper_44_io_out; // @[Math.scala 152:17:@46343.4]
  assign x626_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@46344.4]
  assign RetimeWrapper_45_clock = clock; // @[:@46350.4]
  assign RetimeWrapper_45_reset = reset; // @[:@46351.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46353.4]
  assign RetimeWrapper_45_io_in = ~ x624; // @[package.scala 94:16:@46352.4]
  assign RetimeWrapper_46_clock = clock; // @[:@46364.4]
  assign RetimeWrapper_46_reset = reset; // @[:@46365.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46367.4]
  assign RetimeWrapper_46_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46366.4]
  assign RetimeWrapper_47_clock = clock; // @[:@46385.4]
  assign RetimeWrapper_47_reset = reset; // @[:@46386.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46388.4]
  assign RetimeWrapper_47_io_in = __1_io_result; // @[package.scala 94:16:@46387.4]
  assign RetimeWrapper_48_clock = clock; // @[:@46401.4]
  assign RetimeWrapper_48_reset = reset; // @[:@46402.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46404.4]
  assign RetimeWrapper_48_io_in = $signed(_T_936) < $signed(32'sh0); // @[package.scala 94:16:@46403.4]
  assign RetimeWrapper_49_clock = clock; // @[:@46416.4]
  assign RetimeWrapper_49_reset = reset; // @[:@46417.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46419.4]
  assign RetimeWrapper_49_io_in = {_T_342,_T_343}; // @[package.scala 94:16:@46418.4]
  assign x634_sum_1_clock = clock; // @[:@46425.4]
  assign x634_sum_1_reset = reset; // @[:@46426.4]
  assign x634_sum_1_io_a = {_T_788,_T_789}; // @[Math.scala 151:17:@46427.4]
  assign x634_sum_1_io_b = RetimeWrapper_49_io_out; // @[Math.scala 152:17:@46428.4]
  assign x634_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@46429.4]
  assign RetimeWrapper_50_clock = clock; // @[:@46435.4]
  assign RetimeWrapper_50_reset = reset; // @[:@46436.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46438.4]
  assign RetimeWrapper_50_io_in = ~ x632; // @[package.scala 94:16:@46437.4]
  assign RetimeWrapper_51_clock = clock; // @[:@46449.4]
  assign RetimeWrapper_51_reset = reset; // @[:@46450.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46452.4]
  assign RetimeWrapper_51_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46451.4]
  assign x639_rdcol_1_clock = clock; // @[:@46472.4]
  assign x639_rdcol_1_reset = reset; // @[:@46473.4]
  assign x639_rdcol_1_io_a = RetimeWrapper_47_io_out; // @[Math.scala 151:17:@46474.4]
  assign x639_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@46475.4]
  assign x639_rdcol_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@46476.4]
  assign x645_sum_1_clock = clock; // @[:@46504.4]
  assign x645_sum_1_reset = reset; // @[:@46505.4]
  assign x645_sum_1_io_a = {_T_788,_T_789}; // @[Math.scala 151:17:@46506.4]
  assign x645_sum_1_io_b = {_T_1004,_T_1005}; // @[Math.scala 152:17:@46507.4]
  assign x645_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@46508.4]
  assign RetimeWrapper_52_clock = clock; // @[:@46514.4]
  assign RetimeWrapper_52_reset = reset; // @[:@46515.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46517.4]
  assign RetimeWrapper_52_io_in = ~ x641; // @[package.scala 94:16:@46516.4]
  assign RetimeWrapper_53_clock = clock; // @[:@46528.4]
  assign RetimeWrapper_53_reset = reset; // @[:@46529.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46531.4]
  assign RetimeWrapper_53_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46530.4]
  assign x651_rdcol_1_clock = clock; // @[:@46551.4]
  assign x651_rdcol_1_reset = reset; // @[:@46552.4]
  assign x651_rdcol_1_io_a = RetimeWrapper_47_io_out; // @[Math.scala 151:17:@46553.4]
  assign x651_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@46554.4]
  assign x651_rdcol_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@46555.4]
  assign x657_sum_1_clock = clock; // @[:@46583.4]
  assign x657_sum_1_reset = reset; // @[:@46584.4]
  assign x657_sum_1_io_a = {_T_788,_T_789}; // @[Math.scala 151:17:@46585.4]
  assign x657_sum_1_io_b = {_T_1062,_T_1063}; // @[Math.scala 152:17:@46586.4]
  assign x657_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@46587.4]
  assign RetimeWrapper_54_clock = clock; // @[:@46593.4]
  assign RetimeWrapper_54_reset = reset; // @[:@46594.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46596.4]
  assign RetimeWrapper_54_io_in = ~ x653; // @[package.scala 94:16:@46595.4]
  assign RetimeWrapper_55_clock = clock; // @[:@46607.4]
  assign RetimeWrapper_55_reset = reset; // @[:@46608.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46610.4]
  assign RetimeWrapper_55_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46609.4]
  assign RetimeWrapper_56_clock = clock; // @[:@46628.4]
  assign RetimeWrapper_56_reset = reset; // @[:@46629.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46631.4]
  assign RetimeWrapper_56_io_in = __io_result; // @[package.scala 94:16:@46630.4]
  assign RetimeWrapper_57_clock = clock; // @[:@46655.4]
  assign RetimeWrapper_57_reset = reset; // @[:@46656.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46658.4]
  assign RetimeWrapper_57_io_in = $signed(_T_1104) < $signed(32'sh0); // @[package.scala 94:16:@46657.4]
  assign RetimeWrapper_58_clock = clock; // @[:@46690.4]
  assign RetimeWrapper_58_reset = reset; // @[:@46691.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46693.4]
  assign RetimeWrapper_58_io_in = {_T_1143,_T_1144}; // @[package.scala 94:16:@46692.4]
  assign x669_sum_1_clock = clock; // @[:@46701.4]
  assign x669_sum_1_reset = reset; // @[:@46702.4]
  assign x669_sum_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 151:17:@46703.4]
  assign x669_sum_1_io_b = RetimeWrapper_33_io_out; // @[Math.scala 152:17:@46704.4]
  assign x669_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@46705.4]
  assign RetimeWrapper_59_clock = clock; // @[:@46711.4]
  assign RetimeWrapper_59_reset = reset; // @[:@46712.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46714.4]
  assign RetimeWrapper_59_io_in = ~ x665; // @[package.scala 94:16:@46713.4]
  assign RetimeWrapper_60_clock = clock; // @[:@46720.4]
  assign RetimeWrapper_60_reset = reset; // @[:@46721.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46723.4]
  assign RetimeWrapper_60_io_in = $unsigned(_T_1134); // @[package.scala 94:16:@46722.4]
  assign RetimeWrapper_61_clock = clock; // @[:@46734.4]
  assign RetimeWrapper_61_reset = reset; // @[:@46735.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46737.4]
  assign RetimeWrapper_61_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46736.4]
  assign x677_sum_1_clock = clock; // @[:@46761.4]
  assign x677_sum_1_reset = reset; // @[:@46762.4]
  assign x677_sum_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 151:17:@46763.4]
  assign x677_sum_1_io_b = RetimeWrapper_40_io_out; // @[Math.scala 152:17:@46764.4]
  assign x677_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@46765.4]
  assign RetimeWrapper_62_clock = clock; // @[:@46771.4]
  assign RetimeWrapper_62_reset = reset; // @[:@46772.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46774.4]
  assign RetimeWrapper_62_io_in = ~ x675; // @[package.scala 94:16:@46773.4]
  assign RetimeWrapper_63_clock = clock; // @[:@46785.4]
  assign RetimeWrapper_63_reset = reset; // @[:@46786.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46788.4]
  assign RetimeWrapper_63_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46787.4]
  assign x684_sum_1_clock = clock; // @[:@46812.4]
  assign x684_sum_1_reset = reset; // @[:@46813.4]
  assign x684_sum_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 151:17:@46814.4]
  assign x684_sum_1_io_b = RetimeWrapper_44_io_out; // @[Math.scala 152:17:@46815.4]
  assign x684_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@46816.4]
  assign RetimeWrapper_64_clock = clock; // @[:@46822.4]
  assign RetimeWrapper_64_reset = reset; // @[:@46823.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46825.4]
  assign RetimeWrapper_64_io_in = ~ x682; // @[package.scala 94:16:@46824.4]
  assign RetimeWrapper_65_clock = clock; // @[:@46836.4]
  assign RetimeWrapper_65_reset = reset; // @[:@46837.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46839.4]
  assign RetimeWrapper_65_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46838.4]
  assign RetimeWrapper_66_clock = clock; // @[:@46863.4]
  assign RetimeWrapper_66_reset = reset; // @[:@46864.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46866.4]
  assign RetimeWrapper_66_io_in = {_T_342,_T_343}; // @[package.scala 94:16:@46865.4]
  assign x691_sum_1_clock = clock; // @[:@46872.4]
  assign x691_sum_1_reset = reset; // @[:@46873.4]
  assign x691_sum_1_io_a = {_T_1143,_T_1144}; // @[Math.scala 151:17:@46874.4]
  assign x691_sum_1_io_b = RetimeWrapper_66_io_out; // @[Math.scala 152:17:@46875.4]
  assign x691_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@46876.4]
  assign RetimeWrapper_67_clock = clock; // @[:@46882.4]
  assign RetimeWrapper_67_reset = reset; // @[:@46883.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46885.4]
  assign RetimeWrapper_67_io_in = ~ x689; // @[package.scala 94:16:@46884.4]
  assign RetimeWrapper_68_clock = clock; // @[:@46891.4]
  assign RetimeWrapper_68_reset = reset; // @[:@46892.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46894.4]
  assign RetimeWrapper_68_io_in = x691_sum_1_io_result; // @[package.scala 94:16:@46893.4]
  assign RetimeWrapper_69_clock = clock; // @[:@46905.4]
  assign RetimeWrapper_69_reset = reset; // @[:@46906.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46908.4]
  assign RetimeWrapper_69_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46907.4]
  assign x698_sum_1_clock = clock; // @[:@46932.4]
  assign x698_sum_1_reset = reset; // @[:@46933.4]
  assign x698_sum_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 151:17:@46934.4]
  assign x698_sum_1_io_b = {_T_1004,_T_1005}; // @[Math.scala 152:17:@46935.4]
  assign x698_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@46936.4]
  assign RetimeWrapper_70_clock = clock; // @[:@46942.4]
  assign RetimeWrapper_70_reset = reset; // @[:@46943.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46945.4]
  assign RetimeWrapper_70_io_in = ~ x696; // @[package.scala 94:16:@46944.4]
  assign RetimeWrapper_71_clock = clock; // @[:@46956.4]
  assign RetimeWrapper_71_reset = reset; // @[:@46957.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46959.4]
  assign RetimeWrapper_71_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@46958.4]
  assign x705_sum_1_clock = clock; // @[:@46983.4]
  assign x705_sum_1_reset = reset; // @[:@46984.4]
  assign x705_sum_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 151:17:@46985.4]
  assign x705_sum_1_io_b = {_T_1062,_T_1063}; // @[Math.scala 152:17:@46986.4]
  assign x705_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@46987.4]
  assign RetimeWrapper_72_clock = clock; // @[:@46993.4]
  assign RetimeWrapper_72_reset = reset; // @[:@46994.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@46996.4]
  assign RetimeWrapper_72_io_in = ~ x703; // @[package.scala 94:16:@46995.4]
  assign RetimeWrapper_73_clock = clock; // @[:@47007.4]
  assign RetimeWrapper_73_reset = reset; // @[:@47008.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47010.4]
  assign RetimeWrapper_73_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@47009.4]
  assign x710_rdrow_1_clock = clock; // @[:@47030.4]
  assign x710_rdrow_1_reset = reset; // @[:@47031.4]
  assign x710_rdrow_1_io_a = RetimeWrapper_56_io_out; // @[Math.scala 151:17:@47032.4]
  assign x710_rdrow_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@47033.4]
  assign x710_rdrow_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47034.4]
  assign x717_sum_1_clock = clock; // @[:@47084.4]
  assign x717_sum_1_reset = reset; // @[:@47085.4]
  assign x717_sum_1_io_a = {_T_1404,_T_1405}; // @[Math.scala 151:17:@47086.4]
  assign x717_sum_1_io_b = RetimeWrapper_33_io_out; // @[Math.scala 152:17:@47087.4]
  assign x717_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47088.4]
  assign RetimeWrapper_74_clock = clock; // @[:@47094.4]
  assign RetimeWrapper_74_reset = reset; // @[:@47095.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47097.4]
  assign RetimeWrapper_74_io_in = ~ x713; // @[package.scala 94:16:@47096.4]
  assign RetimeWrapper_75_clock = clock; // @[:@47103.4]
  assign RetimeWrapper_75_reset = reset; // @[:@47104.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47106.4]
  assign RetimeWrapper_75_io_in = $unsigned(_T_1395); // @[package.scala 94:16:@47105.4]
  assign RetimeWrapper_76_clock = clock; // @[:@47117.4]
  assign RetimeWrapper_76_reset = reset; // @[:@47118.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47120.4]
  assign RetimeWrapper_76_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@47119.4]
  assign x725_sum_1_clock = clock; // @[:@47146.4]
  assign x725_sum_1_reset = reset; // @[:@47147.4]
  assign x725_sum_1_io_a = {_T_1404,_T_1405}; // @[Math.scala 151:17:@47148.4]
  assign x725_sum_1_io_b = RetimeWrapper_40_io_out; // @[Math.scala 152:17:@47149.4]
  assign x725_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47150.4]
  assign RetimeWrapper_77_clock = clock; // @[:@47156.4]
  assign RetimeWrapper_77_reset = reset; // @[:@47157.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47159.4]
  assign RetimeWrapper_77_io_in = ~ x723; // @[package.scala 94:16:@47158.4]
  assign RetimeWrapper_78_clock = clock; // @[:@47170.4]
  assign RetimeWrapper_78_reset = reset; // @[:@47171.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47173.4]
  assign RetimeWrapper_78_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@47172.4]
  assign x732_sum_1_clock = clock; // @[:@47197.4]
  assign x732_sum_1_reset = reset; // @[:@47198.4]
  assign x732_sum_1_io_a = {_T_1404,_T_1405}; // @[Math.scala 151:17:@47199.4]
  assign x732_sum_1_io_b = RetimeWrapper_44_io_out; // @[Math.scala 152:17:@47200.4]
  assign x732_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47201.4]
  assign RetimeWrapper_79_clock = clock; // @[:@47207.4]
  assign RetimeWrapper_79_reset = reset; // @[:@47208.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47210.4]
  assign RetimeWrapper_79_io_in = ~ x730; // @[package.scala 94:16:@47209.4]
  assign RetimeWrapper_80_clock = clock; // @[:@47221.4]
  assign RetimeWrapper_80_reset = reset; // @[:@47222.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47224.4]
  assign RetimeWrapper_80_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@47223.4]
  assign x739_sum_1_clock = clock; // @[:@47248.4]
  assign x739_sum_1_reset = reset; // @[:@47249.4]
  assign x739_sum_1_io_a = {_T_1404,_T_1405}; // @[Math.scala 151:17:@47250.4]
  assign x739_sum_1_io_b = RetimeWrapper_49_io_out; // @[Math.scala 152:17:@47251.4]
  assign x739_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47252.4]
  assign RetimeWrapper_81_clock = clock; // @[:@47258.4]
  assign RetimeWrapper_81_reset = reset; // @[:@47259.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47261.4]
  assign RetimeWrapper_81_io_in = ~ x737; // @[package.scala 94:16:@47260.4]
  assign RetimeWrapper_82_clock = clock; // @[:@47272.4]
  assign RetimeWrapper_82_reset = reset; // @[:@47273.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47275.4]
  assign RetimeWrapper_82_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@47274.4]
  assign x746_sum_1_clock = clock; // @[:@47299.4]
  assign x746_sum_1_reset = reset; // @[:@47300.4]
  assign x746_sum_1_io_a = {_T_1404,_T_1405}; // @[Math.scala 151:17:@47301.4]
  assign x746_sum_1_io_b = {_T_1004,_T_1005}; // @[Math.scala 152:17:@47302.4]
  assign x746_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47303.4]
  assign RetimeWrapper_83_clock = clock; // @[:@47309.4]
  assign RetimeWrapper_83_reset = reset; // @[:@47310.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47312.4]
  assign RetimeWrapper_83_io_in = ~ x744; // @[package.scala 94:16:@47311.4]
  assign RetimeWrapper_84_clock = clock; // @[:@47323.4]
  assign RetimeWrapper_84_reset = reset; // @[:@47324.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47326.4]
  assign RetimeWrapper_84_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@47325.4]
  assign x753_sum_1_clock = clock; // @[:@47350.4]
  assign x753_sum_1_reset = reset; // @[:@47351.4]
  assign x753_sum_1_io_a = {_T_1404,_T_1405}; // @[Math.scala 151:17:@47352.4]
  assign x753_sum_1_io_b = {_T_1062,_T_1063}; // @[Math.scala 152:17:@47353.4]
  assign x753_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47354.4]
  assign RetimeWrapper_85_clock = clock; // @[:@47360.4]
  assign RetimeWrapper_85_reset = reset; // @[:@47361.4]
  assign RetimeWrapper_85_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47363.4]
  assign RetimeWrapper_85_io_in = ~ x751; // @[package.scala 94:16:@47362.4]
  assign RetimeWrapper_86_clock = clock; // @[:@47374.4]
  assign RetimeWrapper_86_reset = reset; // @[:@47375.4]
  assign RetimeWrapper_86_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47377.4]
  assign RetimeWrapper_86_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@47376.4]
  assign x758_rdrow_1_clock = clock; // @[:@47397.4]
  assign x758_rdrow_1_reset = reset; // @[:@47398.4]
  assign x758_rdrow_1_io_a = RetimeWrapper_56_io_out; // @[Math.scala 151:17:@47399.4]
  assign x758_rdrow_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@47400.4]
  assign x758_rdrow_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47401.4]
  assign x765_sum_1_clock = clock; // @[:@47451.4]
  assign x765_sum_1_reset = reset; // @[:@47452.4]
  assign x765_sum_1_io_a = {_T_1656,_T_1657}; // @[Math.scala 151:17:@47453.4]
  assign x765_sum_1_io_b = RetimeWrapper_33_io_out; // @[Math.scala 152:17:@47454.4]
  assign x765_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47455.4]
  assign RetimeWrapper_87_clock = clock; // @[:@47461.4]
  assign RetimeWrapper_87_reset = reset; // @[:@47462.4]
  assign RetimeWrapper_87_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47464.4]
  assign RetimeWrapper_87_io_in = ~ x761; // @[package.scala 94:16:@47463.4]
  assign RetimeWrapper_88_clock = clock; // @[:@47470.4]
  assign RetimeWrapper_88_reset = reset; // @[:@47471.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47473.4]
  assign RetimeWrapper_88_io_in = $unsigned(_T_1647); // @[package.scala 94:16:@47472.4]
  assign RetimeWrapper_89_clock = clock; // @[:@47484.4]
  assign RetimeWrapper_89_reset = reset; // @[:@47485.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47487.4]
  assign RetimeWrapper_89_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@47486.4]
  assign x773_sum_1_clock = clock; // @[:@47511.4]
  assign x773_sum_1_reset = reset; // @[:@47512.4]
  assign x773_sum_1_io_a = {_T_1656,_T_1657}; // @[Math.scala 151:17:@47513.4]
  assign x773_sum_1_io_b = RetimeWrapper_40_io_out; // @[Math.scala 152:17:@47514.4]
  assign x773_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47515.4]
  assign RetimeWrapper_90_clock = clock; // @[:@47521.4]
  assign RetimeWrapper_90_reset = reset; // @[:@47522.4]
  assign RetimeWrapper_90_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47524.4]
  assign RetimeWrapper_90_io_in = ~ x771; // @[package.scala 94:16:@47523.4]
  assign RetimeWrapper_91_clock = clock; // @[:@47535.4]
  assign RetimeWrapper_91_reset = reset; // @[:@47536.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47538.4]
  assign RetimeWrapper_91_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@47537.4]
  assign x780_sum_1_clock = clock; // @[:@47564.4]
  assign x780_sum_1_reset = reset; // @[:@47565.4]
  assign x780_sum_1_io_a = {_T_1656,_T_1657}; // @[Math.scala 151:17:@47566.4]
  assign x780_sum_1_io_b = RetimeWrapper_44_io_out; // @[Math.scala 152:17:@47567.4]
  assign x780_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47568.4]
  assign RetimeWrapper_92_clock = clock; // @[:@47574.4]
  assign RetimeWrapper_92_reset = reset; // @[:@47575.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47577.4]
  assign RetimeWrapper_92_io_in = ~ x778; // @[package.scala 94:16:@47576.4]
  assign RetimeWrapper_93_clock = clock; // @[:@47588.4]
  assign RetimeWrapper_93_reset = reset; // @[:@47589.4]
  assign RetimeWrapper_93_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47591.4]
  assign RetimeWrapper_93_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@47590.4]
  assign x787_sum_1_clock = clock; // @[:@47615.4]
  assign x787_sum_1_reset = reset; // @[:@47616.4]
  assign x787_sum_1_io_a = {_T_1656,_T_1657}; // @[Math.scala 151:17:@47617.4]
  assign x787_sum_1_io_b = RetimeWrapper_49_io_out; // @[Math.scala 152:17:@47618.4]
  assign x787_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47619.4]
  assign RetimeWrapper_94_clock = clock; // @[:@47625.4]
  assign RetimeWrapper_94_reset = reset; // @[:@47626.4]
  assign RetimeWrapper_94_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47628.4]
  assign RetimeWrapper_94_io_in = ~ x785; // @[package.scala 94:16:@47627.4]
  assign RetimeWrapper_95_clock = clock; // @[:@47639.4]
  assign RetimeWrapper_95_reset = reset; // @[:@47640.4]
  assign RetimeWrapper_95_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47642.4]
  assign RetimeWrapper_95_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@47641.4]
  assign x794_sum_1_clock = clock; // @[:@47666.4]
  assign x794_sum_1_reset = reset; // @[:@47667.4]
  assign x794_sum_1_io_a = {_T_1656,_T_1657}; // @[Math.scala 151:17:@47668.4]
  assign x794_sum_1_io_b = {_T_1004,_T_1005}; // @[Math.scala 152:17:@47669.4]
  assign x794_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47670.4]
  assign RetimeWrapper_96_clock = clock; // @[:@47676.4]
  assign RetimeWrapper_96_reset = reset; // @[:@47677.4]
  assign RetimeWrapper_96_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47679.4]
  assign RetimeWrapper_96_io_in = ~ x792; // @[package.scala 94:16:@47678.4]
  assign RetimeWrapper_97_clock = clock; // @[:@47690.4]
  assign RetimeWrapper_97_reset = reset; // @[:@47691.4]
  assign RetimeWrapper_97_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47693.4]
  assign RetimeWrapper_97_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@47692.4]
  assign x801_sum_1_clock = clock; // @[:@47717.4]
  assign x801_sum_1_reset = reset; // @[:@47718.4]
  assign x801_sum_1_io_a = {_T_1656,_T_1657}; // @[Math.scala 151:17:@47719.4]
  assign x801_sum_1_io_b = {_T_1062,_T_1063}; // @[Math.scala 152:17:@47720.4]
  assign x801_sum_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47721.4]
  assign RetimeWrapper_98_clock = clock; // @[:@47727.4]
  assign RetimeWrapper_98_reset = reset; // @[:@47728.4]
  assign RetimeWrapper_98_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47730.4]
  assign RetimeWrapper_98_io_in = ~ x799; // @[package.scala 94:16:@47729.4]
  assign RetimeWrapper_99_clock = clock; // @[:@47741.4]
  assign RetimeWrapper_99_reset = reset; // @[:@47742.4]
  assign RetimeWrapper_99_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47744.4]
  assign RetimeWrapper_99_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@47743.4]
  assign x811_x23_1_clock = clock; // @[:@47787.4]
  assign x811_x23_1_reset = reset; // @[:@47788.4]
  assign x811_x23_1_io_a = x524_lb_0_io_rPort_19_output_0; // @[Math.scala 151:17:@47789.4]
  assign x811_x23_1_io_b = _T_1861[7:0]; // @[Math.scala 152:17:@47790.4]
  assign x811_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47791.4]
  assign x812_x24_1_clock = clock; // @[:@47797.4]
  assign x812_x24_1_reset = reset; // @[:@47798.4]
  assign x812_x24_1_io_a = x524_lb_0_io_rPort_0_output_0; // @[Math.scala 151:17:@47799.4]
  assign x812_x24_1_io_b = _T_1865[7:0]; // @[Math.scala 152:17:@47800.4]
  assign x812_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47801.4]
  assign x813_x23_1_clock = clock; // @[:@47807.4]
  assign x813_x23_1_reset = reset; // @[:@47808.4]
  assign x813_x23_1_io_a = _T_1869[7:0]; // @[Math.scala 151:17:@47809.4]
  assign x813_x23_1_io_b = _T_1873[7:0]; // @[Math.scala 152:17:@47810.4]
  assign x813_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47811.4]
  assign x814_x24_1_clock = clock; // @[:@47817.4]
  assign x814_x24_1_reset = reset; // @[:@47818.4]
  assign x814_x24_1_io_a = x524_lb_0_io_rPort_9_output_0; // @[Math.scala 151:17:@47819.4]
  assign x814_x24_1_io_b = _T_1877[7:0]; // @[Math.scala 152:17:@47820.4]
  assign x814_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47821.4]
  assign x815_x23_1_io_a = x811_x23_1_io_result; // @[Math.scala 151:17:@47829.4]
  assign x815_x23_1_io_b = x812_x24_1_io_result; // @[Math.scala 152:17:@47830.4]
  assign x816_x24_1_io_a = x813_x23_1_io_result; // @[Math.scala 151:17:@47839.4]
  assign x816_x24_1_io_b = x814_x24_1_io_result; // @[Math.scala 152:17:@47840.4]
  assign x817_x23_1_io_a = x815_x23_1_io_result; // @[Math.scala 151:17:@47849.4]
  assign x817_x23_1_io_b = x816_x24_1_io_result; // @[Math.scala 152:17:@47850.4]
  assign RetimeWrapper_100_clock = clock; // @[:@47857.4]
  assign RetimeWrapper_100_reset = reset; // @[:@47858.4]
  assign RetimeWrapper_100_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47860.4]
  assign RetimeWrapper_100_io_in = x524_lb_0_io_rPort_21_output_0; // @[package.scala 94:16:@47859.4]
  assign x818_sum_1_io_a = x817_x23_1_io_result; // @[Math.scala 151:17:@47868.4]
  assign x818_sum_1_io_b = RetimeWrapper_100_io_out; // @[Math.scala 152:17:@47869.4]
  assign RetimeWrapper_101_clock = clock; // @[:@47880.4]
  assign RetimeWrapper_101_reset = reset; // @[:@47881.4]
  assign RetimeWrapper_101_io_flow = io_in_x512_TREADY; // @[package.scala 95:18:@47883.4]
  assign RetimeWrapper_101_io_in = {4'h0,_T_1913}; // @[package.scala 94:16:@47882.4]
  assign x825_x23_1_clock = clock; // @[:@47915.4]
  assign x825_x23_1_reset = reset; // @[:@47916.4]
  assign x825_x23_1_io_a = x524_lb_0_io_rPort_13_output_0; // @[Math.scala 151:17:@47917.4]
  assign x825_x23_1_io_b = _T_1920[7:0]; // @[Math.scala 152:17:@47918.4]
  assign x825_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47919.4]
  assign x826_x24_1_clock = clock; // @[:@47925.4]
  assign x826_x24_1_reset = reset; // @[:@47926.4]
  assign x826_x24_1_io_a = x524_lb_0_io_rPort_7_output_0; // @[Math.scala 151:17:@47927.4]
  assign x826_x24_1_io_b = _T_1924[7:0]; // @[Math.scala 152:17:@47928.4]
  assign x826_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47929.4]
  assign x827_x23_1_clock = clock; // @[:@47935.4]
  assign x827_x23_1_reset = reset; // @[:@47936.4]
  assign x827_x23_1_io_a = _T_1928[7:0]; // @[Math.scala 151:17:@47937.4]
  assign x827_x23_1_io_b = _T_1932[7:0]; // @[Math.scala 152:17:@47938.4]
  assign x827_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47939.4]
  assign x828_x24_1_clock = clock; // @[:@47945.4]
  assign x828_x24_1_reset = reset; // @[:@47946.4]
  assign x828_x24_1_io_a = x524_lb_0_io_rPort_22_output_0; // @[Math.scala 151:17:@47947.4]
  assign x828_x24_1_io_b = _T_1936[7:0]; // @[Math.scala 152:17:@47948.4]
  assign x828_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@47949.4]
  assign x829_x23_1_io_a = x825_x23_1_io_result; // @[Math.scala 151:17:@47957.4]
  assign x829_x23_1_io_b = x826_x24_1_io_result; // @[Math.scala 152:17:@47958.4]
  assign x830_x24_1_io_a = x827_x23_1_io_result; // @[Math.scala 151:17:@47967.4]
  assign x830_x24_1_io_b = x828_x24_1_io_result; // @[Math.scala 152:17:@47968.4]
  assign x831_x23_1_io_a = x829_x23_1_io_result; // @[Math.scala 151:17:@47979.4]
  assign x831_x23_1_io_b = x830_x24_1_io_result; // @[Math.scala 152:17:@47980.4]
  assign RetimeWrapper_102_clock = clock; // @[:@47987.4]
  assign RetimeWrapper_102_reset = reset; // @[:@47988.4]
  assign RetimeWrapper_102_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@47990.4]
  assign RetimeWrapper_102_io_in = x524_lb_0_io_rPort_5_output_0; // @[package.scala 94:16:@47989.4]
  assign x832_sum_1_io_a = x831_x23_1_io_result; // @[Math.scala 151:17:@47998.4]
  assign x832_sum_1_io_b = RetimeWrapper_102_io_out; // @[Math.scala 152:17:@47999.4]
  assign RetimeWrapper_103_clock = clock; // @[:@48010.4]
  assign RetimeWrapper_103_reset = reset; // @[:@48011.4]
  assign RetimeWrapper_103_io_flow = io_in_x512_TREADY; // @[package.scala 95:18:@48013.4]
  assign RetimeWrapper_103_io_in = {4'h0,_T_1974}; // @[package.scala 94:16:@48012.4]
  assign x838_x23_1_clock = clock; // @[:@48040.4]
  assign x838_x23_1_reset = reset; // @[:@48041.4]
  assign x838_x23_1_io_a = x524_lb_0_io_rPort_0_output_0; // @[Math.scala 151:17:@48042.4]
  assign x838_x23_1_io_b = _T_1981[7:0]; // @[Math.scala 152:17:@48043.4]
  assign x838_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48044.4]
  assign x839_x24_1_clock = clock; // @[:@48050.4]
  assign x839_x24_1_reset = reset; // @[:@48051.4]
  assign x839_x24_1_io_a = x524_lb_0_io_rPort_12_output_0; // @[Math.scala 151:17:@48052.4]
  assign x839_x24_1_io_b = _T_1873[7:0]; // @[Math.scala 152:17:@48053.4]
  assign x839_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48054.4]
  assign x840_x23_1_clock = clock; // @[:@48060.4]
  assign x840_x23_1_reset = reset; // @[:@48061.4]
  assign x840_x23_1_io_a = _T_1985[7:0]; // @[Math.scala 151:17:@48062.4]
  assign x840_x23_1_io_b = _T_1989[7:0]; // @[Math.scala 152:17:@48063.4]
  assign x840_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48064.4]
  assign x841_x24_1_clock = clock; // @[:@48070.4]
  assign x841_x24_1_reset = reset; // @[:@48071.4]
  assign x841_x24_1_io_a = x524_lb_0_io_rPort_21_output_0; // @[Math.scala 151:17:@48072.4]
  assign x841_x24_1_io_b = _T_1993[7:0]; // @[Math.scala 152:17:@48073.4]
  assign x841_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48074.4]
  assign x842_x23_1_io_a = x838_x23_1_io_result; // @[Math.scala 151:17:@48082.4]
  assign x842_x23_1_io_b = x839_x24_1_io_result; // @[Math.scala 152:17:@48083.4]
  assign x843_x24_1_io_a = x840_x23_1_io_result; // @[Math.scala 151:17:@48092.4]
  assign x843_x24_1_io_b = x841_x24_1_io_result; // @[Math.scala 152:17:@48093.4]
  assign x844_x23_1_io_a = x842_x23_1_io_result; // @[Math.scala 151:17:@48102.4]
  assign x844_x23_1_io_b = x843_x24_1_io_result; // @[Math.scala 152:17:@48103.4]
  assign RetimeWrapper_104_clock = clock; // @[:@48110.4]
  assign RetimeWrapper_104_reset = reset; // @[:@48111.4]
  assign RetimeWrapper_104_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48113.4]
  assign RetimeWrapper_104_io_in = x524_lb_0_io_rPort_16_output_0; // @[package.scala 94:16:@48112.4]
  assign x845_sum_1_io_a = x844_x23_1_io_result; // @[Math.scala 151:17:@48121.4]
  assign x845_sum_1_io_b = RetimeWrapper_104_io_out; // @[Math.scala 152:17:@48122.4]
  assign RetimeWrapper_105_clock = clock; // @[:@48133.4]
  assign RetimeWrapper_105_reset = reset; // @[:@48134.4]
  assign RetimeWrapper_105_io_flow = io_in_x512_TREADY; // @[package.scala 95:18:@48136.4]
  assign RetimeWrapper_105_io_in = {4'h0,_T_2029}; // @[package.scala 94:16:@48135.4]
  assign x851_x23_1_clock = clock; // @[:@48163.4]
  assign x851_x23_1_reset = reset; // @[:@48164.4]
  assign x851_x23_1_io_a = x524_lb_0_io_rPort_7_output_0; // @[Math.scala 151:17:@48165.4]
  assign x851_x23_1_io_b = _T_2036[7:0]; // @[Math.scala 152:17:@48166.4]
  assign x851_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48167.4]
  assign x852_x24_1_clock = clock; // @[:@48173.4]
  assign x852_x24_1_reset = reset; // @[:@48174.4]
  assign x852_x24_1_io_a = x524_lb_0_io_rPort_4_output_0; // @[Math.scala 151:17:@48175.4]
  assign x852_x24_1_io_b = _T_1932[7:0]; // @[Math.scala 152:17:@48176.4]
  assign x852_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48177.4]
  assign x853_x23_1_clock = clock; // @[:@48183.4]
  assign x853_x23_1_reset = reset; // @[:@48184.4]
  assign x853_x23_1_io_a = _T_2040[7:0]; // @[Math.scala 151:17:@48185.4]
  assign x853_x23_1_io_b = _T_2044[7:0]; // @[Math.scala 152:17:@48186.4]
  assign x853_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48187.4]
  assign x854_x24_1_clock = clock; // @[:@48193.4]
  assign x854_x24_1_reset = reset; // @[:@48194.4]
  assign x854_x24_1_io_a = x524_lb_0_io_rPort_5_output_0; // @[Math.scala 151:17:@48195.4]
  assign x854_x24_1_io_b = _T_2048[7:0]; // @[Math.scala 152:17:@48196.4]
  assign x854_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48197.4]
  assign x855_x23_1_io_a = x851_x23_1_io_result; // @[Math.scala 151:17:@48205.4]
  assign x855_x23_1_io_b = x852_x24_1_io_result; // @[Math.scala 152:17:@48206.4]
  assign x856_x24_1_io_a = x853_x23_1_io_result; // @[Math.scala 151:17:@48215.4]
  assign x856_x24_1_io_b = x854_x24_1_io_result; // @[Math.scala 152:17:@48216.4]
  assign x857_x23_1_io_a = x855_x23_1_io_result; // @[Math.scala 151:17:@48225.4]
  assign x857_x23_1_io_b = x856_x24_1_io_result; // @[Math.scala 152:17:@48226.4]
  assign RetimeWrapper_106_clock = clock; // @[:@48233.4]
  assign RetimeWrapper_106_reset = reset; // @[:@48234.4]
  assign RetimeWrapper_106_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48236.4]
  assign RetimeWrapper_106_io_in = x524_lb_0_io_rPort_2_output_0; // @[package.scala 94:16:@48235.4]
  assign x858_sum_1_io_a = x857_x23_1_io_result; // @[Math.scala 151:17:@48244.4]
  assign x858_sum_1_io_b = RetimeWrapper_106_io_out; // @[Math.scala 152:17:@48245.4]
  assign RetimeWrapper_107_clock = clock; // @[:@48256.4]
  assign RetimeWrapper_107_reset = reset; // @[:@48257.4]
  assign RetimeWrapper_107_io_flow = io_in_x512_TREADY; // @[package.scala 95:18:@48259.4]
  assign RetimeWrapper_107_io_in = {4'h0,_T_2084}; // @[package.scala 94:16:@48258.4]
  assign x863_x23_1_clock = clock; // @[:@48281.4]
  assign x863_x23_1_reset = reset; // @[:@48282.4]
  assign x863_x23_1_io_a = x524_lb_0_io_rPort_18_output_0; // @[Math.scala 151:17:@48283.4]
  assign x863_x23_1_io_b = _T_1924[7:0]; // @[Math.scala 152:17:@48284.4]
  assign x863_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48285.4]
  assign x864_x24_1_clock = clock; // @[:@48291.4]
  assign x864_x24_1_reset = reset; // @[:@48292.4]
  assign x864_x24_1_io_a = x524_lb_0_io_rPort_3_output_0; // @[Math.scala 151:17:@48293.4]
  assign x864_x24_1_io_b = _T_2091[7:0]; // @[Math.scala 152:17:@48294.4]
  assign x864_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48295.4]
  assign x865_x23_1_clock = clock; // @[:@48301.4]
  assign x865_x23_1_reset = reset; // @[:@48302.4]
  assign x865_x23_1_io_a = _T_2095[7:0]; // @[Math.scala 151:17:@48303.4]
  assign x865_x23_1_io_b = _T_1936[7:0]; // @[Math.scala 152:17:@48304.4]
  assign x865_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48305.4]
  assign x866_x24_1_clock = clock; // @[:@48311.4]
  assign x866_x24_1_reset = reset; // @[:@48312.4]
  assign x866_x24_1_io_a = x524_lb_0_io_rPort_14_output_0; // @[Math.scala 151:17:@48313.4]
  assign x866_x24_1_io_b = _T_2099[7:0]; // @[Math.scala 152:17:@48314.4]
  assign x866_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48315.4]
  assign x867_x23_1_io_a = x863_x23_1_io_result; // @[Math.scala 151:17:@48323.4]
  assign x867_x23_1_io_b = x864_x24_1_io_result; // @[Math.scala 152:17:@48324.4]
  assign x868_x24_1_io_a = x865_x23_1_io_result; // @[Math.scala 151:17:@48333.4]
  assign x868_x24_1_io_b = x866_x24_1_io_result; // @[Math.scala 152:17:@48334.4]
  assign x869_x23_1_io_a = x867_x23_1_io_result; // @[Math.scala 151:17:@48343.4]
  assign x869_x23_1_io_b = x868_x24_1_io_result; // @[Math.scala 152:17:@48344.4]
  assign RetimeWrapper_108_clock = clock; // @[:@48351.4]
  assign RetimeWrapper_108_reset = reset; // @[:@48352.4]
  assign RetimeWrapper_108_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48354.4]
  assign RetimeWrapper_108_io_in = x524_lb_0_io_rPort_6_output_0; // @[package.scala 94:16:@48353.4]
  assign x870_sum_1_io_a = x869_x23_1_io_result; // @[Math.scala 151:17:@48362.4]
  assign x870_sum_1_io_b = RetimeWrapper_108_io_out; // @[Math.scala 152:17:@48363.4]
  assign RetimeWrapper_109_clock = clock; // @[:@48374.4]
  assign RetimeWrapper_109_reset = reset; // @[:@48375.4]
  assign RetimeWrapper_109_io_flow = io_in_x512_TREADY; // @[package.scala 95:18:@48377.4]
  assign RetimeWrapper_109_io_in = {4'h0,_T_2135}; // @[package.scala 94:16:@48376.4]
  assign x874_x23_1_clock = clock; // @[:@48394.4]
  assign x874_x23_1_reset = reset; // @[:@48395.4]
  assign x874_x23_1_io_a = x524_lb_0_io_rPort_15_output_0; // @[Math.scala 151:17:@48396.4]
  assign x874_x23_1_io_b = _T_1873[7:0]; // @[Math.scala 152:17:@48397.4]
  assign x874_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48398.4]
  assign x875_x24_1_clock = clock; // @[:@48404.4]
  assign x875_x24_1_reset = reset; // @[:@48405.4]
  assign x875_x24_1_io_a = x524_lb_0_io_rPort_10_output_0; // @[Math.scala 151:17:@48406.4]
  assign x875_x24_1_io_b = _T_1877[7:0]; // @[Math.scala 152:17:@48407.4]
  assign x875_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48408.4]
  assign x876_x23_1_clock = clock; // @[:@48416.4]
  assign x876_x23_1_reset = reset; // @[:@48417.4]
  assign x876_x23_1_io_a = _T_2142[7:0]; // @[Math.scala 151:17:@48418.4]
  assign x876_x23_1_io_b = _T_1993[7:0]; // @[Math.scala 152:17:@48419.4]
  assign x876_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48420.4]
  assign x877_x24_1_clock = clock; // @[:@48426.4]
  assign x877_x24_1_reset = reset; // @[:@48427.4]
  assign x877_x24_1_io_a = x524_lb_0_io_rPort_17_output_0; // @[Math.scala 151:17:@48428.4]
  assign x877_x24_1_io_b = _T_2146[7:0]; // @[Math.scala 152:17:@48429.4]
  assign x877_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48430.4]
  assign x878_x23_1_io_a = x874_x23_1_io_result; // @[Math.scala 151:17:@48438.4]
  assign x878_x23_1_io_b = x875_x24_1_io_result; // @[Math.scala 152:17:@48439.4]
  assign x879_x24_1_io_a = x876_x23_1_io_result; // @[Math.scala 151:17:@48448.4]
  assign x879_x24_1_io_b = x877_x24_1_io_result; // @[Math.scala 152:17:@48449.4]
  assign x880_x23_1_io_a = x878_x23_1_io_result; // @[Math.scala 151:17:@48458.4]
  assign x880_x23_1_io_b = x879_x24_1_io_result; // @[Math.scala 152:17:@48459.4]
  assign RetimeWrapper_110_clock = clock; // @[:@48466.4]
  assign RetimeWrapper_110_reset = reset; // @[:@48467.4]
  assign RetimeWrapper_110_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48469.4]
  assign RetimeWrapper_110_io_in = x524_lb_0_io_rPort_20_output_0; // @[package.scala 94:16:@48468.4]
  assign x881_sum_1_io_a = x880_x23_1_io_result; // @[Math.scala 151:17:@48477.4]
  assign x881_sum_1_io_b = RetimeWrapper_110_io_out; // @[Math.scala 152:17:@48478.4]
  assign RetimeWrapper_111_clock = clock; // @[:@48489.4]
  assign RetimeWrapper_111_reset = reset; // @[:@48490.4]
  assign RetimeWrapper_111_io_flow = io_in_x512_TREADY; // @[package.scala 95:18:@48492.4]
  assign RetimeWrapper_111_io_in = {4'h0,_T_2184}; // @[package.scala 94:16:@48491.4]
  assign x885_x23_1_clock = clock; // @[:@48509.4]
  assign x885_x23_1_reset = reset; // @[:@48510.4]
  assign x885_x23_1_io_a = x524_lb_0_io_rPort_3_output_0; // @[Math.scala 151:17:@48511.4]
  assign x885_x23_1_io_b = _T_1932[7:0]; // @[Math.scala 152:17:@48512.4]
  assign x885_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48513.4]
  assign x886_x24_1_clock = clock; // @[:@48519.4]
  assign x886_x24_1_reset = reset; // @[:@48520.4]
  assign x886_x24_1_io_a = x524_lb_0_io_rPort_8_output_0; // @[Math.scala 151:17:@48521.4]
  assign x886_x24_1_io_b = _T_1936[7:0]; // @[Math.scala 152:17:@48522.4]
  assign x886_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48523.4]
  assign x887_x23_1_clock = clock; // @[:@48529.4]
  assign x887_x23_1_reset = reset; // @[:@48530.4]
  assign x887_x23_1_io_a = _T_2191[7:0]; // @[Math.scala 151:17:@48531.4]
  assign x887_x23_1_io_b = _T_2048[7:0]; // @[Math.scala 152:17:@48532.4]
  assign x887_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48533.4]
  assign x888_x24_1_clock = clock; // @[:@48539.4]
  assign x888_x24_1_reset = reset; // @[:@48540.4]
  assign x888_x24_1_io_a = x524_lb_0_io_rPort_6_output_0; // @[Math.scala 151:17:@48541.4]
  assign x888_x24_1_io_b = _T_2195[7:0]; // @[Math.scala 152:17:@48542.4]
  assign x888_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48543.4]
  assign x889_x23_1_io_a = x885_x23_1_io_result; // @[Math.scala 151:17:@48551.4]
  assign x889_x23_1_io_b = x886_x24_1_io_result; // @[Math.scala 152:17:@48552.4]
  assign x890_x24_1_io_a = x887_x23_1_io_result; // @[Math.scala 151:17:@48561.4]
  assign x890_x24_1_io_b = x888_x24_1_io_result; // @[Math.scala 152:17:@48562.4]
  assign x891_x23_1_io_a = x889_x23_1_io_result; // @[Math.scala 151:17:@48571.4]
  assign x891_x23_1_io_b = x890_x24_1_io_result; // @[Math.scala 152:17:@48572.4]
  assign RetimeWrapper_112_clock = clock; // @[:@48579.4]
  assign RetimeWrapper_112_reset = reset; // @[:@48580.4]
  assign RetimeWrapper_112_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48582.4]
  assign RetimeWrapper_112_io_in = x524_lb_0_io_rPort_1_output_0; // @[package.scala 94:16:@48581.4]
  assign x892_sum_1_io_a = x891_x23_1_io_result; // @[Math.scala 151:17:@48590.4]
  assign x892_sum_1_io_b = RetimeWrapper_112_io_out; // @[Math.scala 152:17:@48591.4]
  assign RetimeWrapper_113_clock = clock; // @[:@48602.4]
  assign RetimeWrapper_113_reset = reset; // @[:@48603.4]
  assign RetimeWrapper_113_io_flow = io_in_x512_TREADY; // @[package.scala 95:18:@48605.4]
  assign RetimeWrapper_113_io_in = {4'h0,_T_2231}; // @[package.scala 94:16:@48604.4]
  assign x897_x23_1_clock = clock; // @[:@48627.4]
  assign x897_x23_1_reset = reset; // @[:@48628.4]
  assign x897_x23_1_io_a = x524_lb_0_io_rPort_10_output_0; // @[Math.scala 151:17:@48629.4]
  assign x897_x23_1_io_b = _T_1989[7:0]; // @[Math.scala 152:17:@48630.4]
  assign x897_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48631.4]
  assign x898_x24_1_clock = clock; // @[:@48637.4]
  assign x898_x24_1_reset = reset; // @[:@48638.4]
  assign x898_x24_1_io_a = x524_lb_0_io_rPort_23_output_0; // @[Math.scala 151:17:@48639.4]
  assign x898_x24_1_io_b = _T_1993[7:0]; // @[Math.scala 152:17:@48640.4]
  assign x898_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48641.4]
  assign x899_x23_1_clock = clock; // @[:@48647.4]
  assign x899_x23_1_reset = reset; // @[:@48648.4]
  assign x899_x23_1_io_a = _T_2238[7:0]; // @[Math.scala 151:17:@48649.4]
  assign x899_x23_1_io_b = _T_2242[7:0]; // @[Math.scala 152:17:@48650.4]
  assign x899_x23_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48651.4]
  assign x900_x24_1_clock = clock; // @[:@48657.4]
  assign x900_x24_1_reset = reset; // @[:@48658.4]
  assign x900_x24_1_io_a = x524_lb_0_io_rPort_20_output_0; // @[Math.scala 151:17:@48659.4]
  assign x900_x24_1_io_b = _T_2246[7:0]; // @[Math.scala 152:17:@48660.4]
  assign x900_x24_1_io_flow = io_in_x512_TREADY; // @[Math.scala 153:20:@48661.4]
  assign x901_x23_1_io_a = x897_x23_1_io_result; // @[Math.scala 151:17:@48669.4]
  assign x901_x23_1_io_b = x898_x24_1_io_result; // @[Math.scala 152:17:@48670.4]
  assign x902_x24_1_io_a = x899_x23_1_io_result; // @[Math.scala 151:17:@48679.4]
  assign x902_x24_1_io_b = x900_x24_1_io_result; // @[Math.scala 152:17:@48680.4]
  assign x903_x23_1_io_a = x901_x23_1_io_result; // @[Math.scala 151:17:@48689.4]
  assign x903_x23_1_io_b = x902_x24_1_io_result; // @[Math.scala 152:17:@48690.4]
  assign RetimeWrapper_114_clock = clock; // @[:@48697.4]
  assign RetimeWrapper_114_reset = reset; // @[:@48698.4]
  assign RetimeWrapper_114_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48700.4]
  assign RetimeWrapper_114_io_in = x524_lb_0_io_rPort_11_output_0; // @[package.scala 94:16:@48699.4]
  assign x904_sum_1_io_a = x903_x23_1_io_result; // @[Math.scala 151:17:@48708.4]
  assign x904_sum_1_io_b = RetimeWrapper_114_io_out; // @[Math.scala 152:17:@48709.4]
  assign RetimeWrapper_115_clock = clock; // @[:@48720.4]
  assign RetimeWrapper_115_reset = reset; // @[:@48721.4]
  assign RetimeWrapper_115_io_flow = io_in_x512_TREADY; // @[package.scala 95:18:@48723.4]
  assign RetimeWrapper_115_io_in = {4'h0,_T_2282}; // @[package.scala 94:16:@48722.4]
  assign RetimeWrapper_116_clock = clock; // @[:@48730.4]
  assign RetimeWrapper_116_reset = reset; // @[:@48731.4]
  assign RetimeWrapper_116_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48733.4]
  assign RetimeWrapper_116_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@48732.4]
  assign RetimeWrapper_117_clock = clock; // @[:@48739.4]
  assign RetimeWrapper_117_reset = reset; // @[:@48740.4]
  assign RetimeWrapper_117_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48742.4]
  assign RetimeWrapper_117_io_in = $unsigned(_T_323); // @[package.scala 94:16:@48741.4]
  assign RetimeWrapper_118_clock = clock; // @[:@48748.4]
  assign RetimeWrapper_118_reset = reset; // @[:@48749.4]
  assign RetimeWrapper_118_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48751.4]
  assign RetimeWrapper_118_io_in = RetimeWrapper_115_io_out; // @[package.scala 94:16:@48750.4]
  assign RetimeWrapper_119_clock = clock; // @[:@48757.4]
  assign RetimeWrapper_119_reset = reset; // @[:@48758.4]
  assign RetimeWrapper_119_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48760.4]
  assign RetimeWrapper_119_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@48759.4]
  assign RetimeWrapper_120_clock = clock; // @[:@48766.4]
  assign RetimeWrapper_120_reset = reset; // @[:@48767.4]
  assign RetimeWrapper_120_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48769.4]
  assign RetimeWrapper_120_io_in = x539_sum_1_io_result; // @[package.scala 94:16:@48768.4]
  assign RetimeWrapper_121_clock = clock; // @[:@48779.4]
  assign RetimeWrapper_121_reset = reset; // @[:@48780.4]
  assign RetimeWrapper_121_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48782.4]
  assign RetimeWrapper_121_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@48781.4]
  assign RetimeWrapper_122_clock = clock; // @[:@48800.4]
  assign RetimeWrapper_122_reset = reset; // @[:@48801.4]
  assign RetimeWrapper_122_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48803.4]
  assign RetimeWrapper_122_io_in = RetimeWrapper_113_io_out; // @[package.scala 94:16:@48802.4]
  assign RetimeWrapper_123_clock = clock; // @[:@48809.4]
  assign RetimeWrapper_123_reset = reset; // @[:@48810.4]
  assign RetimeWrapper_123_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48812.4]
  assign RetimeWrapper_123_io_in = x549_sum_1_io_result; // @[package.scala 94:16:@48811.4]
  assign RetimeWrapper_124_clock = clock; // @[:@48822.4]
  assign RetimeWrapper_124_reset = reset; // @[:@48823.4]
  assign RetimeWrapper_124_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48825.4]
  assign RetimeWrapper_124_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@48824.4]
  assign RetimeWrapper_125_clock = clock; // @[:@48843.4]
  assign RetimeWrapper_125_reset = reset; // @[:@48844.4]
  assign RetimeWrapper_125_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48846.4]
  assign RetimeWrapper_125_io_in = x558_sum_1_io_result; // @[package.scala 94:16:@48845.4]
  assign RetimeWrapper_126_clock = clock; // @[:@48852.4]
  assign RetimeWrapper_126_reset = reset; // @[:@48853.4]
  assign RetimeWrapper_126_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48855.4]
  assign RetimeWrapper_126_io_in = RetimeWrapper_111_io_out; // @[package.scala 94:16:@48854.4]
  assign RetimeWrapper_127_clock = clock; // @[:@48865.4]
  assign RetimeWrapper_127_reset = reset; // @[:@48866.4]
  assign RetimeWrapper_127_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48868.4]
  assign RetimeWrapper_127_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@48867.4]
  assign RetimeWrapper_128_clock = clock; // @[:@48886.4]
  assign RetimeWrapper_128_reset = reset; // @[:@48887.4]
  assign RetimeWrapper_128_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48889.4]
  assign RetimeWrapper_128_io_in = x567_sum_1_io_result; // @[package.scala 94:16:@48888.4]
  assign RetimeWrapper_129_clock = clock; // @[:@48895.4]
  assign RetimeWrapper_129_reset = reset; // @[:@48896.4]
  assign RetimeWrapper_129_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48898.4]
  assign RetimeWrapper_129_io_in = RetimeWrapper_109_io_out; // @[package.scala 94:16:@48897.4]
  assign RetimeWrapper_130_clock = clock; // @[:@48908.4]
  assign RetimeWrapper_130_reset = reset; // @[:@48909.4]
  assign RetimeWrapper_130_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48911.4]
  assign RetimeWrapper_130_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@48910.4]
  assign RetimeWrapper_131_clock = clock; // @[:@48929.4]
  assign RetimeWrapper_131_reset = reset; // @[:@48930.4]
  assign RetimeWrapper_131_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48932.4]
  assign RetimeWrapper_131_io_in = $unsigned(_T_602); // @[package.scala 94:16:@48931.4]
  assign RetimeWrapper_132_clock = clock; // @[:@48938.4]
  assign RetimeWrapper_132_reset = reset; // @[:@48939.4]
  assign RetimeWrapper_132_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48941.4]
  assign RetimeWrapper_132_io_in = RetimeWrapper_107_io_out; // @[package.scala 94:16:@48940.4]
  assign RetimeWrapper_133_clock = clock; // @[:@48947.4]
  assign RetimeWrapper_133_reset = reset; // @[:@48948.4]
  assign RetimeWrapper_133_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48950.4]
  assign RetimeWrapper_133_io_in = x581_sum_1_io_result; // @[package.scala 94:16:@48949.4]
  assign RetimeWrapper_134_clock = clock; // @[:@48960.4]
  assign RetimeWrapper_134_reset = reset; // @[:@48961.4]
  assign RetimeWrapper_134_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48963.4]
  assign RetimeWrapper_134_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@48962.4]
  assign RetimeWrapper_135_clock = clock; // @[:@48981.4]
  assign RetimeWrapper_135_reset = reset; // @[:@48982.4]
  assign RetimeWrapper_135_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48984.4]
  assign RetimeWrapper_135_io_in = RetimeWrapper_105_io_out; // @[package.scala 94:16:@48983.4]
  assign RetimeWrapper_136_clock = clock; // @[:@48990.4]
  assign RetimeWrapper_136_reset = reset; // @[:@48991.4]
  assign RetimeWrapper_136_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@48993.4]
  assign RetimeWrapper_136_io_in = x587_sum_1_io_result; // @[package.scala 94:16:@48992.4]
  assign RetimeWrapper_137_clock = clock; // @[:@49003.4]
  assign RetimeWrapper_137_reset = reset; // @[:@49004.4]
  assign RetimeWrapper_137_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49006.4]
  assign RetimeWrapper_137_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49005.4]
  assign RetimeWrapper_138_clock = clock; // @[:@49024.4]
  assign RetimeWrapper_138_reset = reset; // @[:@49025.4]
  assign RetimeWrapper_138_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49027.4]
  assign RetimeWrapper_138_io_in = RetimeWrapper_103_io_out; // @[package.scala 94:16:@49026.4]
  assign RetimeWrapper_139_clock = clock; // @[:@49033.4]
  assign RetimeWrapper_139_reset = reset; // @[:@49034.4]
  assign RetimeWrapper_139_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49036.4]
  assign RetimeWrapper_139_io_in = x592_sum_1_io_result; // @[package.scala 94:16:@49035.4]
  assign RetimeWrapper_140_clock = clock; // @[:@49046.4]
  assign RetimeWrapper_140_reset = reset; // @[:@49047.4]
  assign RetimeWrapper_140_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49049.4]
  assign RetimeWrapper_140_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49048.4]
  assign RetimeWrapper_141_clock = clock; // @[:@49067.4]
  assign RetimeWrapper_141_reset = reset; // @[:@49068.4]
  assign RetimeWrapper_141_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49070.4]
  assign RetimeWrapper_141_io_in = x597_sum_1_io_result; // @[package.scala 94:16:@49069.4]
  assign RetimeWrapper_142_clock = clock; // @[:@49076.4]
  assign RetimeWrapper_142_reset = reset; // @[:@49077.4]
  assign RetimeWrapper_142_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49079.4]
  assign RetimeWrapper_142_io_in = RetimeWrapper_101_io_out; // @[package.scala 94:16:@49078.4]
  assign RetimeWrapper_143_clock = clock; // @[:@49089.4]
  assign RetimeWrapper_143_reset = reset; // @[:@49090.4]
  assign RetimeWrapper_143_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49092.4]
  assign RetimeWrapper_143_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49091.4]
  assign RetimeWrapper_144_clock = clock; // @[:@49110.4]
  assign RetimeWrapper_144_reset = reset; // @[:@49111.4]
  assign RetimeWrapper_144_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49113.4]
  assign RetimeWrapper_144_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@49112.4]
  assign RetimeWrapper_145_clock = clock; // @[:@49119.4]
  assign RetimeWrapper_145_reset = reset; // @[:@49120.4]
  assign RetimeWrapper_145_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49122.4]
  assign RetimeWrapper_145_io_in = ~ x605; // @[package.scala 94:16:@49121.4]
  assign RetimeWrapper_146_clock = clock; // @[:@49128.4]
  assign RetimeWrapper_146_reset = reset; // @[:@49129.4]
  assign RetimeWrapper_146_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49131.4]
  assign RetimeWrapper_146_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@49130.4]
  assign RetimeWrapper_147_clock = clock; // @[:@49137.4]
  assign RetimeWrapper_147_reset = reset; // @[:@49138.4]
  assign RetimeWrapper_147_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49140.4]
  assign RetimeWrapper_147_io_in = $unsigned(_T_779); // @[package.scala 94:16:@49139.4]
  assign RetimeWrapper_148_clock = clock; // @[:@49146.4]
  assign RetimeWrapper_148_reset = reset; // @[:@49147.4]
  assign RetimeWrapper_148_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49149.4]
  assign RetimeWrapper_148_io_in = x609_sum_1_io_result; // @[package.scala 94:16:@49148.4]
  assign RetimeWrapper_149_clock = clock; // @[:@49160.4]
  assign RetimeWrapper_149_reset = reset; // @[:@49161.4]
  assign RetimeWrapper_149_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49163.4]
  assign RetimeWrapper_149_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49162.4]
  assign RetimeWrapper_150_clock = clock; // @[:@49181.4]
  assign RetimeWrapper_150_reset = reset; // @[:@49182.4]
  assign RetimeWrapper_150_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49184.4]
  assign RetimeWrapper_150_io_in = x618_sum_1_io_result; // @[package.scala 94:16:@49183.4]
  assign RetimeWrapper_151_clock = clock; // @[:@49190.4]
  assign RetimeWrapper_151_reset = reset; // @[:@49191.4]
  assign RetimeWrapper_151_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49193.4]
  assign RetimeWrapper_151_io_in = ~ x616; // @[package.scala 94:16:@49192.4]
  assign RetimeWrapper_152_clock = clock; // @[:@49204.4]
  assign RetimeWrapper_152_reset = reset; // @[:@49205.4]
  assign RetimeWrapper_152_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49207.4]
  assign RetimeWrapper_152_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49206.4]
  assign RetimeWrapper_153_clock = clock; // @[:@49225.4]
  assign RetimeWrapper_153_reset = reset; // @[:@49226.4]
  assign RetimeWrapper_153_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49228.4]
  assign RetimeWrapper_153_io_in = ~ x624; // @[package.scala 94:16:@49227.4]
  assign RetimeWrapper_154_clock = clock; // @[:@49234.4]
  assign RetimeWrapper_154_reset = reset; // @[:@49235.4]
  assign RetimeWrapper_154_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49237.4]
  assign RetimeWrapper_154_io_in = x626_sum_1_io_result; // @[package.scala 94:16:@49236.4]
  assign RetimeWrapper_155_clock = clock; // @[:@49248.4]
  assign RetimeWrapper_155_reset = reset; // @[:@49249.4]
  assign RetimeWrapper_155_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49251.4]
  assign RetimeWrapper_155_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49250.4]
  assign RetimeWrapper_156_clock = clock; // @[:@49269.4]
  assign RetimeWrapper_156_reset = reset; // @[:@49270.4]
  assign RetimeWrapper_156_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49272.4]
  assign RetimeWrapper_156_io_in = x634_sum_1_io_result; // @[package.scala 94:16:@49271.4]
  assign RetimeWrapper_157_clock = clock; // @[:@49278.4]
  assign RetimeWrapper_157_reset = reset; // @[:@49279.4]
  assign RetimeWrapper_157_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49281.4]
  assign RetimeWrapper_157_io_in = ~ x632; // @[package.scala 94:16:@49280.4]
  assign RetimeWrapper_158_clock = clock; // @[:@49292.4]
  assign RetimeWrapper_158_reset = reset; // @[:@49293.4]
  assign RetimeWrapper_158_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49295.4]
  assign RetimeWrapper_158_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49294.4]
  assign RetimeWrapper_159_clock = clock; // @[:@49313.4]
  assign RetimeWrapper_159_reset = reset; // @[:@49314.4]
  assign RetimeWrapper_159_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49316.4]
  assign RetimeWrapper_159_io_in = x645_sum_1_io_result; // @[package.scala 94:16:@49315.4]
  assign RetimeWrapper_160_clock = clock; // @[:@49322.4]
  assign RetimeWrapper_160_reset = reset; // @[:@49323.4]
  assign RetimeWrapper_160_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49325.4]
  assign RetimeWrapper_160_io_in = ~ x641; // @[package.scala 94:16:@49324.4]
  assign RetimeWrapper_161_clock = clock; // @[:@49336.4]
  assign RetimeWrapper_161_reset = reset; // @[:@49337.4]
  assign RetimeWrapper_161_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49339.4]
  assign RetimeWrapper_161_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49338.4]
  assign RetimeWrapper_162_clock = clock; // @[:@49357.4]
  assign RetimeWrapper_162_reset = reset; // @[:@49358.4]
  assign RetimeWrapper_162_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49360.4]
  assign RetimeWrapper_162_io_in = ~ x665; // @[package.scala 94:16:@49359.4]
  assign RetimeWrapper_163_clock = clock; // @[:@49366.4]
  assign RetimeWrapper_163_reset = reset; // @[:@49367.4]
  assign RetimeWrapper_163_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49369.4]
  assign RetimeWrapper_163_io_in = x669_sum_1_io_result; // @[package.scala 94:16:@49368.4]
  assign RetimeWrapper_164_clock = clock; // @[:@49375.4]
  assign RetimeWrapper_164_reset = reset; // @[:@49376.4]
  assign RetimeWrapper_164_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49378.4]
  assign RetimeWrapper_164_io_in = $unsigned(_T_1134); // @[package.scala 94:16:@49377.4]
  assign RetimeWrapper_165_clock = clock; // @[:@49389.4]
  assign RetimeWrapper_165_reset = reset; // @[:@49390.4]
  assign RetimeWrapper_165_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49392.4]
  assign RetimeWrapper_165_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49391.4]
  assign RetimeWrapper_166_clock = clock; // @[:@49410.4]
  assign RetimeWrapper_166_reset = reset; // @[:@49411.4]
  assign RetimeWrapper_166_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49413.4]
  assign RetimeWrapper_166_io_in = x677_sum_1_io_result; // @[package.scala 94:16:@49412.4]
  assign RetimeWrapper_167_clock = clock; // @[:@49419.4]
  assign RetimeWrapper_167_reset = reset; // @[:@49420.4]
  assign RetimeWrapper_167_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49422.4]
  assign RetimeWrapper_167_io_in = ~ x675; // @[package.scala 94:16:@49421.4]
  assign RetimeWrapper_168_clock = clock; // @[:@49433.4]
  assign RetimeWrapper_168_reset = reset; // @[:@49434.4]
  assign RetimeWrapper_168_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49436.4]
  assign RetimeWrapper_168_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49435.4]
  assign RetimeWrapper_169_clock = clock; // @[:@49454.4]
  assign RetimeWrapper_169_reset = reset; // @[:@49455.4]
  assign RetimeWrapper_169_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49457.4]
  assign RetimeWrapper_169_io_in = ~ x682; // @[package.scala 94:16:@49456.4]
  assign RetimeWrapper_170_clock = clock; // @[:@49463.4]
  assign RetimeWrapper_170_reset = reset; // @[:@49464.4]
  assign RetimeWrapper_170_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49466.4]
  assign RetimeWrapper_170_io_in = x684_sum_1_io_result; // @[package.scala 94:16:@49465.4]
  assign RetimeWrapper_171_clock = clock; // @[:@49477.4]
  assign RetimeWrapper_171_reset = reset; // @[:@49478.4]
  assign RetimeWrapper_171_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49480.4]
  assign RetimeWrapper_171_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49479.4]
  assign RetimeWrapper_172_clock = clock; // @[:@49498.4]
  assign RetimeWrapper_172_reset = reset; // @[:@49499.4]
  assign RetimeWrapper_172_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49501.4]
  assign RetimeWrapper_172_io_in = ~ x689; // @[package.scala 94:16:@49500.4]
  assign RetimeWrapper_173_clock = clock; // @[:@49507.4]
  assign RetimeWrapper_173_reset = reset; // @[:@49508.4]
  assign RetimeWrapper_173_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49510.4]
  assign RetimeWrapper_173_io_in = x691_sum_1_io_result; // @[package.scala 94:16:@49509.4]
  assign RetimeWrapper_174_clock = clock; // @[:@49521.4]
  assign RetimeWrapper_174_reset = reset; // @[:@49522.4]
  assign RetimeWrapper_174_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49524.4]
  assign RetimeWrapper_174_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49523.4]
  assign RetimeWrapper_175_clock = clock; // @[:@49542.4]
  assign RetimeWrapper_175_reset = reset; // @[:@49543.4]
  assign RetimeWrapper_175_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49545.4]
  assign RetimeWrapper_175_io_in = x698_sum_1_io_result; // @[package.scala 94:16:@49544.4]
  assign RetimeWrapper_176_clock = clock; // @[:@49551.4]
  assign RetimeWrapper_176_reset = reset; // @[:@49552.4]
  assign RetimeWrapper_176_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49554.4]
  assign RetimeWrapper_176_io_in = ~ x696; // @[package.scala 94:16:@49553.4]
  assign RetimeWrapper_177_clock = clock; // @[:@49565.4]
  assign RetimeWrapper_177_reset = reset; // @[:@49566.4]
  assign RetimeWrapper_177_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49568.4]
  assign RetimeWrapper_177_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49567.4]
  assign RetimeWrapper_178_clock = clock; // @[:@49586.4]
  assign RetimeWrapper_178_reset = reset; // @[:@49587.4]
  assign RetimeWrapper_178_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49589.4]
  assign RetimeWrapper_178_io_in = ~ x713; // @[package.scala 94:16:@49588.4]
  assign RetimeWrapper_179_clock = clock; // @[:@49595.4]
  assign RetimeWrapper_179_reset = reset; // @[:@49596.4]
  assign RetimeWrapper_179_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49598.4]
  assign RetimeWrapper_179_io_in = $unsigned(_T_1395); // @[package.scala 94:16:@49597.4]
  assign RetimeWrapper_180_clock = clock; // @[:@49604.4]
  assign RetimeWrapper_180_reset = reset; // @[:@49605.4]
  assign RetimeWrapper_180_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49607.4]
  assign RetimeWrapper_180_io_in = x717_sum_1_io_result; // @[package.scala 94:16:@49606.4]
  assign RetimeWrapper_181_clock = clock; // @[:@49618.4]
  assign RetimeWrapper_181_reset = reset; // @[:@49619.4]
  assign RetimeWrapper_181_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49621.4]
  assign RetimeWrapper_181_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49620.4]
  assign RetimeWrapper_182_clock = clock; // @[:@49639.4]
  assign RetimeWrapper_182_reset = reset; // @[:@49640.4]
  assign RetimeWrapper_182_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49642.4]
  assign RetimeWrapper_182_io_in = ~ x723; // @[package.scala 94:16:@49641.4]
  assign RetimeWrapper_183_clock = clock; // @[:@49648.4]
  assign RetimeWrapper_183_reset = reset; // @[:@49649.4]
  assign RetimeWrapper_183_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49651.4]
  assign RetimeWrapper_183_io_in = x725_sum_1_io_result; // @[package.scala 94:16:@49650.4]
  assign RetimeWrapper_184_clock = clock; // @[:@49662.4]
  assign RetimeWrapper_184_reset = reset; // @[:@49663.4]
  assign RetimeWrapper_184_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49665.4]
  assign RetimeWrapper_184_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49664.4]
  assign RetimeWrapper_185_clock = clock; // @[:@49683.4]
  assign RetimeWrapper_185_reset = reset; // @[:@49684.4]
  assign RetimeWrapper_185_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49686.4]
  assign RetimeWrapper_185_io_in = x732_sum_1_io_result; // @[package.scala 94:16:@49685.4]
  assign RetimeWrapper_186_clock = clock; // @[:@49692.4]
  assign RetimeWrapper_186_reset = reset; // @[:@49693.4]
  assign RetimeWrapper_186_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49695.4]
  assign RetimeWrapper_186_io_in = ~ x730; // @[package.scala 94:16:@49694.4]
  assign RetimeWrapper_187_clock = clock; // @[:@49706.4]
  assign RetimeWrapper_187_reset = reset; // @[:@49707.4]
  assign RetimeWrapper_187_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49709.4]
  assign RetimeWrapper_187_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49708.4]
  assign RetimeWrapper_188_clock = clock; // @[:@49727.4]
  assign RetimeWrapper_188_reset = reset; // @[:@49728.4]
  assign RetimeWrapper_188_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49730.4]
  assign RetimeWrapper_188_io_in = ~ x737; // @[package.scala 94:16:@49729.4]
  assign RetimeWrapper_189_clock = clock; // @[:@49736.4]
  assign RetimeWrapper_189_reset = reset; // @[:@49737.4]
  assign RetimeWrapper_189_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49739.4]
  assign RetimeWrapper_189_io_in = x739_sum_1_io_result; // @[package.scala 94:16:@49738.4]
  assign RetimeWrapper_190_clock = clock; // @[:@49750.4]
  assign RetimeWrapper_190_reset = reset; // @[:@49751.4]
  assign RetimeWrapper_190_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49753.4]
  assign RetimeWrapper_190_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49752.4]
  assign RetimeWrapper_191_clock = clock; // @[:@49771.4]
  assign RetimeWrapper_191_reset = reset; // @[:@49772.4]
  assign RetimeWrapper_191_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49774.4]
  assign RetimeWrapper_191_io_in = x746_sum_1_io_result; // @[package.scala 94:16:@49773.4]
  assign RetimeWrapper_192_clock = clock; // @[:@49780.4]
  assign RetimeWrapper_192_reset = reset; // @[:@49781.4]
  assign RetimeWrapper_192_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49783.4]
  assign RetimeWrapper_192_io_in = ~ x744; // @[package.scala 94:16:@49782.4]
  assign RetimeWrapper_193_clock = clock; // @[:@49794.4]
  assign RetimeWrapper_193_reset = reset; // @[:@49795.4]
  assign RetimeWrapper_193_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@49797.4]
  assign RetimeWrapper_193_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49796.4]
  assign x948_x25_1_io_a = x525_lb2_0_io_rPort_5_output_0; // @[Math.scala 151:17:@49829.4]
  assign x948_x25_1_io_b = _T_2945[7:0]; // @[Math.scala 152:17:@49830.4]
  assign x949_x26_1_io_a = _T_2949[7:0]; // @[Math.scala 151:17:@49839.4]
  assign x949_x26_1_io_b = x525_lb2_0_io_rPort_13_output_0; // @[Math.scala 152:17:@49840.4]
  assign x950_sum_1_io_a = x948_x25_1_io_result; // @[Math.scala 151:17:@49849.4]
  assign x950_sum_1_io_b = x949_x26_1_io_result; // @[Math.scala 152:17:@49850.4]
  assign x951_div_1_clock = clock; // @[:@49859.4]
  assign x951_div_1_reset = reset; // @[:@49860.4]
  assign x951_div_1_io_a = x950_sum_1_io_result; // @[Math.scala 328:17:@49861.4]
  assign x951_div_1_io_flow = io_in_x512_TREADY; // @[Math.scala 330:20:@49863.4]
  assign x954_x25_1_io_a = x525_lb2_0_io_rPort_12_output_0; // @[Math.scala 151:17:@49881.4]
  assign x954_x25_1_io_b = _T_2969[7:0]; // @[Math.scala 152:17:@49882.4]
  assign x955_x26_1_io_a = _T_2973[7:0]; // @[Math.scala 151:17:@49891.4]
  assign x955_x26_1_io_b = x525_lb2_0_io_rPort_0_output_0; // @[Math.scala 152:17:@49892.4]
  assign x956_sum_1_io_a = x954_x25_1_io_result; // @[Math.scala 151:17:@49901.4]
  assign x956_sum_1_io_b = x955_x26_1_io_result; // @[Math.scala 152:17:@49902.4]
  assign x957_div_1_clock = clock; // @[:@49911.4]
  assign x957_div_1_reset = reset; // @[:@49912.4]
  assign x957_div_1_io_a = x956_sum_1_io_result; // @[Math.scala 328:17:@49913.4]
  assign x957_div_1_io_flow = io_in_x512_TREADY; // @[Math.scala 330:20:@49915.4]
  assign x960_x25_1_io_a = x525_lb2_0_io_rPort_3_output_0; // @[Math.scala 151:17:@49933.4]
  assign x960_x25_1_io_b = _T_2993[7:0]; // @[Math.scala 152:17:@49934.4]
  assign x961_x26_1_io_a = _T_2997[7:0]; // @[Math.scala 151:17:@49943.4]
  assign x961_x26_1_io_b = x525_lb2_0_io_rPort_9_output_0; // @[Math.scala 152:17:@49944.4]
  assign x962_sum_1_io_a = x960_x25_1_io_result; // @[Math.scala 151:17:@49953.4]
  assign x962_sum_1_io_b = x961_x26_1_io_result; // @[Math.scala 152:17:@49954.4]
  assign x963_div_1_clock = clock; // @[:@49963.4]
  assign x963_div_1_reset = reset; // @[:@49964.4]
  assign x963_div_1_io_a = x962_sum_1_io_result; // @[Math.scala 328:17:@49965.4]
  assign x963_div_1_io_flow = io_in_x512_TREADY; // @[Math.scala 330:20:@49967.4]
  assign x966_x25_1_io_a = x525_lb2_0_io_rPort_10_output_0; // @[Math.scala 151:17:@49987.4]
  assign x966_x25_1_io_b = _T_3017[7:0]; // @[Math.scala 152:17:@49988.4]
  assign x967_x26_1_io_a = _T_3023[7:0]; // @[Math.scala 151:17:@49997.4]
  assign x967_x26_1_io_b = x525_lb2_0_io_rPort_1_output_0; // @[Math.scala 152:17:@49998.4]
  assign x968_sum_1_io_a = x966_x25_1_io_result; // @[Math.scala 151:17:@50007.4]
  assign x968_sum_1_io_b = x967_x26_1_io_result; // @[Math.scala 152:17:@50008.4]
  assign x969_div_1_clock = clock; // @[:@50017.4]
  assign x969_div_1_reset = reset; // @[:@50018.4]
  assign x969_div_1_io_a = x968_sum_1_io_result; // @[Math.scala 328:17:@50019.4]
  assign x969_div_1_io_flow = io_in_x512_TREADY; // @[Math.scala 330:20:@50021.4]
  assign x971_x25_1_io_a = x525_lb2_0_io_rPort_7_output_0; // @[Math.scala 151:17:@50034.4]
  assign x971_x25_1_io_b = _T_2973[7:0]; // @[Math.scala 152:17:@50035.4]
  assign x972_x26_1_io_a = _T_3043[7:0]; // @[Math.scala 151:17:@50044.4]
  assign x972_x26_1_io_b = x525_lb2_0_io_rPort_6_output_0; // @[Math.scala 152:17:@50045.4]
  assign x973_sum_1_io_a = x971_x25_1_io_result; // @[Math.scala 151:17:@50054.4]
  assign x973_sum_1_io_b = x972_x26_1_io_result; // @[Math.scala 152:17:@50055.4]
  assign x974_div_1_clock = clock; // @[:@50064.4]
  assign x974_div_1_reset = reset; // @[:@50065.4]
  assign x974_div_1_io_a = x973_sum_1_io_result; // @[Math.scala 328:17:@50066.4]
  assign x974_div_1_io_flow = io_in_x512_TREADY; // @[Math.scala 330:20:@50068.4]
  assign x976_x25_1_io_a = x525_lb2_0_io_rPort_13_output_0; // @[Math.scala 151:17:@50081.4]
  assign x976_x25_1_io_b = _T_2997[7:0]; // @[Math.scala 152:17:@50082.4]
  assign x977_x26_1_io_a = _T_3063[7:0]; // @[Math.scala 151:17:@50091.4]
  assign x977_x26_1_io_b = x525_lb2_0_io_rPort_14_output_0; // @[Math.scala 152:17:@50092.4]
  assign x978_sum_1_io_a = x976_x25_1_io_result; // @[Math.scala 151:17:@50101.4]
  assign x978_sum_1_io_b = x977_x26_1_io_result; // @[Math.scala 152:17:@50102.4]
  assign x979_div_1_clock = clock; // @[:@50111.4]
  assign x979_div_1_reset = reset; // @[:@50112.4]
  assign x979_div_1_io_a = x978_sum_1_io_result; // @[Math.scala 328:17:@50113.4]
  assign x979_div_1_io_flow = io_in_x512_TREADY; // @[Math.scala 330:20:@50115.4]
  assign x981_x25_1_io_a = x525_lb2_0_io_rPort_0_output_0; // @[Math.scala 151:17:@50128.4]
  assign x981_x25_1_io_b = _T_3023[7:0]; // @[Math.scala 152:17:@50129.4]
  assign x982_x26_1_io_a = _T_3083[7:0]; // @[Math.scala 151:17:@50138.4]
  assign x982_x26_1_io_b = x525_lb2_0_io_rPort_4_output_0; // @[Math.scala 152:17:@50139.4]
  assign x983_sum_1_io_a = x981_x25_1_io_result; // @[Math.scala 151:17:@50148.4]
  assign x983_sum_1_io_b = x982_x26_1_io_result; // @[Math.scala 152:17:@50149.4]
  assign x984_div_1_clock = clock; // @[:@50158.4]
  assign x984_div_1_reset = reset; // @[:@50159.4]
  assign x984_div_1_io_a = x983_sum_1_io_result; // @[Math.scala 328:17:@50160.4]
  assign x984_div_1_io_flow = io_in_x512_TREADY; // @[Math.scala 330:20:@50162.4]
  assign x987_x25_1_io_a = x525_lb2_0_io_rPort_9_output_0; // @[Math.scala 151:17:@50180.4]
  assign x987_x25_1_io_b = _T_3103[7:0]; // @[Math.scala 152:17:@50181.4]
  assign x988_x26_1_io_a = _T_3107[7:0]; // @[Math.scala 151:17:@50190.4]
  assign x988_x26_1_io_b = x525_lb2_0_io_rPort_11_output_0; // @[Math.scala 152:17:@50191.4]
  assign x989_sum_1_io_a = x987_x25_1_io_result; // @[Math.scala 151:17:@50200.4]
  assign x989_sum_1_io_b = x988_x26_1_io_result; // @[Math.scala 152:17:@50201.4]
  assign x990_div_1_clock = clock; // @[:@50210.4]
  assign x990_div_1_reset = reset; // @[:@50211.4]
  assign x990_div_1_io_a = x989_sum_1_io_result; // @[Math.scala 328:17:@50212.4]
  assign x990_div_1_io_flow = io_in_x512_TREADY; // @[Math.scala 330:20:@50214.4]
  assign RetimeWrapper_194_clock = clock; // @[:@50238.4]
  assign RetimeWrapper_194_reset = reset; // @[:@50239.4]
  assign RetimeWrapper_194_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@50241.4]
  assign RetimeWrapper_194_io_in = {_T_3144,_T_3141}; // @[package.scala 94:16:@50240.4]
  assign RetimeWrapper_195_clock = clock; // @[:@50247.4]
  assign RetimeWrapper_195_reset = reset; // @[:@50248.4]
  assign RetimeWrapper_195_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@50250.4]
  assign RetimeWrapper_195_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@50249.4]
  assign RetimeWrapper_196_clock = clock; // @[:@50256.4]
  assign RetimeWrapper_196_reset = reset; // @[:@50257.4]
  assign RetimeWrapper_196_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@50259.4]
  assign RetimeWrapper_196_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@50258.4]
  assign RetimeWrapper_197_clock = clock; // @[:@50265.4]
  assign RetimeWrapper_197_reset = reset; // @[:@50266.4]
  assign RetimeWrapper_197_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@50268.4]
  assign RetimeWrapper_197_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@50267.4]
endmodule
module x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1( // @[:@50286.2]
  input          clock, // @[:@50287.4]
  input          reset, // @[:@50288.4]
  input          io_in_x511_TVALID, // @[:@50289.4]
  output         io_in_x511_TREADY, // @[:@50289.4]
  input  [255:0] io_in_x511_TDATA, // @[:@50289.4]
  input  [7:0]   io_in_x511_TID, // @[:@50289.4]
  input  [7:0]   io_in_x511_TDEST, // @[:@50289.4]
  output         io_in_x512_TVALID, // @[:@50289.4]
  input          io_in_x512_TREADY, // @[:@50289.4]
  output [255:0] io_in_x512_TDATA, // @[:@50289.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@50289.4]
  input          io_sigsIn_smChildAcks_0, // @[:@50289.4]
  output         io_sigsOut_smDoneIn_0, // @[:@50289.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@50289.4]
  input          io_rr // @[:@50289.4]
);
  wire  x519_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@50299.4]
  wire  x519_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@50299.4]
  wire  x519_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@50299.4]
  wire  x519_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@50299.4]
  wire [31:0] x519_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@50299.4]
  wire [31:0] x519_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@50299.4]
  wire  x519_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@50299.4]
  wire  x519_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@50299.4]
  wire  x519_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@50299.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 32:18:@50358.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 32:18:@50358.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 32:18:@50358.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 32:18:@50358.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 32:18:@50358.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 32:18:@50358.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 32:18:@50358.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 32:18:@50358.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 32:18:@50358.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 32:18:@50358.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 32:18:@50358.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 32:18:@50358.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@50386.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@50386.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@50386.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@50386.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@50386.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@50428.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@50428.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@50428.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@50428.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@50428.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@50436.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@50436.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@50436.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@50436.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@50436.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x511_TREADY; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire [255:0] x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x511_TDATA; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire [7:0] x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x511_TID; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire [7:0] x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x511_TDEST; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x512_TVALID; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x512_TREADY; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire [255:0] x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x512_TDATA; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire [31:0] x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire [31:0] x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
  wire  _T_239; // @[package.scala 96:25:@50391.4 package.scala 96:25:@50392.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x996_outr_UnitPipe.scala 68:66:@50397.4]
  wire  _T_252; // @[package.scala 96:25:@50433.4 package.scala 96:25:@50434.4]
  wire  _T_258; // @[package.scala 96:25:@50441.4 package.scala 96:25:@50442.4]
  wire  _T_261; // @[SpatialBlocks.scala 110:93:@50444.4]
  wire  x995_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 110:90:@50445.4]
  wire  _T_263; // @[SpatialBlocks.scala 128:36:@50453.4]
  wire  _T_264; // @[SpatialBlocks.scala 128:78:@50454.4]
  wire  _T_269; // @[SpatialBlocks.scala 130:61:@50463.4]
  x519_ctrchain x519_ctrchain ( // @[SpatialBlocks.scala 37:22:@50299.4]
    .clock(x519_ctrchain_clock),
    .reset(x519_ctrchain_reset),
    .io_input_reset(x519_ctrchain_io_input_reset),
    .io_input_enable(x519_ctrchain_io_input_enable),
    .io_output_counts_1(x519_ctrchain_io_output_counts_1),
    .io_output_counts_0(x519_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x519_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x519_ctrchain_io_output_oobs_1),
    .io_output_done(x519_ctrchain_io_output_done)
  );
  x995_inr_Foreach_SAMPLER_BOX_sm x995_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 32:18:@50358.4]
    .clock(x995_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x995_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x995_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x995_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x995_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x995_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x995_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x995_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x995_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x995_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x995_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x995_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@50386.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@50428.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@50436.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1 x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1362:24:@50468.4]
    .clock(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x511_TREADY(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x511_TREADY),
    .io_in_x511_TDATA(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x511_TDATA),
    .io_in_x511_TID(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x511_TID),
    .io_in_x511_TDEST(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x511_TDEST),
    .io_in_x512_TVALID(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x512_TVALID),
    .io_in_x512_TREADY(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x512_TREADY),
    .io_in_x512_TDATA(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x512_TDATA),
    .io_sigsIn_backpressure(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_239 = RetimeWrapper_io_out; // @[package.scala 96:25:@50391.4 package.scala 96:25:@50392.4]
  assign x995_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x511_TVALID | x995_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x996_outr_UnitPipe.scala 68:66:@50397.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@50433.4 package.scala 96:25:@50434.4]
  assign _T_258 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@50441.4 package.scala 96:25:@50442.4]
  assign _T_261 = ~ _T_258; // @[SpatialBlocks.scala 110:93:@50444.4]
  assign x995_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_252 & _T_261; // @[SpatialBlocks.scala 110:90:@50445.4]
  assign _T_263 = x995_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@50453.4]
  assign _T_264 = ~ x995_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@50454.4]
  assign _T_269 = x995_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 130:61:@50463.4]
  assign io_in_x511_TREADY = x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x511_TREADY; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 48:23:@50525.4]
  assign io_in_x512_TVALID = x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x512_TVALID; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 49:23:@50535.4]
  assign io_in_x512_TDATA = x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x512_TDATA; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 49:23:@50533.4]
  assign io_sigsOut_smDoneIn_0 = x995_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 127:53:@50451.4]
  assign io_sigsOut_smCtrCopyDone_0 = x995_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 139:125:@50467.4]
  assign x519_ctrchain_clock = clock; // @[:@50300.4]
  assign x519_ctrchain_reset = reset; // @[:@50301.4]
  assign x519_ctrchain_io_input_reset = x995_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@50466.4]
  assign x519_ctrchain_io_input_enable = _T_269 & x995_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 104:75:@50421.4 SpatialBlocks.scala 130:45:@50465.4]
  assign x995_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@50359.4]
  assign x995_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@50360.4]
  assign x995_inr_Foreach_SAMPLER_BOX_sm_io_enable = x995_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x995_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 112:18:@50448.4]
  assign x995_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_239 : 1'h0; // @[sm_x996_outr_UnitPipe.scala 66:50:@50394.4]
  assign x995_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@50450.4]
  assign x995_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x512_TREADY | x995_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 105:24:@50422.4]
  assign x995_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x996_outr_UnitPipe.scala 70:48:@50400.4]
  assign RetimeWrapper_clock = clock; // @[:@50387.4]
  assign RetimeWrapper_reset = reset; // @[:@50388.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@50390.4]
  assign RetimeWrapper_io_in = x519_ctrchain_io_output_done; // @[package.scala 94:16:@50389.4]
  assign RetimeWrapper_1_clock = clock; // @[:@50429.4]
  assign RetimeWrapper_1_reset = reset; // @[:@50430.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@50432.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@50431.4]
  assign RetimeWrapper_2_clock = clock; // @[:@50437.4]
  assign RetimeWrapper_2_reset = reset; // @[:@50438.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@50440.4]
  assign RetimeWrapper_2_io_in = x995_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@50439.4]
  assign x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@50469.4]
  assign x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@50470.4]
  assign x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x511_TDATA = io_in_x511_TDATA; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 48:23:@50524.4]
  assign x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x511_TID = io_in_x511_TID; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 48:23:@50520.4]
  assign x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x511_TDEST = io_in_x511_TDEST; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 48:23:@50519.4]
  assign x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x512_TREADY = io_in_x512_TREADY; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 49:23:@50534.4]
  assign x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x512_TREADY | x995_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1366:22:@50552.4]
  assign x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_263 & _T_264; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1366:22:@50550.4]
  assign x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x995_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1366:22:@50548.4]
  assign x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = x519_ctrchain_io_output_counts_1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1366:22:@50543.4]
  assign x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x519_ctrchain_io_output_counts_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1366:22:@50542.4]
  assign x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x519_ctrchain_io_output_oobs_0; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1366:22:@50540.4]
  assign x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x519_ctrchain_io_output_oobs_1; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1366:22:@50541.4]
  assign x995_inr_Foreach_SAMPLER_BOX_kernelx995_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x995_inr_Foreach_SAMPLER_BOX.scala 1365:18:@50536.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@50565.2]
  input          clock, // @[:@50566.4]
  input          reset, // @[:@50567.4]
  input          io_in_x511_TVALID, // @[:@50568.4]
  output         io_in_x511_TREADY, // @[:@50568.4]
  input  [255:0] io_in_x511_TDATA, // @[:@50568.4]
  input  [7:0]   io_in_x511_TID, // @[:@50568.4]
  input  [7:0]   io_in_x511_TDEST, // @[:@50568.4]
  output         io_in_x512_TVALID, // @[:@50568.4]
  input          io_in_x512_TREADY, // @[:@50568.4]
  output [255:0] io_in_x512_TDATA, // @[:@50568.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@50568.4]
  input          io_sigsIn_smChildAcks_0, // @[:@50568.4]
  output         io_sigsOut_smDoneIn_0, // @[:@50568.4]
  input          io_rr // @[:@50568.4]
);
  wire  x996_outr_UnitPipe_sm_clock; // @[sm_x996_outr_UnitPipe.scala 32:18:@50709.4]
  wire  x996_outr_UnitPipe_sm_reset; // @[sm_x996_outr_UnitPipe.scala 32:18:@50709.4]
  wire  x996_outr_UnitPipe_sm_io_enable; // @[sm_x996_outr_UnitPipe.scala 32:18:@50709.4]
  wire  x996_outr_UnitPipe_sm_io_done; // @[sm_x996_outr_UnitPipe.scala 32:18:@50709.4]
  wire  x996_outr_UnitPipe_sm_io_parentAck; // @[sm_x996_outr_UnitPipe.scala 32:18:@50709.4]
  wire  x996_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x996_outr_UnitPipe.scala 32:18:@50709.4]
  wire  x996_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x996_outr_UnitPipe.scala 32:18:@50709.4]
  wire  x996_outr_UnitPipe_sm_io_childAck_0; // @[sm_x996_outr_UnitPipe.scala 32:18:@50709.4]
  wire  x996_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x996_outr_UnitPipe.scala 32:18:@50709.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@50761.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@50761.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@50761.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@50761.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@50761.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@50769.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@50769.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@50769.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@50769.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@50769.4]
  wire  x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_clock; // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
  wire  x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_reset; // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
  wire  x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x511_TVALID; // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
  wire  x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x511_TREADY; // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
  wire [255:0] x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x511_TDATA; // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
  wire [7:0] x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x511_TID; // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
  wire [7:0] x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x511_TDEST; // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
  wire  x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x512_TVALID; // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
  wire  x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x512_TREADY; // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
  wire [255:0] x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x512_TDATA; // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
  wire  x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
  wire  x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
  wire  x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
  wire  x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
  wire  x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_rr; // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
  wire  _T_246; // @[package.scala 96:25:@50766.4 package.scala 96:25:@50767.4]
  wire  _T_252; // @[package.scala 96:25:@50774.4 package.scala 96:25:@50775.4]
  wire  _T_255; // @[SpatialBlocks.scala 110:93:@50777.4]
  x996_outr_UnitPipe_sm x996_outr_UnitPipe_sm ( // @[sm_x996_outr_UnitPipe.scala 32:18:@50709.4]
    .clock(x996_outr_UnitPipe_sm_clock),
    .reset(x996_outr_UnitPipe_sm_reset),
    .io_enable(x996_outr_UnitPipe_sm_io_enable),
    .io_done(x996_outr_UnitPipe_sm_io_done),
    .io_parentAck(x996_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x996_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x996_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x996_outr_UnitPipe_sm_io_childAck_0),
    .io_ctrCopyDone_0(x996_outr_UnitPipe_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@50761.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@50769.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1 x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1 ( // @[sm_x996_outr_UnitPipe.scala 75:24:@50796.4]
    .clock(x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_clock),
    .reset(x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_reset),
    .io_in_x511_TVALID(x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x511_TVALID),
    .io_in_x511_TREADY(x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x511_TREADY),
    .io_in_x511_TDATA(x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x511_TDATA),
    .io_in_x511_TID(x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x511_TID),
    .io_in_x511_TDEST(x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x511_TDEST),
    .io_in_x512_TVALID(x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x512_TVALID),
    .io_in_x512_TREADY(x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x512_TREADY),
    .io_in_x512_TDATA(x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x512_TDATA),
    .io_sigsIn_smEnableOuts_0(x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_246 = RetimeWrapper_io_out; // @[package.scala 96:25:@50766.4 package.scala 96:25:@50767.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@50774.4 package.scala 96:25:@50775.4]
  assign _T_255 = ~ _T_252; // @[SpatialBlocks.scala 110:93:@50777.4]
  assign io_in_x511_TREADY = x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x511_TREADY; // @[sm_x996_outr_UnitPipe.scala 48:23:@50851.4]
  assign io_in_x512_TVALID = x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x512_TVALID; // @[sm_x996_outr_UnitPipe.scala 49:23:@50861.4]
  assign io_in_x512_TDATA = x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x512_TDATA; // @[sm_x996_outr_UnitPipe.scala 49:23:@50859.4]
  assign io_sigsOut_smDoneIn_0 = x996_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@50784.4]
  assign x996_outr_UnitPipe_sm_clock = clock; // @[:@50710.4]
  assign x996_outr_UnitPipe_sm_reset = reset; // @[:@50711.4]
  assign x996_outr_UnitPipe_sm_io_enable = _T_246 & _T_255; // @[SpatialBlocks.scala 112:18:@50781.4]
  assign x996_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@50783.4]
  assign x996_outr_UnitPipe_sm_io_doneIn_0 = x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@50753.4]
  assign x996_outr_UnitPipe_sm_io_ctrCopyDone_0 = x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 132:80:@50795.4]
  assign RetimeWrapper_clock = clock; // @[:@50762.4]
  assign RetimeWrapper_reset = reset; // @[:@50763.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@50765.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@50764.4]
  assign RetimeWrapper_1_clock = clock; // @[:@50770.4]
  assign RetimeWrapper_1_reset = reset; // @[:@50771.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@50773.4]
  assign RetimeWrapper_1_io_in = x996_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@50772.4]
  assign x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_clock = clock; // @[:@50797.4]
  assign x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_reset = reset; // @[:@50798.4]
  assign x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x511_TVALID = io_in_x511_TVALID; // @[sm_x996_outr_UnitPipe.scala 48:23:@50852.4]
  assign x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x511_TDATA = io_in_x511_TDATA; // @[sm_x996_outr_UnitPipe.scala 48:23:@50850.4]
  assign x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x511_TID = io_in_x511_TID; // @[sm_x996_outr_UnitPipe.scala 48:23:@50846.4]
  assign x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x511_TDEST = io_in_x511_TDEST; // @[sm_x996_outr_UnitPipe.scala 48:23:@50845.4]
  assign x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_in_x512_TREADY = io_in_x512_TREADY; // @[sm_x996_outr_UnitPipe.scala 49:23:@50860.4]
  assign x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x996_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x996_outr_UnitPipe.scala 79:22:@50870.4]
  assign x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x996_outr_UnitPipe_sm_io_childAck_0; // @[sm_x996_outr_UnitPipe.scala 79:22:@50868.4]
  assign x996_outr_UnitPipe_kernelx996_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x996_outr_UnitPipe.scala 78:18:@50862.4]
endmodule
module AccelUnit( // @[:@50889.2]
  input          clock, // @[:@50890.4]
  input          reset, // @[:@50891.4]
  input          io_enable, // @[:@50892.4]
  output         io_done, // @[:@50892.4]
  input          io_reset, // @[:@50892.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@50892.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@50892.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@50892.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@50892.4]
  output         io_memStreams_loads_0_data_ready, // @[:@50892.4]
  input          io_memStreams_loads_0_data_valid, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@50892.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@50892.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@50892.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@50892.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@50892.4]
  input          io_memStreams_stores_0_data_ready, // @[:@50892.4]
  output         io_memStreams_stores_0_data_valid, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_1, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_2, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_3, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_4, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_5, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_6, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_7, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_8, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_9, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_10, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_11, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_12, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_13, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_14, // @[:@50892.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_15, // @[:@50892.4]
  output [15:0]  io_memStreams_stores_0_data_bits_wstrb, // @[:@50892.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@50892.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@50892.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@50892.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@50892.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@50892.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@50892.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@50892.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@50892.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@50892.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@50892.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@50892.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@50892.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@50892.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@50892.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@50892.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@50892.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@50892.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@50892.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@50892.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@50892.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@50892.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@50892.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@50892.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@50892.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@50892.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@50892.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@50892.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@50892.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@50892.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@50892.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@50892.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@50892.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@50892.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@50892.4]
  output         io_heap_0_req_valid, // @[:@50892.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@50892.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@50892.4]
  input          io_heap_0_resp_valid, // @[:@50892.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@50892.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@50892.4]
  input  [63:0]  io_argIns_0, // @[:@50892.4]
  input  [63:0]  io_argIns_1, // @[:@50892.4]
  input          io_argOuts_0_port_ready, // @[:@50892.4]
  output         io_argOuts_0_port_valid, // @[:@50892.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@50892.4]
  input  [63:0]  io_argOuts_0_echo // @[:@50892.4]
);
  wire  SingleCounter_clock; // @[Main.scala 35:32:@51055.4]
  wire  SingleCounter_reset; // @[Main.scala 35:32:@51055.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 35:32:@51055.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 35:32:@51055.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@51073.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@51073.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@51073.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@51073.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@51073.4]
  wire  SRFF_clock; // @[Main.scala 39:28:@51082.4]
  wire  SRFF_reset; // @[Main.scala 39:28:@51082.4]
  wire  SRFF_io_input_set; // @[Main.scala 39:28:@51082.4]
  wire  SRFF_io_input_reset; // @[Main.scala 39:28:@51082.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 39:28:@51082.4]
  wire  SRFF_io_output; // @[Main.scala 39:28:@51082.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@51120.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@51120.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@51120.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@51120.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@51120.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@51120.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@51120.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 32:18:@51120.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 32:18:@51120.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 32:18:@51120.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@51152.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@51152.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@51152.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@51152.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@51152.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 73:24:@51211.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 73:24:@51211.4]
  wire  RootController_kernelRootController_concrete1_io_in_x511_TVALID; // @[sm_RootController.scala 73:24:@51211.4]
  wire  RootController_kernelRootController_concrete1_io_in_x511_TREADY; // @[sm_RootController.scala 73:24:@51211.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x511_TDATA; // @[sm_RootController.scala 73:24:@51211.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x511_TID; // @[sm_RootController.scala 73:24:@51211.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x511_TDEST; // @[sm_RootController.scala 73:24:@51211.4]
  wire  RootController_kernelRootController_concrete1_io_in_x512_TVALID; // @[sm_RootController.scala 73:24:@51211.4]
  wire  RootController_kernelRootController_concrete1_io_in_x512_TREADY; // @[sm_RootController.scala 73:24:@51211.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x512_TDATA; // @[sm_RootController.scala 73:24:@51211.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 73:24:@51211.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 73:24:@51211.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 73:24:@51211.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 73:24:@51211.4]
  wire  _T_599; // @[package.scala 96:25:@51078.4 package.scala 96:25:@51079.4]
  wire  _T_664; // @[Main.scala 41:50:@51148.4]
  wire  _T_665; // @[Main.scala 41:59:@51149.4]
  wire  _T_677; // @[package.scala 100:49:@51169.4]
  reg  _T_680; // @[package.scala 48:56:@51170.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 35:32:@51055.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@51073.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 39:28:@51082.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@51120.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@51152.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 73:24:@51211.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x511_TVALID(RootController_kernelRootController_concrete1_io_in_x511_TVALID),
    .io_in_x511_TREADY(RootController_kernelRootController_concrete1_io_in_x511_TREADY),
    .io_in_x511_TDATA(RootController_kernelRootController_concrete1_io_in_x511_TDATA),
    .io_in_x511_TID(RootController_kernelRootController_concrete1_io_in_x511_TID),
    .io_in_x511_TDEST(RootController_kernelRootController_concrete1_io_in_x511_TDEST),
    .io_in_x512_TVALID(RootController_kernelRootController_concrete1_io_in_x512_TVALID),
    .io_in_x512_TREADY(RootController_kernelRootController_concrete1_io_in_x512_TREADY),
    .io_in_x512_TDATA(RootController_kernelRootController_concrete1_io_in_x512_TDATA),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@51078.4 package.scala 96:25:@51079.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 41:50:@51148.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 41:59:@51149.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@51169.4]
  assign io_done = SRFF_io_output; // @[Main.scala 48:23:@51168.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x511_TREADY; // @[sm_RootController.scala 48:23:@51266.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x512_TVALID; // @[sm_RootController.scala 49:23:@51276.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x512_TDATA; // @[sm_RootController.scala 49:23:@51274.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 49:23:@51273.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 49:23:@51272.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 49:23:@51271.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 49:23:@51270.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 49:23:@51269.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 49:23:@51268.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@51056.4]
  assign SingleCounter_reset = reset; // @[:@51057.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 36:79:@51071.4]
  assign RetimeWrapper_clock = clock; // @[:@51074.4]
  assign RetimeWrapper_reset = reset; // @[:@51075.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@51077.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@51076.4]
  assign SRFF_clock = clock; // @[:@51083.4]
  assign SRFF_reset = reset; // @[:@51084.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 57:29:@51303.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 46:31:@51166.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 47:36:@51167.4]
  assign RootController_sm_clock = clock; // @[:@51121.4]
  assign RootController_sm_reset = reset; // @[:@51122.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 45:33:@51165.4 SpatialBlocks.scala 112:18:@51199.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 106:15:@51193.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 49:34:@51173.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@51190.4]
  assign RetimeWrapper_1_clock = clock; // @[:@51153.4]
  assign RetimeWrapper_1_reset = reset; // @[:@51154.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@51156.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@51155.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@51212.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@51213.4]
  assign RootController_kernelRootController_concrete1_io_in_x511_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 48:23:@51267.4]
  assign RootController_kernelRootController_concrete1_io_in_x511_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 48:23:@51265.4]
  assign RootController_kernelRootController_concrete1_io_in_x511_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 48:23:@51261.4]
  assign RootController_kernelRootController_concrete1_io_in_x511_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 48:23:@51260.4]
  assign RootController_kernelRootController_concrete1_io_in_x512_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 49:23:@51275.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 77:22:@51285.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 77:22:@51283.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 76:18:@51277.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module SpatialIP( // @[:@51305.2]
  input         clock, // @[:@51306.4]
  input         reset, // @[:@51307.4]
  input  [31:0] io_raddr, // @[:@51308.4]
  input         io_wen, // @[:@51308.4]
  input  [31:0] io_waddr, // @[:@51308.4]
  input  [63:0] io_wdata, // @[:@51308.4]
  output [63:0] io_rdata // @[:@51308.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 53:44:@51310.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@51310.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@51310.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@51310.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@51310.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@51310.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@51310.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@51310.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@51310.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@51310.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@51310.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@51310.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  assign io_rdata = 64'h0;
  assign accel_clock = clock; // @[:@51311.4]
  assign accel_reset = reset; // @[:@51312.4]
  assign accel_io_enable = 1'h0;
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_loads_0_data_valid = 1'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0;
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_stores_0_data_ready = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0;
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0;
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0;
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0;
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = 1'h0;
  assign accel_io_heap_0_resp_bits_allocDealloc = 1'h0;
  assign accel_io_heap_0_resp_bits_sizeAddr = 64'h0;
  assign accel_io_argIns_0 = 64'h0;
  assign accel_io_argIns_1 = 64'h0;
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0;
endmodule
