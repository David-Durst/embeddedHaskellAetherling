module FIFO(
  input        clock,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_1_0_0,
  input  [7:0] I_2_0_0,
  input  [7:0] I_3_0_0,
  input  [7:0] I_4_0_0,
  input  [7:0] I_5_0_0,
  input  [7:0] I_6_0_0,
  input  [7:0] I_7_0_0,
  input  [7:0] I_8_0_0,
  input  [7:0] I_9_0_0,
  input  [7:0] I_10_0_0,
  input  [7:0] I_11_0_0,
  input  [7:0] I_12_0_0,
  input  [7:0] I_13_0_0,
  input  [7:0] I_14_0_0,
  input  [7:0] I_15_0_0,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0,
  output [7:0] O_8_0_0,
  output [7:0] O_9_0_0,
  output [7:0] O_10_0_0,
  output [7:0] O_11_0_0,
  output [7:0] O_12_0_0,
  output [7:0] O_13_0_0,
  output [7:0] O_14_0_0,
  output [7:0] O_15_0_0
);
  reg [7:0] _T__0_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [7:0] _T__1_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg [7:0] _T__2_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg [7:0] _T__3_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg [7:0] _T__4_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_4;
  reg [7:0] _T__5_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_5;
  reg [7:0] _T__6_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_6;
  reg [7:0] _T__7_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_7;
  reg [7:0] _T__8_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_8;
  reg [7:0] _T__9_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_9;
  reg [7:0] _T__10_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_10;
  reg [7:0] _T__11_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_11;
  reg [7:0] _T__12_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_12;
  reg [7:0] _T__13_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_13;
  reg [7:0] _T__14_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_14;
  reg [7:0] _T__15_0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_15;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_16;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0_0_0 = _T__0_0_0; // @[FIFO.scala 14:7]
  assign O_1_0_0 = _T__1_0_0; // @[FIFO.scala 14:7]
  assign O_2_0_0 = _T__2_0_0; // @[FIFO.scala 14:7]
  assign O_3_0_0 = _T__3_0_0; // @[FIFO.scala 14:7]
  assign O_4_0_0 = _T__4_0_0; // @[FIFO.scala 14:7]
  assign O_5_0_0 = _T__5_0_0; // @[FIFO.scala 14:7]
  assign O_6_0_0 = _T__6_0_0; // @[FIFO.scala 14:7]
  assign O_7_0_0 = _T__7_0_0; // @[FIFO.scala 14:7]
  assign O_8_0_0 = _T__8_0_0; // @[FIFO.scala 14:7]
  assign O_9_0_0 = _T__9_0_0; // @[FIFO.scala 14:7]
  assign O_10_0_0 = _T__10_0_0; // @[FIFO.scala 14:7]
  assign O_11_0_0 = _T__11_0_0; // @[FIFO.scala 14:7]
  assign O_12_0_0 = _T__12_0_0; // @[FIFO.scala 14:7]
  assign O_13_0_0 = _T__13_0_0; // @[FIFO.scala 14:7]
  assign O_14_0_0 = _T__14_0_0; // @[FIFO.scala 14:7]
  assign O_15_0_0 = _T__15_0_0; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0_0_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__1_0_0 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__2_0_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__3_0_0 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T__4_0_0 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T__5_0_0 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__6_0_0 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__7_0_0 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T__8_0_0 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T__9_0_0 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__10_0_0 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__11_0_0 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T__12_0_0 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T__13_0_0 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__14_0_0 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__15_0_0 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0_0_0 <= I_0_0_0;
    _T__1_0_0 <= I_1_0_0;
    _T__2_0_0 <= I_2_0_0;
    _T__3_0_0 <= I_3_0_0;
    _T__4_0_0 <= I_4_0_0;
    _T__5_0_0 <= I_5_0_0;
    _T__6_0_0 <= I_6_0_0;
    _T__7_0_0 <= I_7_0_0;
    _T__8_0_0 <= I_8_0_0;
    _T__9_0_0 <= I_9_0_0;
    _T__10_0_0 <= I_10_0_0;
    _T__11_0_0 <= I_11_0_0;
    _T__12_0_0 <= I_12_0_0;
    _T__13_0_0 <= I_13_0_0;
    _T__14_0_0 <= I_14_0_0;
    _T__15_0_0 <= I_15_0_0;
    _T_1 <= valid_up;
  end
endmodule
module NestedCounters(
  input   CE,
  output  valid
);
  assign valid = CE; // @[NestedCounters.scala 65:13]
endmodule
module NestedCounters_1(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 53:31]
  wire  NestedCounters_valid; // @[NestedCounters.scala 53:31]
  NestedCounters NestedCounters ( // @[NestedCounters.scala 53:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 56:11]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 57:22]
endmodule
module NestedCounters_2(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 53:31]
  wire  NestedCounters_valid; // @[NestedCounters.scala 53:31]
  NestedCounters_1 NestedCounters ( // @[NestedCounters.scala 53:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 56:11]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 57:22]
endmodule
module NestedCountersWithNumValid(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 20:44]
  wire  NestedCounters_valid; // @[NestedCounters.scala 20:44]
  NestedCounters_2 NestedCounters ( // @[NestedCounters.scala 20:44]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 22:9]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 21:27]
endmodule
module RAM_ST(
  input        clock,
  input        RE,
  input  [6:0] RADDR,
  output [7:0] RDATA_0_0,
  input        WE,
  input  [6:0] WADDR,
  input  [7:0] WDATA_0_0
);
  wire  write_elem_counter_CE; // @[RAM_ST.scala 20:34]
  wire  write_elem_counter_valid; // @[RAM_ST.scala 20:34]
  wire  read_elem_counter_CE; // @[RAM_ST.scala 21:33]
  wire  read_elem_counter_valid; // @[RAM_ST.scala 21:33]
  reg [7:0] ram_0_0 [0:119]; // @[RAM_ST.scala 29:24]
  reg [31:0] _RAND_0;
  wire [7:0] ram_0_0__T_8_data; // @[RAM_ST.scala 29:24]
  wire [6:0] ram_0_0__T_8_addr; // @[RAM_ST.scala 29:24]
  reg [31:0] _RAND_1;
  wire [7:0] ram_0_0__T_2_data; // @[RAM_ST.scala 29:24]
  wire [6:0] ram_0_0__T_2_addr; // @[RAM_ST.scala 29:24]
  wire  ram_0_0__T_2_mask; // @[RAM_ST.scala 29:24]
  wire  ram_0_0__T_2_en; // @[RAM_ST.scala 29:24]
  reg  ram_0_0__T_8_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [6:0] ram_0_0__T_8_addr_pipe_0;
  reg [31:0] _RAND_3;
  wire [6:0] _GEN_1; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_2; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_3; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_4; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_5; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_6; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_7; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_8; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_9; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_10; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_11; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_12; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_13; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_14; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_15; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_16; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_17; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_18; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_19; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_20; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_21; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_22; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_23; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_24; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_25; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_26; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_27; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_28; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_29; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_30; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_31; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_32; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_33; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_34; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_35; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_36; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_37; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_38; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_39; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_40; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_41; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_42; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_43; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_44; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_45; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_46; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_47; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_48; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_49; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_50; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_51; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_52; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_53; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_54; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_55; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_56; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_57; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_58; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_59; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_60; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_61; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_62; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_63; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_64; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_65; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_66; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_67; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_68; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_69; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_70; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_71; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_72; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_73; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_74; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_75; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_76; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_77; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_78; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_79; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_80; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_81; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_82; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_83; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_84; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_85; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_86; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_87; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_88; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_89; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_90; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_91; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_92; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_93; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_94; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_95; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_96; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_97; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_98; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_99; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_100; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_101; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_102; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_103; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_104; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_105; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_106; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_107; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_108; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_109; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_110; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_111; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_112; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_113; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_114; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_115; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_116; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_117; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_118; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_119; // @[RAM_ST.scala 31:71]
  wire [7:0] _T; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_126; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_127; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_128; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_129; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_130; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_131; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_132; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_133; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_134; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_135; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_136; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_137; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_138; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_139; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_140; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_141; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_142; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_143; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_144; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_145; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_146; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_147; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_148; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_149; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_150; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_151; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_152; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_153; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_154; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_155; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_156; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_157; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_158; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_159; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_160; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_161; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_162; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_163; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_164; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_165; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_166; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_167; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_168; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_169; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_170; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_171; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_172; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_173; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_174; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_175; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_176; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_177; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_178; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_179; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_180; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_181; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_182; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_183; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_184; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_185; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_186; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_187; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_188; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_189; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_190; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_191; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_192; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_193; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_194; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_195; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_196; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_197; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_198; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_199; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_200; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_201; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_202; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_203; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_204; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_205; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_206; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_207; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_208; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_209; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_210; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_211; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_212; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_213; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_214; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_215; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_216; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_217; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_218; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_219; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_220; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_221; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_222; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_223; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_224; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_225; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_226; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_227; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_228; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_229; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_230; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_231; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_232; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_233; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_234; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_235; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_236; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_237; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_238; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_239; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_240; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_241; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_242; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_243; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_244; // @[RAM_ST.scala 32:46]
  wire [7:0] _T_3; // @[RAM_ST.scala 32:46]
  NestedCountersWithNumValid write_elem_counter ( // @[RAM_ST.scala 20:34]
    .CE(write_elem_counter_CE),
    .valid(write_elem_counter_valid)
  );
  NestedCountersWithNumValid read_elem_counter ( // @[RAM_ST.scala 21:33]
    .CE(read_elem_counter_CE),
    .valid(read_elem_counter_valid)
  );
  assign ram_0_0__T_8_addr = ram_0_0__T_8_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_0_0__T_8_data = ram_0_0[ram_0_0__T_8_addr]; // @[RAM_ST.scala 29:24]
  `else
  assign ram_0_0__T_8_data = ram_0_0__T_8_addr >= 7'h78 ? _RAND_1[7:0] : ram_0_0[ram_0_0__T_8_addr]; // @[RAM_ST.scala 29:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_0_0__T_2_data = WDATA_0_0;
  assign ram_0_0__T_2_addr = _T[6:0];
  assign ram_0_0__T_2_mask = 1'h1;
  assign ram_0_0__T_2_en = write_elem_counter_valid;
  assign _GEN_1 = 7'h1 == WADDR ? 7'h1 : 7'h0; // @[RAM_ST.scala 31:71]
  assign _GEN_2 = 7'h2 == WADDR ? 7'h2 : _GEN_1; // @[RAM_ST.scala 31:71]
  assign _GEN_3 = 7'h3 == WADDR ? 7'h3 : _GEN_2; // @[RAM_ST.scala 31:71]
  assign _GEN_4 = 7'h4 == WADDR ? 7'h4 : _GEN_3; // @[RAM_ST.scala 31:71]
  assign _GEN_5 = 7'h5 == WADDR ? 7'h5 : _GEN_4; // @[RAM_ST.scala 31:71]
  assign _GEN_6 = 7'h6 == WADDR ? 7'h6 : _GEN_5; // @[RAM_ST.scala 31:71]
  assign _GEN_7 = 7'h7 == WADDR ? 7'h7 : _GEN_6; // @[RAM_ST.scala 31:71]
  assign _GEN_8 = 7'h8 == WADDR ? 7'h8 : _GEN_7; // @[RAM_ST.scala 31:71]
  assign _GEN_9 = 7'h9 == WADDR ? 7'h9 : _GEN_8; // @[RAM_ST.scala 31:71]
  assign _GEN_10 = 7'ha == WADDR ? 7'ha : _GEN_9; // @[RAM_ST.scala 31:71]
  assign _GEN_11 = 7'hb == WADDR ? 7'hb : _GEN_10; // @[RAM_ST.scala 31:71]
  assign _GEN_12 = 7'hc == WADDR ? 7'hc : _GEN_11; // @[RAM_ST.scala 31:71]
  assign _GEN_13 = 7'hd == WADDR ? 7'hd : _GEN_12; // @[RAM_ST.scala 31:71]
  assign _GEN_14 = 7'he == WADDR ? 7'he : _GEN_13; // @[RAM_ST.scala 31:71]
  assign _GEN_15 = 7'hf == WADDR ? 7'hf : _GEN_14; // @[RAM_ST.scala 31:71]
  assign _GEN_16 = 7'h10 == WADDR ? 7'h10 : _GEN_15; // @[RAM_ST.scala 31:71]
  assign _GEN_17 = 7'h11 == WADDR ? 7'h11 : _GEN_16; // @[RAM_ST.scala 31:71]
  assign _GEN_18 = 7'h12 == WADDR ? 7'h12 : _GEN_17; // @[RAM_ST.scala 31:71]
  assign _GEN_19 = 7'h13 == WADDR ? 7'h13 : _GEN_18; // @[RAM_ST.scala 31:71]
  assign _GEN_20 = 7'h14 == WADDR ? 7'h14 : _GEN_19; // @[RAM_ST.scala 31:71]
  assign _GEN_21 = 7'h15 == WADDR ? 7'h15 : _GEN_20; // @[RAM_ST.scala 31:71]
  assign _GEN_22 = 7'h16 == WADDR ? 7'h16 : _GEN_21; // @[RAM_ST.scala 31:71]
  assign _GEN_23 = 7'h17 == WADDR ? 7'h17 : _GEN_22; // @[RAM_ST.scala 31:71]
  assign _GEN_24 = 7'h18 == WADDR ? 7'h18 : _GEN_23; // @[RAM_ST.scala 31:71]
  assign _GEN_25 = 7'h19 == WADDR ? 7'h19 : _GEN_24; // @[RAM_ST.scala 31:71]
  assign _GEN_26 = 7'h1a == WADDR ? 7'h1a : _GEN_25; // @[RAM_ST.scala 31:71]
  assign _GEN_27 = 7'h1b == WADDR ? 7'h1b : _GEN_26; // @[RAM_ST.scala 31:71]
  assign _GEN_28 = 7'h1c == WADDR ? 7'h1c : _GEN_27; // @[RAM_ST.scala 31:71]
  assign _GEN_29 = 7'h1d == WADDR ? 7'h1d : _GEN_28; // @[RAM_ST.scala 31:71]
  assign _GEN_30 = 7'h1e == WADDR ? 7'h1e : _GEN_29; // @[RAM_ST.scala 31:71]
  assign _GEN_31 = 7'h1f == WADDR ? 7'h1f : _GEN_30; // @[RAM_ST.scala 31:71]
  assign _GEN_32 = 7'h20 == WADDR ? 7'h20 : _GEN_31; // @[RAM_ST.scala 31:71]
  assign _GEN_33 = 7'h21 == WADDR ? 7'h21 : _GEN_32; // @[RAM_ST.scala 31:71]
  assign _GEN_34 = 7'h22 == WADDR ? 7'h22 : _GEN_33; // @[RAM_ST.scala 31:71]
  assign _GEN_35 = 7'h23 == WADDR ? 7'h23 : _GEN_34; // @[RAM_ST.scala 31:71]
  assign _GEN_36 = 7'h24 == WADDR ? 7'h24 : _GEN_35; // @[RAM_ST.scala 31:71]
  assign _GEN_37 = 7'h25 == WADDR ? 7'h25 : _GEN_36; // @[RAM_ST.scala 31:71]
  assign _GEN_38 = 7'h26 == WADDR ? 7'h26 : _GEN_37; // @[RAM_ST.scala 31:71]
  assign _GEN_39 = 7'h27 == WADDR ? 7'h27 : _GEN_38; // @[RAM_ST.scala 31:71]
  assign _GEN_40 = 7'h28 == WADDR ? 7'h28 : _GEN_39; // @[RAM_ST.scala 31:71]
  assign _GEN_41 = 7'h29 == WADDR ? 7'h29 : _GEN_40; // @[RAM_ST.scala 31:71]
  assign _GEN_42 = 7'h2a == WADDR ? 7'h2a : _GEN_41; // @[RAM_ST.scala 31:71]
  assign _GEN_43 = 7'h2b == WADDR ? 7'h2b : _GEN_42; // @[RAM_ST.scala 31:71]
  assign _GEN_44 = 7'h2c == WADDR ? 7'h2c : _GEN_43; // @[RAM_ST.scala 31:71]
  assign _GEN_45 = 7'h2d == WADDR ? 7'h2d : _GEN_44; // @[RAM_ST.scala 31:71]
  assign _GEN_46 = 7'h2e == WADDR ? 7'h2e : _GEN_45; // @[RAM_ST.scala 31:71]
  assign _GEN_47 = 7'h2f == WADDR ? 7'h2f : _GEN_46; // @[RAM_ST.scala 31:71]
  assign _GEN_48 = 7'h30 == WADDR ? 7'h30 : _GEN_47; // @[RAM_ST.scala 31:71]
  assign _GEN_49 = 7'h31 == WADDR ? 7'h31 : _GEN_48; // @[RAM_ST.scala 31:71]
  assign _GEN_50 = 7'h32 == WADDR ? 7'h32 : _GEN_49; // @[RAM_ST.scala 31:71]
  assign _GEN_51 = 7'h33 == WADDR ? 7'h33 : _GEN_50; // @[RAM_ST.scala 31:71]
  assign _GEN_52 = 7'h34 == WADDR ? 7'h34 : _GEN_51; // @[RAM_ST.scala 31:71]
  assign _GEN_53 = 7'h35 == WADDR ? 7'h35 : _GEN_52; // @[RAM_ST.scala 31:71]
  assign _GEN_54 = 7'h36 == WADDR ? 7'h36 : _GEN_53; // @[RAM_ST.scala 31:71]
  assign _GEN_55 = 7'h37 == WADDR ? 7'h37 : _GEN_54; // @[RAM_ST.scala 31:71]
  assign _GEN_56 = 7'h38 == WADDR ? 7'h38 : _GEN_55; // @[RAM_ST.scala 31:71]
  assign _GEN_57 = 7'h39 == WADDR ? 7'h39 : _GEN_56; // @[RAM_ST.scala 31:71]
  assign _GEN_58 = 7'h3a == WADDR ? 7'h3a : _GEN_57; // @[RAM_ST.scala 31:71]
  assign _GEN_59 = 7'h3b == WADDR ? 7'h3b : _GEN_58; // @[RAM_ST.scala 31:71]
  assign _GEN_60 = 7'h3c == WADDR ? 7'h3c : _GEN_59; // @[RAM_ST.scala 31:71]
  assign _GEN_61 = 7'h3d == WADDR ? 7'h3d : _GEN_60; // @[RAM_ST.scala 31:71]
  assign _GEN_62 = 7'h3e == WADDR ? 7'h3e : _GEN_61; // @[RAM_ST.scala 31:71]
  assign _GEN_63 = 7'h3f == WADDR ? 7'h3f : _GEN_62; // @[RAM_ST.scala 31:71]
  assign _GEN_64 = 7'h40 == WADDR ? 7'h40 : _GEN_63; // @[RAM_ST.scala 31:71]
  assign _GEN_65 = 7'h41 == WADDR ? 7'h41 : _GEN_64; // @[RAM_ST.scala 31:71]
  assign _GEN_66 = 7'h42 == WADDR ? 7'h42 : _GEN_65; // @[RAM_ST.scala 31:71]
  assign _GEN_67 = 7'h43 == WADDR ? 7'h43 : _GEN_66; // @[RAM_ST.scala 31:71]
  assign _GEN_68 = 7'h44 == WADDR ? 7'h44 : _GEN_67; // @[RAM_ST.scala 31:71]
  assign _GEN_69 = 7'h45 == WADDR ? 7'h45 : _GEN_68; // @[RAM_ST.scala 31:71]
  assign _GEN_70 = 7'h46 == WADDR ? 7'h46 : _GEN_69; // @[RAM_ST.scala 31:71]
  assign _GEN_71 = 7'h47 == WADDR ? 7'h47 : _GEN_70; // @[RAM_ST.scala 31:71]
  assign _GEN_72 = 7'h48 == WADDR ? 7'h48 : _GEN_71; // @[RAM_ST.scala 31:71]
  assign _GEN_73 = 7'h49 == WADDR ? 7'h49 : _GEN_72; // @[RAM_ST.scala 31:71]
  assign _GEN_74 = 7'h4a == WADDR ? 7'h4a : _GEN_73; // @[RAM_ST.scala 31:71]
  assign _GEN_75 = 7'h4b == WADDR ? 7'h4b : _GEN_74; // @[RAM_ST.scala 31:71]
  assign _GEN_76 = 7'h4c == WADDR ? 7'h4c : _GEN_75; // @[RAM_ST.scala 31:71]
  assign _GEN_77 = 7'h4d == WADDR ? 7'h4d : _GEN_76; // @[RAM_ST.scala 31:71]
  assign _GEN_78 = 7'h4e == WADDR ? 7'h4e : _GEN_77; // @[RAM_ST.scala 31:71]
  assign _GEN_79 = 7'h4f == WADDR ? 7'h4f : _GEN_78; // @[RAM_ST.scala 31:71]
  assign _GEN_80 = 7'h50 == WADDR ? 7'h50 : _GEN_79; // @[RAM_ST.scala 31:71]
  assign _GEN_81 = 7'h51 == WADDR ? 7'h51 : _GEN_80; // @[RAM_ST.scala 31:71]
  assign _GEN_82 = 7'h52 == WADDR ? 7'h52 : _GEN_81; // @[RAM_ST.scala 31:71]
  assign _GEN_83 = 7'h53 == WADDR ? 7'h53 : _GEN_82; // @[RAM_ST.scala 31:71]
  assign _GEN_84 = 7'h54 == WADDR ? 7'h54 : _GEN_83; // @[RAM_ST.scala 31:71]
  assign _GEN_85 = 7'h55 == WADDR ? 7'h55 : _GEN_84; // @[RAM_ST.scala 31:71]
  assign _GEN_86 = 7'h56 == WADDR ? 7'h56 : _GEN_85; // @[RAM_ST.scala 31:71]
  assign _GEN_87 = 7'h57 == WADDR ? 7'h57 : _GEN_86; // @[RAM_ST.scala 31:71]
  assign _GEN_88 = 7'h58 == WADDR ? 7'h58 : _GEN_87; // @[RAM_ST.scala 31:71]
  assign _GEN_89 = 7'h59 == WADDR ? 7'h59 : _GEN_88; // @[RAM_ST.scala 31:71]
  assign _GEN_90 = 7'h5a == WADDR ? 7'h5a : _GEN_89; // @[RAM_ST.scala 31:71]
  assign _GEN_91 = 7'h5b == WADDR ? 7'h5b : _GEN_90; // @[RAM_ST.scala 31:71]
  assign _GEN_92 = 7'h5c == WADDR ? 7'h5c : _GEN_91; // @[RAM_ST.scala 31:71]
  assign _GEN_93 = 7'h5d == WADDR ? 7'h5d : _GEN_92; // @[RAM_ST.scala 31:71]
  assign _GEN_94 = 7'h5e == WADDR ? 7'h5e : _GEN_93; // @[RAM_ST.scala 31:71]
  assign _GEN_95 = 7'h5f == WADDR ? 7'h5f : _GEN_94; // @[RAM_ST.scala 31:71]
  assign _GEN_96 = 7'h60 == WADDR ? 7'h60 : _GEN_95; // @[RAM_ST.scala 31:71]
  assign _GEN_97 = 7'h61 == WADDR ? 7'h61 : _GEN_96; // @[RAM_ST.scala 31:71]
  assign _GEN_98 = 7'h62 == WADDR ? 7'h62 : _GEN_97; // @[RAM_ST.scala 31:71]
  assign _GEN_99 = 7'h63 == WADDR ? 7'h63 : _GEN_98; // @[RAM_ST.scala 31:71]
  assign _GEN_100 = 7'h64 == WADDR ? 7'h64 : _GEN_99; // @[RAM_ST.scala 31:71]
  assign _GEN_101 = 7'h65 == WADDR ? 7'h65 : _GEN_100; // @[RAM_ST.scala 31:71]
  assign _GEN_102 = 7'h66 == WADDR ? 7'h66 : _GEN_101; // @[RAM_ST.scala 31:71]
  assign _GEN_103 = 7'h67 == WADDR ? 7'h67 : _GEN_102; // @[RAM_ST.scala 31:71]
  assign _GEN_104 = 7'h68 == WADDR ? 7'h68 : _GEN_103; // @[RAM_ST.scala 31:71]
  assign _GEN_105 = 7'h69 == WADDR ? 7'h69 : _GEN_104; // @[RAM_ST.scala 31:71]
  assign _GEN_106 = 7'h6a == WADDR ? 7'h6a : _GEN_105; // @[RAM_ST.scala 31:71]
  assign _GEN_107 = 7'h6b == WADDR ? 7'h6b : _GEN_106; // @[RAM_ST.scala 31:71]
  assign _GEN_108 = 7'h6c == WADDR ? 7'h6c : _GEN_107; // @[RAM_ST.scala 31:71]
  assign _GEN_109 = 7'h6d == WADDR ? 7'h6d : _GEN_108; // @[RAM_ST.scala 31:71]
  assign _GEN_110 = 7'h6e == WADDR ? 7'h6e : _GEN_109; // @[RAM_ST.scala 31:71]
  assign _GEN_111 = 7'h6f == WADDR ? 7'h6f : _GEN_110; // @[RAM_ST.scala 31:71]
  assign _GEN_112 = 7'h70 == WADDR ? 7'h70 : _GEN_111; // @[RAM_ST.scala 31:71]
  assign _GEN_113 = 7'h71 == WADDR ? 7'h71 : _GEN_112; // @[RAM_ST.scala 31:71]
  assign _GEN_114 = 7'h72 == WADDR ? 7'h72 : _GEN_113; // @[RAM_ST.scala 31:71]
  assign _GEN_115 = 7'h73 == WADDR ? 7'h73 : _GEN_114; // @[RAM_ST.scala 31:71]
  assign _GEN_116 = 7'h74 == WADDR ? 7'h74 : _GEN_115; // @[RAM_ST.scala 31:71]
  assign _GEN_117 = 7'h75 == WADDR ? 7'h75 : _GEN_116; // @[RAM_ST.scala 31:71]
  assign _GEN_118 = 7'h76 == WADDR ? 7'h76 : _GEN_117; // @[RAM_ST.scala 31:71]
  assign _GEN_119 = 7'h77 == WADDR ? 7'h77 : _GEN_118; // @[RAM_ST.scala 31:71]
  assign _T = {{1'd0}, _GEN_119}; // @[RAM_ST.scala 31:71]
  assign _GEN_126 = 7'h1 == RADDR ? 7'h1 : 7'h0; // @[RAM_ST.scala 32:46]
  assign _GEN_127 = 7'h2 == RADDR ? 7'h2 : _GEN_126; // @[RAM_ST.scala 32:46]
  assign _GEN_128 = 7'h3 == RADDR ? 7'h3 : _GEN_127; // @[RAM_ST.scala 32:46]
  assign _GEN_129 = 7'h4 == RADDR ? 7'h4 : _GEN_128; // @[RAM_ST.scala 32:46]
  assign _GEN_130 = 7'h5 == RADDR ? 7'h5 : _GEN_129; // @[RAM_ST.scala 32:46]
  assign _GEN_131 = 7'h6 == RADDR ? 7'h6 : _GEN_130; // @[RAM_ST.scala 32:46]
  assign _GEN_132 = 7'h7 == RADDR ? 7'h7 : _GEN_131; // @[RAM_ST.scala 32:46]
  assign _GEN_133 = 7'h8 == RADDR ? 7'h8 : _GEN_132; // @[RAM_ST.scala 32:46]
  assign _GEN_134 = 7'h9 == RADDR ? 7'h9 : _GEN_133; // @[RAM_ST.scala 32:46]
  assign _GEN_135 = 7'ha == RADDR ? 7'ha : _GEN_134; // @[RAM_ST.scala 32:46]
  assign _GEN_136 = 7'hb == RADDR ? 7'hb : _GEN_135; // @[RAM_ST.scala 32:46]
  assign _GEN_137 = 7'hc == RADDR ? 7'hc : _GEN_136; // @[RAM_ST.scala 32:46]
  assign _GEN_138 = 7'hd == RADDR ? 7'hd : _GEN_137; // @[RAM_ST.scala 32:46]
  assign _GEN_139 = 7'he == RADDR ? 7'he : _GEN_138; // @[RAM_ST.scala 32:46]
  assign _GEN_140 = 7'hf == RADDR ? 7'hf : _GEN_139; // @[RAM_ST.scala 32:46]
  assign _GEN_141 = 7'h10 == RADDR ? 7'h10 : _GEN_140; // @[RAM_ST.scala 32:46]
  assign _GEN_142 = 7'h11 == RADDR ? 7'h11 : _GEN_141; // @[RAM_ST.scala 32:46]
  assign _GEN_143 = 7'h12 == RADDR ? 7'h12 : _GEN_142; // @[RAM_ST.scala 32:46]
  assign _GEN_144 = 7'h13 == RADDR ? 7'h13 : _GEN_143; // @[RAM_ST.scala 32:46]
  assign _GEN_145 = 7'h14 == RADDR ? 7'h14 : _GEN_144; // @[RAM_ST.scala 32:46]
  assign _GEN_146 = 7'h15 == RADDR ? 7'h15 : _GEN_145; // @[RAM_ST.scala 32:46]
  assign _GEN_147 = 7'h16 == RADDR ? 7'h16 : _GEN_146; // @[RAM_ST.scala 32:46]
  assign _GEN_148 = 7'h17 == RADDR ? 7'h17 : _GEN_147; // @[RAM_ST.scala 32:46]
  assign _GEN_149 = 7'h18 == RADDR ? 7'h18 : _GEN_148; // @[RAM_ST.scala 32:46]
  assign _GEN_150 = 7'h19 == RADDR ? 7'h19 : _GEN_149; // @[RAM_ST.scala 32:46]
  assign _GEN_151 = 7'h1a == RADDR ? 7'h1a : _GEN_150; // @[RAM_ST.scala 32:46]
  assign _GEN_152 = 7'h1b == RADDR ? 7'h1b : _GEN_151; // @[RAM_ST.scala 32:46]
  assign _GEN_153 = 7'h1c == RADDR ? 7'h1c : _GEN_152; // @[RAM_ST.scala 32:46]
  assign _GEN_154 = 7'h1d == RADDR ? 7'h1d : _GEN_153; // @[RAM_ST.scala 32:46]
  assign _GEN_155 = 7'h1e == RADDR ? 7'h1e : _GEN_154; // @[RAM_ST.scala 32:46]
  assign _GEN_156 = 7'h1f == RADDR ? 7'h1f : _GEN_155; // @[RAM_ST.scala 32:46]
  assign _GEN_157 = 7'h20 == RADDR ? 7'h20 : _GEN_156; // @[RAM_ST.scala 32:46]
  assign _GEN_158 = 7'h21 == RADDR ? 7'h21 : _GEN_157; // @[RAM_ST.scala 32:46]
  assign _GEN_159 = 7'h22 == RADDR ? 7'h22 : _GEN_158; // @[RAM_ST.scala 32:46]
  assign _GEN_160 = 7'h23 == RADDR ? 7'h23 : _GEN_159; // @[RAM_ST.scala 32:46]
  assign _GEN_161 = 7'h24 == RADDR ? 7'h24 : _GEN_160; // @[RAM_ST.scala 32:46]
  assign _GEN_162 = 7'h25 == RADDR ? 7'h25 : _GEN_161; // @[RAM_ST.scala 32:46]
  assign _GEN_163 = 7'h26 == RADDR ? 7'h26 : _GEN_162; // @[RAM_ST.scala 32:46]
  assign _GEN_164 = 7'h27 == RADDR ? 7'h27 : _GEN_163; // @[RAM_ST.scala 32:46]
  assign _GEN_165 = 7'h28 == RADDR ? 7'h28 : _GEN_164; // @[RAM_ST.scala 32:46]
  assign _GEN_166 = 7'h29 == RADDR ? 7'h29 : _GEN_165; // @[RAM_ST.scala 32:46]
  assign _GEN_167 = 7'h2a == RADDR ? 7'h2a : _GEN_166; // @[RAM_ST.scala 32:46]
  assign _GEN_168 = 7'h2b == RADDR ? 7'h2b : _GEN_167; // @[RAM_ST.scala 32:46]
  assign _GEN_169 = 7'h2c == RADDR ? 7'h2c : _GEN_168; // @[RAM_ST.scala 32:46]
  assign _GEN_170 = 7'h2d == RADDR ? 7'h2d : _GEN_169; // @[RAM_ST.scala 32:46]
  assign _GEN_171 = 7'h2e == RADDR ? 7'h2e : _GEN_170; // @[RAM_ST.scala 32:46]
  assign _GEN_172 = 7'h2f == RADDR ? 7'h2f : _GEN_171; // @[RAM_ST.scala 32:46]
  assign _GEN_173 = 7'h30 == RADDR ? 7'h30 : _GEN_172; // @[RAM_ST.scala 32:46]
  assign _GEN_174 = 7'h31 == RADDR ? 7'h31 : _GEN_173; // @[RAM_ST.scala 32:46]
  assign _GEN_175 = 7'h32 == RADDR ? 7'h32 : _GEN_174; // @[RAM_ST.scala 32:46]
  assign _GEN_176 = 7'h33 == RADDR ? 7'h33 : _GEN_175; // @[RAM_ST.scala 32:46]
  assign _GEN_177 = 7'h34 == RADDR ? 7'h34 : _GEN_176; // @[RAM_ST.scala 32:46]
  assign _GEN_178 = 7'h35 == RADDR ? 7'h35 : _GEN_177; // @[RAM_ST.scala 32:46]
  assign _GEN_179 = 7'h36 == RADDR ? 7'h36 : _GEN_178; // @[RAM_ST.scala 32:46]
  assign _GEN_180 = 7'h37 == RADDR ? 7'h37 : _GEN_179; // @[RAM_ST.scala 32:46]
  assign _GEN_181 = 7'h38 == RADDR ? 7'h38 : _GEN_180; // @[RAM_ST.scala 32:46]
  assign _GEN_182 = 7'h39 == RADDR ? 7'h39 : _GEN_181; // @[RAM_ST.scala 32:46]
  assign _GEN_183 = 7'h3a == RADDR ? 7'h3a : _GEN_182; // @[RAM_ST.scala 32:46]
  assign _GEN_184 = 7'h3b == RADDR ? 7'h3b : _GEN_183; // @[RAM_ST.scala 32:46]
  assign _GEN_185 = 7'h3c == RADDR ? 7'h3c : _GEN_184; // @[RAM_ST.scala 32:46]
  assign _GEN_186 = 7'h3d == RADDR ? 7'h3d : _GEN_185; // @[RAM_ST.scala 32:46]
  assign _GEN_187 = 7'h3e == RADDR ? 7'h3e : _GEN_186; // @[RAM_ST.scala 32:46]
  assign _GEN_188 = 7'h3f == RADDR ? 7'h3f : _GEN_187; // @[RAM_ST.scala 32:46]
  assign _GEN_189 = 7'h40 == RADDR ? 7'h40 : _GEN_188; // @[RAM_ST.scala 32:46]
  assign _GEN_190 = 7'h41 == RADDR ? 7'h41 : _GEN_189; // @[RAM_ST.scala 32:46]
  assign _GEN_191 = 7'h42 == RADDR ? 7'h42 : _GEN_190; // @[RAM_ST.scala 32:46]
  assign _GEN_192 = 7'h43 == RADDR ? 7'h43 : _GEN_191; // @[RAM_ST.scala 32:46]
  assign _GEN_193 = 7'h44 == RADDR ? 7'h44 : _GEN_192; // @[RAM_ST.scala 32:46]
  assign _GEN_194 = 7'h45 == RADDR ? 7'h45 : _GEN_193; // @[RAM_ST.scala 32:46]
  assign _GEN_195 = 7'h46 == RADDR ? 7'h46 : _GEN_194; // @[RAM_ST.scala 32:46]
  assign _GEN_196 = 7'h47 == RADDR ? 7'h47 : _GEN_195; // @[RAM_ST.scala 32:46]
  assign _GEN_197 = 7'h48 == RADDR ? 7'h48 : _GEN_196; // @[RAM_ST.scala 32:46]
  assign _GEN_198 = 7'h49 == RADDR ? 7'h49 : _GEN_197; // @[RAM_ST.scala 32:46]
  assign _GEN_199 = 7'h4a == RADDR ? 7'h4a : _GEN_198; // @[RAM_ST.scala 32:46]
  assign _GEN_200 = 7'h4b == RADDR ? 7'h4b : _GEN_199; // @[RAM_ST.scala 32:46]
  assign _GEN_201 = 7'h4c == RADDR ? 7'h4c : _GEN_200; // @[RAM_ST.scala 32:46]
  assign _GEN_202 = 7'h4d == RADDR ? 7'h4d : _GEN_201; // @[RAM_ST.scala 32:46]
  assign _GEN_203 = 7'h4e == RADDR ? 7'h4e : _GEN_202; // @[RAM_ST.scala 32:46]
  assign _GEN_204 = 7'h4f == RADDR ? 7'h4f : _GEN_203; // @[RAM_ST.scala 32:46]
  assign _GEN_205 = 7'h50 == RADDR ? 7'h50 : _GEN_204; // @[RAM_ST.scala 32:46]
  assign _GEN_206 = 7'h51 == RADDR ? 7'h51 : _GEN_205; // @[RAM_ST.scala 32:46]
  assign _GEN_207 = 7'h52 == RADDR ? 7'h52 : _GEN_206; // @[RAM_ST.scala 32:46]
  assign _GEN_208 = 7'h53 == RADDR ? 7'h53 : _GEN_207; // @[RAM_ST.scala 32:46]
  assign _GEN_209 = 7'h54 == RADDR ? 7'h54 : _GEN_208; // @[RAM_ST.scala 32:46]
  assign _GEN_210 = 7'h55 == RADDR ? 7'h55 : _GEN_209; // @[RAM_ST.scala 32:46]
  assign _GEN_211 = 7'h56 == RADDR ? 7'h56 : _GEN_210; // @[RAM_ST.scala 32:46]
  assign _GEN_212 = 7'h57 == RADDR ? 7'h57 : _GEN_211; // @[RAM_ST.scala 32:46]
  assign _GEN_213 = 7'h58 == RADDR ? 7'h58 : _GEN_212; // @[RAM_ST.scala 32:46]
  assign _GEN_214 = 7'h59 == RADDR ? 7'h59 : _GEN_213; // @[RAM_ST.scala 32:46]
  assign _GEN_215 = 7'h5a == RADDR ? 7'h5a : _GEN_214; // @[RAM_ST.scala 32:46]
  assign _GEN_216 = 7'h5b == RADDR ? 7'h5b : _GEN_215; // @[RAM_ST.scala 32:46]
  assign _GEN_217 = 7'h5c == RADDR ? 7'h5c : _GEN_216; // @[RAM_ST.scala 32:46]
  assign _GEN_218 = 7'h5d == RADDR ? 7'h5d : _GEN_217; // @[RAM_ST.scala 32:46]
  assign _GEN_219 = 7'h5e == RADDR ? 7'h5e : _GEN_218; // @[RAM_ST.scala 32:46]
  assign _GEN_220 = 7'h5f == RADDR ? 7'h5f : _GEN_219; // @[RAM_ST.scala 32:46]
  assign _GEN_221 = 7'h60 == RADDR ? 7'h60 : _GEN_220; // @[RAM_ST.scala 32:46]
  assign _GEN_222 = 7'h61 == RADDR ? 7'h61 : _GEN_221; // @[RAM_ST.scala 32:46]
  assign _GEN_223 = 7'h62 == RADDR ? 7'h62 : _GEN_222; // @[RAM_ST.scala 32:46]
  assign _GEN_224 = 7'h63 == RADDR ? 7'h63 : _GEN_223; // @[RAM_ST.scala 32:46]
  assign _GEN_225 = 7'h64 == RADDR ? 7'h64 : _GEN_224; // @[RAM_ST.scala 32:46]
  assign _GEN_226 = 7'h65 == RADDR ? 7'h65 : _GEN_225; // @[RAM_ST.scala 32:46]
  assign _GEN_227 = 7'h66 == RADDR ? 7'h66 : _GEN_226; // @[RAM_ST.scala 32:46]
  assign _GEN_228 = 7'h67 == RADDR ? 7'h67 : _GEN_227; // @[RAM_ST.scala 32:46]
  assign _GEN_229 = 7'h68 == RADDR ? 7'h68 : _GEN_228; // @[RAM_ST.scala 32:46]
  assign _GEN_230 = 7'h69 == RADDR ? 7'h69 : _GEN_229; // @[RAM_ST.scala 32:46]
  assign _GEN_231 = 7'h6a == RADDR ? 7'h6a : _GEN_230; // @[RAM_ST.scala 32:46]
  assign _GEN_232 = 7'h6b == RADDR ? 7'h6b : _GEN_231; // @[RAM_ST.scala 32:46]
  assign _GEN_233 = 7'h6c == RADDR ? 7'h6c : _GEN_232; // @[RAM_ST.scala 32:46]
  assign _GEN_234 = 7'h6d == RADDR ? 7'h6d : _GEN_233; // @[RAM_ST.scala 32:46]
  assign _GEN_235 = 7'h6e == RADDR ? 7'h6e : _GEN_234; // @[RAM_ST.scala 32:46]
  assign _GEN_236 = 7'h6f == RADDR ? 7'h6f : _GEN_235; // @[RAM_ST.scala 32:46]
  assign _GEN_237 = 7'h70 == RADDR ? 7'h70 : _GEN_236; // @[RAM_ST.scala 32:46]
  assign _GEN_238 = 7'h71 == RADDR ? 7'h71 : _GEN_237; // @[RAM_ST.scala 32:46]
  assign _GEN_239 = 7'h72 == RADDR ? 7'h72 : _GEN_238; // @[RAM_ST.scala 32:46]
  assign _GEN_240 = 7'h73 == RADDR ? 7'h73 : _GEN_239; // @[RAM_ST.scala 32:46]
  assign _GEN_241 = 7'h74 == RADDR ? 7'h74 : _GEN_240; // @[RAM_ST.scala 32:46]
  assign _GEN_242 = 7'h75 == RADDR ? 7'h75 : _GEN_241; // @[RAM_ST.scala 32:46]
  assign _GEN_243 = 7'h76 == RADDR ? 7'h76 : _GEN_242; // @[RAM_ST.scala 32:46]
  assign _GEN_244 = 7'h77 == RADDR ? 7'h77 : _GEN_243; // @[RAM_ST.scala 32:46]
  assign _T_3 = {{1'd0}, _GEN_244}; // @[RAM_ST.scala 32:46]
  assign RDATA_0_0 = ram_0_0__T_8_data; // @[RAM_ST.scala 32:9]
  assign write_elem_counter_CE = WE; // @[RAM_ST.scala 23:25]
  assign read_elem_counter_CE = RE; // @[RAM_ST.scala 24:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 120; initvar = initvar+1)
    ram_0_0[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_0_0__T_8_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ram_0_0__T_8_addr_pipe_0 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_0_0__T_2_en & ram_0_0__T_2_mask) begin
      ram_0_0[ram_0_0__T_2_addr] <= ram_0_0__T_2_data; // @[RAM_ST.scala 29:24]
    end
    ram_0_0__T_8_en_pipe_0 <= read_elem_counter_valid;
    if (read_elem_counter_valid) begin
      ram_0_0__T_8_addr_pipe_0 <= _T_3[6:0];
    end
  end
endmodule
module ShiftT(
  input        clock,
  input        reset,
  input        valid_up,
  input  [7:0] I_0_0,
  output [7:0] O_0_0
);
  wire  RAM_ST_clock; // @[ShiftT.scala 39:29]
  wire  RAM_ST_RE; // @[ShiftT.scala 39:29]
  wire [6:0] RAM_ST_RADDR; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_RDATA_0_0; // @[ShiftT.scala 39:29]
  wire  RAM_ST_WE; // @[ShiftT.scala 39:29]
  wire [6:0] RAM_ST_WADDR; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_WDATA_0_0; // @[ShiftT.scala 39:29]
  wire  NestedCounters_CE; // @[ShiftT.scala 41:31]
  wire  NestedCounters_valid; // @[ShiftT.scala 41:31]
  reg [6:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[Counter.scala 37:24]
  wire [6:0] _T_3; // @[Counter.scala 38:22]
  RAM_ST RAM_ST ( // @[ShiftT.scala 39:29]
    .clock(RAM_ST_clock),
    .RE(RAM_ST_RE),
    .RADDR(RAM_ST_RADDR),
    .RDATA_0_0(RAM_ST_RDATA_0_0),
    .WE(RAM_ST_WE),
    .WADDR(RAM_ST_WADDR),
    .WDATA_0_0(RAM_ST_WDATA_0_0)
  );
  NestedCounters_2 NestedCounters ( // @[ShiftT.scala 41:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign _T_1 = value == 7'h77; // @[Counter.scala 37:24]
  assign _T_3 = value + 7'h1; // @[Counter.scala 38:22]
  assign O_0_0 = RAM_ST_RDATA_0_0; // @[ShiftT.scala 51:7]
  assign RAM_ST_clock = clock;
  assign RAM_ST_RE = valid_up; // @[ShiftT.scala 49:20]
  assign RAM_ST_RADDR = _T_1 ? 7'h0 : _T_3; // @[ShiftT.scala 46:76 ShiftT.scala 47:38]
  assign RAM_ST_WE = valid_up; // @[ShiftT.scala 48:20]
  assign RAM_ST_WADDR = value; // @[ShiftT.scala 45:23]
  assign RAM_ST_WDATA_0_0 = I_0_0; // @[ShiftT.scala 50:23]
  assign NestedCounters_CE = valid_up; // @[ShiftT.scala 42:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 7'h0;
    end else if (valid_up) begin
      if (_T_1) begin
        value <= 7'h0;
      end else begin
        value <= _T_3;
      end
    end
  end
endmodule
module ShiftTS(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_1_0_0,
  input  [7:0] I_2_0_0,
  input  [7:0] I_3_0_0,
  input  [7:0] I_4_0_0,
  input  [7:0] I_5_0_0,
  input  [7:0] I_6_0_0,
  input  [7:0] I_7_0_0,
  input  [7:0] I_8_0_0,
  input  [7:0] I_9_0_0,
  input  [7:0] I_10_0_0,
  input  [7:0] I_11_0_0,
  input  [7:0] I_12_0_0,
  input  [7:0] I_13_0_0,
  input  [7:0] I_14_0_0,
  input  [7:0] I_15_0_0,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0,
  output [7:0] O_8_0_0,
  output [7:0] O_9_0_0,
  output [7:0] O_10_0_0,
  output [7:0] O_11_0_0,
  output [7:0] O_12_0_0,
  output [7:0] O_13_0_0,
  output [7:0] O_14_0_0,
  output [7:0] O_15_0_0
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_1_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_1_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_1_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_1_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_1_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_2_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_2_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_2_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_2_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_2_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_3_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_3_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_3_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_3_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_3_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_4_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_4_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_4_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_4_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_4_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_5_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_5_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_5_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_5_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_5_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_6_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_6_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_6_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_6_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_6_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_7_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_7_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_7_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_7_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_7_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_8_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_8_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_8_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_8_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_8_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_9_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_9_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_9_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_9_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_9_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_10_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_10_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_10_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_10_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_10_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_11_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_11_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_11_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_11_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_11_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_12_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_12_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_12_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_12_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_12_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_13_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_13_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_13_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_13_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_13_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_14_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_14_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_14_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_14_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_14_O_0_0; // @[ShiftTS.scala 32:34]
  wire  ShiftT_15_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_15_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_15_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_15_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_15_O_0_0; // @[ShiftTS.scala 32:34]
  ShiftT ShiftT ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_clock),
    .reset(ShiftT_reset),
    .valid_up(ShiftT_valid_up),
    .I_0_0(ShiftT_I_0_0),
    .O_0_0(ShiftT_O_0_0)
  );
  ShiftT ShiftT_1 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_1_clock),
    .reset(ShiftT_1_reset),
    .valid_up(ShiftT_1_valid_up),
    .I_0_0(ShiftT_1_I_0_0),
    .O_0_0(ShiftT_1_O_0_0)
  );
  ShiftT ShiftT_2 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_2_clock),
    .reset(ShiftT_2_reset),
    .valid_up(ShiftT_2_valid_up),
    .I_0_0(ShiftT_2_I_0_0),
    .O_0_0(ShiftT_2_O_0_0)
  );
  ShiftT ShiftT_3 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_3_clock),
    .reset(ShiftT_3_reset),
    .valid_up(ShiftT_3_valid_up),
    .I_0_0(ShiftT_3_I_0_0),
    .O_0_0(ShiftT_3_O_0_0)
  );
  ShiftT ShiftT_4 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_4_clock),
    .reset(ShiftT_4_reset),
    .valid_up(ShiftT_4_valid_up),
    .I_0_0(ShiftT_4_I_0_0),
    .O_0_0(ShiftT_4_O_0_0)
  );
  ShiftT ShiftT_5 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_5_clock),
    .reset(ShiftT_5_reset),
    .valid_up(ShiftT_5_valid_up),
    .I_0_0(ShiftT_5_I_0_0),
    .O_0_0(ShiftT_5_O_0_0)
  );
  ShiftT ShiftT_6 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_6_clock),
    .reset(ShiftT_6_reset),
    .valid_up(ShiftT_6_valid_up),
    .I_0_0(ShiftT_6_I_0_0),
    .O_0_0(ShiftT_6_O_0_0)
  );
  ShiftT ShiftT_7 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_7_clock),
    .reset(ShiftT_7_reset),
    .valid_up(ShiftT_7_valid_up),
    .I_0_0(ShiftT_7_I_0_0),
    .O_0_0(ShiftT_7_O_0_0)
  );
  ShiftT ShiftT_8 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_8_clock),
    .reset(ShiftT_8_reset),
    .valid_up(ShiftT_8_valid_up),
    .I_0_0(ShiftT_8_I_0_0),
    .O_0_0(ShiftT_8_O_0_0)
  );
  ShiftT ShiftT_9 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_9_clock),
    .reset(ShiftT_9_reset),
    .valid_up(ShiftT_9_valid_up),
    .I_0_0(ShiftT_9_I_0_0),
    .O_0_0(ShiftT_9_O_0_0)
  );
  ShiftT ShiftT_10 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_10_clock),
    .reset(ShiftT_10_reset),
    .valid_up(ShiftT_10_valid_up),
    .I_0_0(ShiftT_10_I_0_0),
    .O_0_0(ShiftT_10_O_0_0)
  );
  ShiftT ShiftT_11 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_11_clock),
    .reset(ShiftT_11_reset),
    .valid_up(ShiftT_11_valid_up),
    .I_0_0(ShiftT_11_I_0_0),
    .O_0_0(ShiftT_11_O_0_0)
  );
  ShiftT ShiftT_12 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_12_clock),
    .reset(ShiftT_12_reset),
    .valid_up(ShiftT_12_valid_up),
    .I_0_0(ShiftT_12_I_0_0),
    .O_0_0(ShiftT_12_O_0_0)
  );
  ShiftT ShiftT_13 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_13_clock),
    .reset(ShiftT_13_reset),
    .valid_up(ShiftT_13_valid_up),
    .I_0_0(ShiftT_13_I_0_0),
    .O_0_0(ShiftT_13_O_0_0)
  );
  ShiftT ShiftT_14 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_14_clock),
    .reset(ShiftT_14_reset),
    .valid_up(ShiftT_14_valid_up),
    .I_0_0(ShiftT_14_I_0_0),
    .O_0_0(ShiftT_14_O_0_0)
  );
  ShiftT ShiftT_15 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_15_clock),
    .reset(ShiftT_15_reset),
    .valid_up(ShiftT_15_valid_up),
    .I_0_0(ShiftT_15_I_0_0),
    .O_0_0(ShiftT_15_O_0_0)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 39:14]
  assign O_0_0_0 = ShiftT_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_1_0_0 = ShiftT_1_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_2_0_0 = ShiftT_2_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_3_0_0 = ShiftT_3_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_4_0_0 = ShiftT_4_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_5_0_0 = ShiftT_5_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_6_0_0 = ShiftT_6_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_7_0_0 = ShiftT_7_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_8_0_0 = ShiftT_8_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_9_0_0 = ShiftT_9_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_10_0_0 = ShiftT_10_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_11_0_0 = ShiftT_11_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_12_0_0 = ShiftT_12_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_13_0_0 = ShiftT_13_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_14_0_0 = ShiftT_14_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_15_0_0 = ShiftT_15_O_0_0; // @[ShiftTS.scala 34:36]
  assign ShiftT_clock = clock;
  assign ShiftT_reset = reset;
  assign ShiftT_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_I_0_0 = I_0_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_1_clock = clock;
  assign ShiftT_1_reset = reset;
  assign ShiftT_1_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_1_I_0_0 = I_1_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_2_clock = clock;
  assign ShiftT_2_reset = reset;
  assign ShiftT_2_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_2_I_0_0 = I_2_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_3_clock = clock;
  assign ShiftT_3_reset = reset;
  assign ShiftT_3_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_3_I_0_0 = I_3_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_4_clock = clock;
  assign ShiftT_4_reset = reset;
  assign ShiftT_4_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_4_I_0_0 = I_4_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_5_clock = clock;
  assign ShiftT_5_reset = reset;
  assign ShiftT_5_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_5_I_0_0 = I_5_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_6_clock = clock;
  assign ShiftT_6_reset = reset;
  assign ShiftT_6_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_6_I_0_0 = I_6_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_7_clock = clock;
  assign ShiftT_7_reset = reset;
  assign ShiftT_7_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_7_I_0_0 = I_7_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_8_clock = clock;
  assign ShiftT_8_reset = reset;
  assign ShiftT_8_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_8_I_0_0 = I_8_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_9_clock = clock;
  assign ShiftT_9_reset = reset;
  assign ShiftT_9_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_9_I_0_0 = I_9_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_10_clock = clock;
  assign ShiftT_10_reset = reset;
  assign ShiftT_10_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_10_I_0_0 = I_10_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_11_clock = clock;
  assign ShiftT_11_reset = reset;
  assign ShiftT_11_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_11_I_0_0 = I_11_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_12_clock = clock;
  assign ShiftT_12_reset = reset;
  assign ShiftT_12_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_12_I_0_0 = I_12_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_13_clock = clock;
  assign ShiftT_13_reset = reset;
  assign ShiftT_13_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_13_I_0_0 = I_13_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_14_clock = clock;
  assign ShiftT_14_reset = reset;
  assign ShiftT_14_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_14_I_0_0 = I_14_0_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_15_clock = clock;
  assign ShiftT_15_reset = reset;
  assign ShiftT_15_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_15_I_0_0 = I_15_0_0; // @[ShiftTS.scala 33:24]
endmodule
module ShiftT_32(
  input        clock,
  input  [7:0] I_0_0,
  output [7:0] O_0_0
);
  reg [7:0] _T_0_0; // @[ShiftT.scala 24:82]
  reg [31:0] _RAND_0;
  assign O_0_0 = _T_0_0; // @[ShiftT.scala 24:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0_0 <= I_0_0;
  end
endmodule
module ShiftTS_2(
  input        clock,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_1_0_0,
  input  [7:0] I_2_0_0,
  input  [7:0] I_3_0_0,
  input  [7:0] I_4_0_0,
  input  [7:0] I_5_0_0,
  input  [7:0] I_6_0_0,
  input  [7:0] I_7_0_0,
  input  [7:0] I_8_0_0,
  input  [7:0] I_9_0_0,
  input  [7:0] I_10_0_0,
  input  [7:0] I_11_0_0,
  input  [7:0] I_12_0_0,
  input  [7:0] I_13_0_0,
  input  [7:0] I_14_0_0,
  input  [7:0] I_15_0_0,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0,
  output [7:0] O_8_0_0,
  output [7:0] O_9_0_0,
  output [7:0] O_10_0_0,
  output [7:0] O_11_0_0,
  output [7:0] O_12_0_0,
  output [7:0] O_13_0_0,
  output [7:0] O_14_0_0,
  output [7:0] O_15_0_0
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_I_0_0; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_O_0_0; // @[ShiftTS.scala 32:34]
  ShiftT_32 ShiftT ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_clock),
    .I_0_0(ShiftT_I_0_0),
    .O_0_0(ShiftT_O_0_0)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 39:14]
  assign O_0_0_0 = ShiftT_O_0_0; // @[ShiftTS.scala 34:36]
  assign O_1_0_0 = I_0_0_0; // @[ShiftTS.scala 29:36]
  assign O_2_0_0 = I_1_0_0; // @[ShiftTS.scala 29:36]
  assign O_3_0_0 = I_2_0_0; // @[ShiftTS.scala 29:36]
  assign O_4_0_0 = I_3_0_0; // @[ShiftTS.scala 29:36]
  assign O_5_0_0 = I_4_0_0; // @[ShiftTS.scala 29:36]
  assign O_6_0_0 = I_5_0_0; // @[ShiftTS.scala 29:36]
  assign O_7_0_0 = I_6_0_0; // @[ShiftTS.scala 29:36]
  assign O_8_0_0 = I_7_0_0; // @[ShiftTS.scala 29:36]
  assign O_9_0_0 = I_8_0_0; // @[ShiftTS.scala 29:36]
  assign O_10_0_0 = I_9_0_0; // @[ShiftTS.scala 29:36]
  assign O_11_0_0 = I_10_0_0; // @[ShiftTS.scala 29:36]
  assign O_12_0_0 = I_11_0_0; // @[ShiftTS.scala 29:36]
  assign O_13_0_0 = I_12_0_0; // @[ShiftTS.scala 29:36]
  assign O_14_0_0 = I_13_0_0; // @[ShiftTS.scala 29:36]
  assign O_15_0_0 = I_14_0_0; // @[ShiftTS.scala 29:36]
  assign ShiftT_clock = clock;
  assign ShiftT_I_0_0 = I_15_0_0; // @[ShiftTS.scala 33:24]
endmodule
module SSeqTupleCreator(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0 = I0; // @[Tuple.scala 12:32]
  assign O_1 = I1; // @[Tuple.scala 13:32]
endmodule
module Map2S(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I1_0,
  output [7:0] O_0_0,
  output [7:0] O_0_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1; // @[Map2S.scala 9:22]
  SSeqTupleCreator fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I1_0_0,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  Map2S fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I1_0(fst_op_I1_0),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_2(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_1_0_0,
  input  [7:0] I0_2_0_0,
  input  [7:0] I0_3_0_0,
  input  [7:0] I0_4_0_0,
  input  [7:0] I0_5_0_0,
  input  [7:0] I0_6_0_0,
  input  [7:0] I0_7_0_0,
  input  [7:0] I0_8_0_0,
  input  [7:0] I0_9_0_0,
  input  [7:0] I0_10_0_0,
  input  [7:0] I0_11_0_0,
  input  [7:0] I0_12_0_0,
  input  [7:0] I0_13_0_0,
  input  [7:0] I0_14_0_0,
  input  [7:0] I0_15_0_0,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_7_0_0,
  input  [7:0] I1_8_0_0,
  input  [7:0] I1_9_0_0,
  input  [7:0] I1_10_0_0,
  input  [7:0] I1_11_0_0,
  input  [7:0] I1_12_0_0,
  input  [7:0] I1_13_0_0,
  input  [7:0] I1_14_0_0,
  input  [7:0] I1_15_0_0,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_8_0_0_0,
  output [7:0] O_8_0_0_1,
  output [7:0] O_9_0_0_0,
  output [7:0] O_9_0_0_1,
  output [7:0] O_10_0_0_0,
  output [7:0] O_10_0_0_1,
  output [7:0] O_11_0_0_0,
  output [7:0] O_11_0_0_1,
  output [7:0] O_12_0_0_0,
  output [7:0] O_12_0_0_1,
  output [7:0] O_13_0_0_0,
  output [7:0] O_13_0_0_1,
  output [7:0] O_14_0_0_0,
  output [7:0] O_14_0_0_1,
  output [7:0] O_15_0_0_0,
  output [7:0] O_15_0_0_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_1; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0_1; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0_1; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  Map2S_1 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I1_0_0(fst_op_I1_0_0),
    .O_0_0_0(fst_op_O_0_0_0),
    .O_0_0_1(fst_op_O_0_0_1)
  );
  Map2S_1 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0(other_ops_0_I0_0_0),
    .I1_0_0(other_ops_0_I1_0_0),
    .O_0_0_0(other_ops_0_O_0_0_0),
    .O_0_0_1(other_ops_0_O_0_0_1)
  );
  Map2S_1 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0(other_ops_1_I0_0_0),
    .I1_0_0(other_ops_1_I1_0_0),
    .O_0_0_0(other_ops_1_O_0_0_0),
    .O_0_0_1(other_ops_1_O_0_0_1)
  );
  Map2S_1 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0(other_ops_2_I0_0_0),
    .I1_0_0(other_ops_2_I1_0_0),
    .O_0_0_0(other_ops_2_O_0_0_0),
    .O_0_0_1(other_ops_2_O_0_0_1)
  );
  Map2S_1 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0(other_ops_3_I0_0_0),
    .I1_0_0(other_ops_3_I1_0_0),
    .O_0_0_0(other_ops_3_O_0_0_0),
    .O_0_0_1(other_ops_3_O_0_0_1)
  );
  Map2S_1 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0(other_ops_4_I0_0_0),
    .I1_0_0(other_ops_4_I1_0_0),
    .O_0_0_0(other_ops_4_O_0_0_0),
    .O_0_0_1(other_ops_4_O_0_0_1)
  );
  Map2S_1 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0(other_ops_5_I0_0_0),
    .I1_0_0(other_ops_5_I1_0_0),
    .O_0_0_0(other_ops_5_O_0_0_0),
    .O_0_0_1(other_ops_5_O_0_0_1)
  );
  Map2S_1 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0(other_ops_6_I0_0_0),
    .I1_0_0(other_ops_6_I1_0_0),
    .O_0_0_0(other_ops_6_O_0_0_0),
    .O_0_0_1(other_ops_6_O_0_0_1)
  );
  Map2S_1 other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0_0(other_ops_7_I0_0_0),
    .I1_0_0(other_ops_7_I1_0_0),
    .O_0_0_0(other_ops_7_O_0_0_0),
    .O_0_0_1(other_ops_7_O_0_0_1)
  );
  Map2S_1 other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0_0(other_ops_8_I0_0_0),
    .I1_0_0(other_ops_8_I1_0_0),
    .O_0_0_0(other_ops_8_O_0_0_0),
    .O_0_0_1(other_ops_8_O_0_0_1)
  );
  Map2S_1 other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0_0(other_ops_9_I0_0_0),
    .I1_0_0(other_ops_9_I1_0_0),
    .O_0_0_0(other_ops_9_O_0_0_0),
    .O_0_0_1(other_ops_9_O_0_0_1)
  );
  Map2S_1 other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0_0(other_ops_10_I0_0_0),
    .I1_0_0(other_ops_10_I1_0_0),
    .O_0_0_0(other_ops_10_O_0_0_0),
    .O_0_0_1(other_ops_10_O_0_0_1)
  );
  Map2S_1 other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0_0(other_ops_11_I0_0_0),
    .I1_0_0(other_ops_11_I1_0_0),
    .O_0_0_0(other_ops_11_O_0_0_0),
    .O_0_0_1(other_ops_11_O_0_0_1)
  );
  Map2S_1 other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0_0(other_ops_12_I0_0_0),
    .I1_0_0(other_ops_12_I1_0_0),
    .O_0_0_0(other_ops_12_O_0_0_0),
    .O_0_0_1(other_ops_12_O_0_0_1)
  );
  Map2S_1 other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0_0(other_ops_13_I0_0_0),
    .I1_0_0(other_ops_13_I1_0_0),
    .O_0_0_0(other_ops_13_O_0_0_0),
    .O_0_0_1(other_ops_13_O_0_0_1)
  );
  Map2S_1 other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0_0(other_ops_14_I0_0_0),
    .I1_0_0(other_ops_14_I1_0_0),
    .O_0_0_0(other_ops_14_O_0_0_0),
    .O_0_0_1(other_ops_14_O_0_0_1)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0_0 = fst_op_O_0_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_0_1 = fst_op_O_0_0_1; // @[Map2S.scala 19:8]
  assign O_1_0_0_0 = other_ops_0_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_0_1 = other_ops_0_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_0_0 = other_ops_1_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_0_1 = other_ops_1_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_0_0 = other_ops_2_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_0_1 = other_ops_2_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_0_0 = other_ops_3_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_0_1 = other_ops_3_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_0_0 = other_ops_4_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_0_1 = other_ops_4_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_0_0 = other_ops_5_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_0_1 = other_ops_5_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_0_0 = other_ops_6_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_0_1 = other_ops_6_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_8_0_0_0 = other_ops_7_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_8_0_0_1 = other_ops_7_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_9_0_0_0 = other_ops_8_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_9_0_0_1 = other_ops_8_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_10_0_0_0 = other_ops_9_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_10_0_0_1 = other_ops_9_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_11_0_0_0 = other_ops_10_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_11_0_0_1 = other_ops_10_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_12_0_0_0 = other_ops_11_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_12_0_0_1 = other_ops_11_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_13_0_0_0 = other_ops_12_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_13_0_0_1 = other_ops_12_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_14_0_0_0 = other_ops_13_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_14_0_0_1 = other_ops_13_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_15_0_0_0 = other_ops_14_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_15_0_0_1 = other_ops_14_O_0_0_1; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_0 = I1_0_0_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0 = I0_1_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0_0 = I1_1_0_0; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0 = I0_2_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0_0 = I1_2_0_0; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0 = I0_3_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0_0 = I1_3_0_0; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0 = I0_4_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0_0 = I1_4_0_0; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0 = I0_5_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0_0 = I1_5_0_0; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0 = I0_6_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0_0 = I1_6_0_0; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0 = I0_7_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0_0 = I1_7_0_0; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0_0 = I0_8_0_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I1_0_0 = I1_8_0_0; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0_0 = I0_9_0_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I1_0_0 = I1_9_0_0; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0_0 = I0_10_0_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I1_0_0 = I1_10_0_0; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0_0 = I0_11_0_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I1_0_0 = I1_11_0_0; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0_0 = I0_12_0_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I1_0_0 = I1_12_0_0; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0_0 = I0_13_0_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I1_0_0 = I1_13_0_0; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0_0 = I0_14_0_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I1_0_0 = I1_14_0_0; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0_0 = I0_15_0_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I1_0_0 = I1_15_0_0; // @[Map2S.scala 23:43]
endmodule
module Map2T(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_1_0_0,
  input  [7:0] I0_2_0_0,
  input  [7:0] I0_3_0_0,
  input  [7:0] I0_4_0_0,
  input  [7:0] I0_5_0_0,
  input  [7:0] I0_6_0_0,
  input  [7:0] I0_7_0_0,
  input  [7:0] I0_8_0_0,
  input  [7:0] I0_9_0_0,
  input  [7:0] I0_10_0_0,
  input  [7:0] I0_11_0_0,
  input  [7:0] I0_12_0_0,
  input  [7:0] I0_13_0_0,
  input  [7:0] I0_14_0_0,
  input  [7:0] I0_15_0_0,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_7_0_0,
  input  [7:0] I1_8_0_0,
  input  [7:0] I1_9_0_0,
  input  [7:0] I1_10_0_0,
  input  [7:0] I1_11_0_0,
  input  [7:0] I1_12_0_0,
  input  [7:0] I1_13_0_0,
  input  [7:0] I1_14_0_0,
  input  [7:0] I1_15_0_0,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_8_0_0_0,
  output [7:0] O_8_0_0_1,
  output [7:0] O_9_0_0_0,
  output [7:0] O_9_0_0_1,
  output [7:0] O_10_0_0_0,
  output [7:0] O_10_0_0_1,
  output [7:0] O_11_0_0_0,
  output [7:0] O_11_0_0_1,
  output [7:0] O_12_0_0_0,
  output [7:0] O_12_0_0_1,
  output [7:0] O_13_0_0_0,
  output [7:0] O_13_0_0_1,
  output [7:0] O_14_0_0_0,
  output [7:0] O_14_0_0_1,
  output [7:0] O_15_0_0_0,
  output [7:0] O_15_0_0_1
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_0_1; // @[Map2T.scala 8:20]
  Map2S_2 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0(op_I0_0_0_0),
    .I0_1_0_0(op_I0_1_0_0),
    .I0_2_0_0(op_I0_2_0_0),
    .I0_3_0_0(op_I0_3_0_0),
    .I0_4_0_0(op_I0_4_0_0),
    .I0_5_0_0(op_I0_5_0_0),
    .I0_6_0_0(op_I0_6_0_0),
    .I0_7_0_0(op_I0_7_0_0),
    .I0_8_0_0(op_I0_8_0_0),
    .I0_9_0_0(op_I0_9_0_0),
    .I0_10_0_0(op_I0_10_0_0),
    .I0_11_0_0(op_I0_11_0_0),
    .I0_12_0_0(op_I0_12_0_0),
    .I0_13_0_0(op_I0_13_0_0),
    .I0_14_0_0(op_I0_14_0_0),
    .I0_15_0_0(op_I0_15_0_0),
    .I1_0_0_0(op_I1_0_0_0),
    .I1_1_0_0(op_I1_1_0_0),
    .I1_2_0_0(op_I1_2_0_0),
    .I1_3_0_0(op_I1_3_0_0),
    .I1_4_0_0(op_I1_4_0_0),
    .I1_5_0_0(op_I1_5_0_0),
    .I1_6_0_0(op_I1_6_0_0),
    .I1_7_0_0(op_I1_7_0_0),
    .I1_8_0_0(op_I1_8_0_0),
    .I1_9_0_0(op_I1_9_0_0),
    .I1_10_0_0(op_I1_10_0_0),
    .I1_11_0_0(op_I1_11_0_0),
    .I1_12_0_0(op_I1_12_0_0),
    .I1_13_0_0(op_I1_13_0_0),
    .I1_14_0_0(op_I1_14_0_0),
    .I1_15_0_0(op_I1_15_0_0),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_4_0_0_0(op_O_4_0_0_0),
    .O_4_0_0_1(op_O_4_0_0_1),
    .O_5_0_0_0(op_O_5_0_0_0),
    .O_5_0_0_1(op_O_5_0_0_1),
    .O_6_0_0_0(op_O_6_0_0_0),
    .O_6_0_0_1(op_O_6_0_0_1),
    .O_7_0_0_0(op_O_7_0_0_0),
    .O_7_0_0_1(op_O_7_0_0_1),
    .O_8_0_0_0(op_O_8_0_0_0),
    .O_8_0_0_1(op_O_8_0_0_1),
    .O_9_0_0_0(op_O_9_0_0_0),
    .O_9_0_0_1(op_O_9_0_0_1),
    .O_10_0_0_0(op_O_10_0_0_0),
    .O_10_0_0_1(op_O_10_0_0_1),
    .O_11_0_0_0(op_O_11_0_0_0),
    .O_11_0_0_1(op_O_11_0_0_1),
    .O_12_0_0_0(op_O_12_0_0_0),
    .O_12_0_0_1(op_O_12_0_0_1),
    .O_13_0_0_0(op_O_13_0_0_0),
    .O_13_0_0_1(op_O_13_0_0_1),
    .O_14_0_0_0(op_O_14_0_0_0),
    .O_14_0_0_1(op_O_14_0_0_1),
    .O_15_0_0_0(op_O_15_0_0_0),
    .O_15_0_0_1(op_O_15_0_0_1)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_0_0 = op_O_4_0_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_0_1 = op_O_4_0_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_0_0 = op_O_5_0_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_0_1 = op_O_5_0_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_0_0 = op_O_6_0_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_0_1 = op_O_6_0_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_0_0 = op_O_7_0_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_0_1 = op_O_7_0_0_1; // @[Map2T.scala 17:7]
  assign O_8_0_0_0 = op_O_8_0_0_0; // @[Map2T.scala 17:7]
  assign O_8_0_0_1 = op_O_8_0_0_1; // @[Map2T.scala 17:7]
  assign O_9_0_0_0 = op_O_9_0_0_0; // @[Map2T.scala 17:7]
  assign O_9_0_0_1 = op_O_9_0_0_1; // @[Map2T.scala 17:7]
  assign O_10_0_0_0 = op_O_10_0_0_0; // @[Map2T.scala 17:7]
  assign O_10_0_0_1 = op_O_10_0_0_1; // @[Map2T.scala 17:7]
  assign O_11_0_0_0 = op_O_11_0_0_0; // @[Map2T.scala 17:7]
  assign O_11_0_0_1 = op_O_11_0_0_1; // @[Map2T.scala 17:7]
  assign O_12_0_0_0 = op_O_12_0_0_0; // @[Map2T.scala 17:7]
  assign O_12_0_0_1 = op_O_12_0_0_1; // @[Map2T.scala 17:7]
  assign O_13_0_0_0 = op_O_13_0_0_0; // @[Map2T.scala 17:7]
  assign O_13_0_0_1 = op_O_13_0_0_1; // @[Map2T.scala 17:7]
  assign O_14_0_0_0 = op_O_14_0_0_0; // @[Map2T.scala 17:7]
  assign O_14_0_0_1 = op_O_14_0_0_1; // @[Map2T.scala 17:7]
  assign O_15_0_0_0 = op_O_15_0_0_0; // @[Map2T.scala 17:7]
  assign O_15_0_0_1 = op_O_15_0_0_1; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0 = I0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0 = I0_1_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0 = I0_2_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0 = I0_3_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0 = I0_4_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0 = I0_5_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0 = I0_6_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0 = I0_7_0_0; // @[Map2T.scala 15:11]
  assign op_I0_8_0_0 = I0_8_0_0; // @[Map2T.scala 15:11]
  assign op_I0_9_0_0 = I0_9_0_0; // @[Map2T.scala 15:11]
  assign op_I0_10_0_0 = I0_10_0_0; // @[Map2T.scala 15:11]
  assign op_I0_11_0_0 = I0_11_0_0; // @[Map2T.scala 15:11]
  assign op_I0_12_0_0 = I0_12_0_0; // @[Map2T.scala 15:11]
  assign op_I0_13_0_0 = I0_13_0_0; // @[Map2T.scala 15:11]
  assign op_I0_14_0_0 = I0_14_0_0; // @[Map2T.scala 15:11]
  assign op_I0_15_0_0 = I0_15_0_0; // @[Map2T.scala 15:11]
  assign op_I1_0_0_0 = I1_0_0_0; // @[Map2T.scala 16:11]
  assign op_I1_1_0_0 = I1_1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_2_0_0 = I1_2_0_0; // @[Map2T.scala 16:11]
  assign op_I1_3_0_0 = I1_3_0_0; // @[Map2T.scala 16:11]
  assign op_I1_4_0_0 = I1_4_0_0; // @[Map2T.scala 16:11]
  assign op_I1_5_0_0 = I1_5_0_0; // @[Map2T.scala 16:11]
  assign op_I1_6_0_0 = I1_6_0_0; // @[Map2T.scala 16:11]
  assign op_I1_7_0_0 = I1_7_0_0; // @[Map2T.scala 16:11]
  assign op_I1_8_0_0 = I1_8_0_0; // @[Map2T.scala 16:11]
  assign op_I1_9_0_0 = I1_9_0_0; // @[Map2T.scala 16:11]
  assign op_I1_10_0_0 = I1_10_0_0; // @[Map2T.scala 16:11]
  assign op_I1_11_0_0 = I1_11_0_0; // @[Map2T.scala 16:11]
  assign op_I1_12_0_0 = I1_12_0_0; // @[Map2T.scala 16:11]
  assign op_I1_13_0_0 = I1_13_0_0; // @[Map2T.scala 16:11]
  assign op_I1_14_0_0 = I1_14_0_0; // @[Map2T.scala 16:11]
  assign op_I1_15_0_0 = I1_15_0_0; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0 = I0_0; // @[Tuple.scala 24:34]
  assign O_1 = I0_1; // @[Tuple.scala 24:34]
  assign O_2 = I1; // @[Tuple.scala 26:32]
endmodule
module Map2S_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I1_0,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2; // @[Map2S.scala 9:22]
  SSeqTupleAppender fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_0_2 = fst_op_O_2; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_0_0_1,
  input  [7:0] I1_0_0,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  Map2S_3 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I1_0(fst_op_I1_0),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_5(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0_0,
  input  [7:0] I0_0_0_0_1,
  input  [7:0] I0_1_0_0_0,
  input  [7:0] I0_1_0_0_1,
  input  [7:0] I0_2_0_0_0,
  input  [7:0] I0_2_0_0_1,
  input  [7:0] I0_3_0_0_0,
  input  [7:0] I0_3_0_0_1,
  input  [7:0] I0_4_0_0_0,
  input  [7:0] I0_4_0_0_1,
  input  [7:0] I0_5_0_0_0,
  input  [7:0] I0_5_0_0_1,
  input  [7:0] I0_6_0_0_0,
  input  [7:0] I0_6_0_0_1,
  input  [7:0] I0_7_0_0_0,
  input  [7:0] I0_7_0_0_1,
  input  [7:0] I0_8_0_0_0,
  input  [7:0] I0_8_0_0_1,
  input  [7:0] I0_9_0_0_0,
  input  [7:0] I0_9_0_0_1,
  input  [7:0] I0_10_0_0_0,
  input  [7:0] I0_10_0_0_1,
  input  [7:0] I0_11_0_0_0,
  input  [7:0] I0_11_0_0_1,
  input  [7:0] I0_12_0_0_0,
  input  [7:0] I0_12_0_0_1,
  input  [7:0] I0_13_0_0_0,
  input  [7:0] I0_13_0_0_1,
  input  [7:0] I0_14_0_0_0,
  input  [7:0] I0_14_0_0_1,
  input  [7:0] I0_15_0_0_0,
  input  [7:0] I0_15_0_0_1,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_7_0_0,
  input  [7:0] I1_8_0_0,
  input  [7:0] I1_9_0_0,
  input  [7:0] I1_10_0_0,
  input  [7:0] I1_11_0_0,
  input  [7:0] I1_12_0_0,
  input  [7:0] I1_13_0_0,
  input  [7:0] I1_14_0_0,
  input  [7:0] I1_15_0_0,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_0_2,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_0_2,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_0_2,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_0_2,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_0_2,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_0_2,
  output [7:0] O_8_0_0_0,
  output [7:0] O_8_0_0_1,
  output [7:0] O_8_0_0_2,
  output [7:0] O_9_0_0_0,
  output [7:0] O_9_0_0_1,
  output [7:0] O_9_0_0_2,
  output [7:0] O_10_0_0_0,
  output [7:0] O_10_0_0_1,
  output [7:0] O_10_0_0_2,
  output [7:0] O_11_0_0_0,
  output [7:0] O_11_0_0_1,
  output [7:0] O_11_0_0_2,
  output [7:0] O_12_0_0_0,
  output [7:0] O_12_0_0_1,
  output [7:0] O_12_0_0_2,
  output [7:0] O_13_0_0_0,
  output [7:0] O_13_0_0_1,
  output [7:0] O_13_0_0_2,
  output [7:0] O_14_0_0_0,
  output [7:0] O_14_0_0_1,
  output [7:0] O_14_0_0_2,
  output [7:0] O_15_0_0_0,
  output [7:0] O_15_0_0_1,
  output [7:0] O_15_0_0_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  Map2S_4 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0_0(fst_op_I0_0_0_0),
    .I0_0_0_1(fst_op_I0_0_0_1),
    .I1_0_0(fst_op_I1_0_0),
    .O_0_0_0(fst_op_O_0_0_0),
    .O_0_0_1(fst_op_O_0_0_1),
    .O_0_0_2(fst_op_O_0_0_2)
  );
  Map2S_4 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0_0(other_ops_0_I0_0_0_0),
    .I0_0_0_1(other_ops_0_I0_0_0_1),
    .I1_0_0(other_ops_0_I1_0_0),
    .O_0_0_0(other_ops_0_O_0_0_0),
    .O_0_0_1(other_ops_0_O_0_0_1),
    .O_0_0_2(other_ops_0_O_0_0_2)
  );
  Map2S_4 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0_0(other_ops_1_I0_0_0_0),
    .I0_0_0_1(other_ops_1_I0_0_0_1),
    .I1_0_0(other_ops_1_I1_0_0),
    .O_0_0_0(other_ops_1_O_0_0_0),
    .O_0_0_1(other_ops_1_O_0_0_1),
    .O_0_0_2(other_ops_1_O_0_0_2)
  );
  Map2S_4 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0_0(other_ops_2_I0_0_0_0),
    .I0_0_0_1(other_ops_2_I0_0_0_1),
    .I1_0_0(other_ops_2_I1_0_0),
    .O_0_0_0(other_ops_2_O_0_0_0),
    .O_0_0_1(other_ops_2_O_0_0_1),
    .O_0_0_2(other_ops_2_O_0_0_2)
  );
  Map2S_4 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0_0(other_ops_3_I0_0_0_0),
    .I0_0_0_1(other_ops_3_I0_0_0_1),
    .I1_0_0(other_ops_3_I1_0_0),
    .O_0_0_0(other_ops_3_O_0_0_0),
    .O_0_0_1(other_ops_3_O_0_0_1),
    .O_0_0_2(other_ops_3_O_0_0_2)
  );
  Map2S_4 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0_0(other_ops_4_I0_0_0_0),
    .I0_0_0_1(other_ops_4_I0_0_0_1),
    .I1_0_0(other_ops_4_I1_0_0),
    .O_0_0_0(other_ops_4_O_0_0_0),
    .O_0_0_1(other_ops_4_O_0_0_1),
    .O_0_0_2(other_ops_4_O_0_0_2)
  );
  Map2S_4 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0_0(other_ops_5_I0_0_0_0),
    .I0_0_0_1(other_ops_5_I0_0_0_1),
    .I1_0_0(other_ops_5_I1_0_0),
    .O_0_0_0(other_ops_5_O_0_0_0),
    .O_0_0_1(other_ops_5_O_0_0_1),
    .O_0_0_2(other_ops_5_O_0_0_2)
  );
  Map2S_4 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0_0(other_ops_6_I0_0_0_0),
    .I0_0_0_1(other_ops_6_I0_0_0_1),
    .I1_0_0(other_ops_6_I1_0_0),
    .O_0_0_0(other_ops_6_O_0_0_0),
    .O_0_0_1(other_ops_6_O_0_0_1),
    .O_0_0_2(other_ops_6_O_0_0_2)
  );
  Map2S_4 other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0_0_0(other_ops_7_I0_0_0_0),
    .I0_0_0_1(other_ops_7_I0_0_0_1),
    .I1_0_0(other_ops_7_I1_0_0),
    .O_0_0_0(other_ops_7_O_0_0_0),
    .O_0_0_1(other_ops_7_O_0_0_1),
    .O_0_0_2(other_ops_7_O_0_0_2)
  );
  Map2S_4 other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0_0_0(other_ops_8_I0_0_0_0),
    .I0_0_0_1(other_ops_8_I0_0_0_1),
    .I1_0_0(other_ops_8_I1_0_0),
    .O_0_0_0(other_ops_8_O_0_0_0),
    .O_0_0_1(other_ops_8_O_0_0_1),
    .O_0_0_2(other_ops_8_O_0_0_2)
  );
  Map2S_4 other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0_0_0(other_ops_9_I0_0_0_0),
    .I0_0_0_1(other_ops_9_I0_0_0_1),
    .I1_0_0(other_ops_9_I1_0_0),
    .O_0_0_0(other_ops_9_O_0_0_0),
    .O_0_0_1(other_ops_9_O_0_0_1),
    .O_0_0_2(other_ops_9_O_0_0_2)
  );
  Map2S_4 other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0_0_0(other_ops_10_I0_0_0_0),
    .I0_0_0_1(other_ops_10_I0_0_0_1),
    .I1_0_0(other_ops_10_I1_0_0),
    .O_0_0_0(other_ops_10_O_0_0_0),
    .O_0_0_1(other_ops_10_O_0_0_1),
    .O_0_0_2(other_ops_10_O_0_0_2)
  );
  Map2S_4 other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0_0_0(other_ops_11_I0_0_0_0),
    .I0_0_0_1(other_ops_11_I0_0_0_1),
    .I1_0_0(other_ops_11_I1_0_0),
    .O_0_0_0(other_ops_11_O_0_0_0),
    .O_0_0_1(other_ops_11_O_0_0_1),
    .O_0_0_2(other_ops_11_O_0_0_2)
  );
  Map2S_4 other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0_0_0(other_ops_12_I0_0_0_0),
    .I0_0_0_1(other_ops_12_I0_0_0_1),
    .I1_0_0(other_ops_12_I1_0_0),
    .O_0_0_0(other_ops_12_O_0_0_0),
    .O_0_0_1(other_ops_12_O_0_0_1),
    .O_0_0_2(other_ops_12_O_0_0_2)
  );
  Map2S_4 other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0_0_0(other_ops_13_I0_0_0_0),
    .I0_0_0_1(other_ops_13_I0_0_0_1),
    .I1_0_0(other_ops_13_I1_0_0),
    .O_0_0_0(other_ops_13_O_0_0_0),
    .O_0_0_1(other_ops_13_O_0_0_1),
    .O_0_0_2(other_ops_13_O_0_0_2)
  );
  Map2S_4 other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0_0_0(other_ops_14_I0_0_0_0),
    .I0_0_0_1(other_ops_14_I0_0_0_1),
    .I1_0_0(other_ops_14_I1_0_0),
    .O_0_0_0(other_ops_14_O_0_0_0),
    .O_0_0_1(other_ops_14_O_0_0_1),
    .O_0_0_2(other_ops_14_O_0_0_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0_0 = fst_op_O_0_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_0_1 = fst_op_O_0_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_0_2 = fst_op_O_0_0_2; // @[Map2S.scala 19:8]
  assign O_1_0_0_0 = other_ops_0_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_0_1 = other_ops_0_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_0_2 = other_ops_0_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_2_0_0_0 = other_ops_1_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_0_1 = other_ops_1_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_0_2 = other_ops_1_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_3_0_0_0 = other_ops_2_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_0_1 = other_ops_2_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_0_2 = other_ops_2_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_4_0_0_0 = other_ops_3_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_0_1 = other_ops_3_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_0_2 = other_ops_3_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_5_0_0_0 = other_ops_4_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_0_1 = other_ops_4_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_0_2 = other_ops_4_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_6_0_0_0 = other_ops_5_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_0_1 = other_ops_5_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_0_2 = other_ops_5_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_7_0_0_0 = other_ops_6_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_0_1 = other_ops_6_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_0_2 = other_ops_6_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_8_0_0_0 = other_ops_7_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_8_0_0_1 = other_ops_7_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_8_0_0_2 = other_ops_7_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_9_0_0_0 = other_ops_8_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_9_0_0_1 = other_ops_8_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_9_0_0_2 = other_ops_8_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_10_0_0_0 = other_ops_9_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_10_0_0_1 = other_ops_9_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_10_0_0_2 = other_ops_9_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_11_0_0_0 = other_ops_10_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_11_0_0_1 = other_ops_10_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_11_0_0_2 = other_ops_10_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_12_0_0_0 = other_ops_11_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_12_0_0_1 = other_ops_11_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_12_0_0_2 = other_ops_11_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_13_0_0_0 = other_ops_12_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_13_0_0_1 = other_ops_12_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_13_0_0_2 = other_ops_12_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_14_0_0_0 = other_ops_13_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_14_0_0_1 = other_ops_13_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_14_0_0_2 = other_ops_13_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_15_0_0_0 = other_ops_14_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_15_0_0_1 = other_ops_14_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_15_0_0_2 = other_ops_14_O_0_0_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0_0 = I0_0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_0_1 = I0_0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_0 = I1_0_0_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0_0 = I0_1_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_0_1 = I0_1_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0_0 = I1_1_0_0; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0_0 = I0_2_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_0_1 = I0_2_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0_0 = I1_2_0_0; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0_0 = I0_3_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_0_1 = I0_3_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0_0 = I1_3_0_0; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0_0 = I0_4_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_0_1 = I0_4_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0_0 = I1_4_0_0; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0_0 = I0_5_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_0_1 = I0_5_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0_0 = I1_5_0_0; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0_0 = I0_6_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_0_1 = I0_6_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0_0 = I1_6_0_0; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0_0 = I0_7_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_0_1 = I0_7_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0_0 = I1_7_0_0; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0_0_0 = I0_8_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_0_1 = I0_8_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I1_0_0 = I1_8_0_0; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0_0_0 = I0_9_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_0_1 = I0_9_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I1_0_0 = I1_9_0_0; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0_0_0 = I0_10_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_0_1 = I0_10_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I1_0_0 = I1_10_0_0; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0_0_0 = I0_11_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_0_1 = I0_11_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I1_0_0 = I1_11_0_0; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0_0_0 = I0_12_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_0_1 = I0_12_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I1_0_0 = I1_12_0_0; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0_0_0 = I0_13_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_0_1 = I0_13_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I1_0_0 = I1_13_0_0; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0_0_0 = I0_14_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_0_1 = I0_14_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I1_0_0 = I1_14_0_0; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0_0_0 = I0_15_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_0_1 = I0_15_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I1_0_0 = I1_15_0_0; // @[Map2S.scala 23:43]
endmodule
module Map2T_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0_0,
  input  [7:0] I0_0_0_0_1,
  input  [7:0] I0_1_0_0_0,
  input  [7:0] I0_1_0_0_1,
  input  [7:0] I0_2_0_0_0,
  input  [7:0] I0_2_0_0_1,
  input  [7:0] I0_3_0_0_0,
  input  [7:0] I0_3_0_0_1,
  input  [7:0] I0_4_0_0_0,
  input  [7:0] I0_4_0_0_1,
  input  [7:0] I0_5_0_0_0,
  input  [7:0] I0_5_0_0_1,
  input  [7:0] I0_6_0_0_0,
  input  [7:0] I0_6_0_0_1,
  input  [7:0] I0_7_0_0_0,
  input  [7:0] I0_7_0_0_1,
  input  [7:0] I0_8_0_0_0,
  input  [7:0] I0_8_0_0_1,
  input  [7:0] I0_9_0_0_0,
  input  [7:0] I0_9_0_0_1,
  input  [7:0] I0_10_0_0_0,
  input  [7:0] I0_10_0_0_1,
  input  [7:0] I0_11_0_0_0,
  input  [7:0] I0_11_0_0_1,
  input  [7:0] I0_12_0_0_0,
  input  [7:0] I0_12_0_0_1,
  input  [7:0] I0_13_0_0_0,
  input  [7:0] I0_13_0_0_1,
  input  [7:0] I0_14_0_0_0,
  input  [7:0] I0_14_0_0_1,
  input  [7:0] I0_15_0_0_0,
  input  [7:0] I0_15_0_0_1,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_7_0_0,
  input  [7:0] I1_8_0_0,
  input  [7:0] I1_9_0_0,
  input  [7:0] I1_10_0_0,
  input  [7:0] I1_11_0_0,
  input  [7:0] I1_12_0_0,
  input  [7:0] I1_13_0_0,
  input  [7:0] I1_14_0_0,
  input  [7:0] I1_15_0_0,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_0_2,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_0_2,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_0_2,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_0_2,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_0_2,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_0_2,
  output [7:0] O_8_0_0_0,
  output [7:0] O_8_0_0_1,
  output [7:0] O_8_0_0_2,
  output [7:0] O_9_0_0_0,
  output [7:0] O_9_0_0_1,
  output [7:0] O_9_0_0_2,
  output [7:0] O_10_0_0_0,
  output [7:0] O_10_0_0_1,
  output [7:0] O_10_0_0_2,
  output [7:0] O_11_0_0_0,
  output [7:0] O_11_0_0_1,
  output [7:0] O_11_0_0_2,
  output [7:0] O_12_0_0_0,
  output [7:0] O_12_0_0_1,
  output [7:0] O_12_0_0_2,
  output [7:0] O_13_0_0_0,
  output [7:0] O_13_0_0_1,
  output [7:0] O_13_0_0_2,
  output [7:0] O_14_0_0_0,
  output [7:0] O_14_0_0_1,
  output [7:0] O_14_0_0_2,
  output [7:0] O_15_0_0_0,
  output [7:0] O_15_0_0_1,
  output [7:0] O_15_0_0_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_0_2; // @[Map2T.scala 8:20]
  Map2S_5 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0_0(op_I0_0_0_0_0),
    .I0_0_0_0_1(op_I0_0_0_0_1),
    .I0_1_0_0_0(op_I0_1_0_0_0),
    .I0_1_0_0_1(op_I0_1_0_0_1),
    .I0_2_0_0_0(op_I0_2_0_0_0),
    .I0_2_0_0_1(op_I0_2_0_0_1),
    .I0_3_0_0_0(op_I0_3_0_0_0),
    .I0_3_0_0_1(op_I0_3_0_0_1),
    .I0_4_0_0_0(op_I0_4_0_0_0),
    .I0_4_0_0_1(op_I0_4_0_0_1),
    .I0_5_0_0_0(op_I0_5_0_0_0),
    .I0_5_0_0_1(op_I0_5_0_0_1),
    .I0_6_0_0_0(op_I0_6_0_0_0),
    .I0_6_0_0_1(op_I0_6_0_0_1),
    .I0_7_0_0_0(op_I0_7_0_0_0),
    .I0_7_0_0_1(op_I0_7_0_0_1),
    .I0_8_0_0_0(op_I0_8_0_0_0),
    .I0_8_0_0_1(op_I0_8_0_0_1),
    .I0_9_0_0_0(op_I0_9_0_0_0),
    .I0_9_0_0_1(op_I0_9_0_0_1),
    .I0_10_0_0_0(op_I0_10_0_0_0),
    .I0_10_0_0_1(op_I0_10_0_0_1),
    .I0_11_0_0_0(op_I0_11_0_0_0),
    .I0_11_0_0_1(op_I0_11_0_0_1),
    .I0_12_0_0_0(op_I0_12_0_0_0),
    .I0_12_0_0_1(op_I0_12_0_0_1),
    .I0_13_0_0_0(op_I0_13_0_0_0),
    .I0_13_0_0_1(op_I0_13_0_0_1),
    .I0_14_0_0_0(op_I0_14_0_0_0),
    .I0_14_0_0_1(op_I0_14_0_0_1),
    .I0_15_0_0_0(op_I0_15_0_0_0),
    .I0_15_0_0_1(op_I0_15_0_0_1),
    .I1_0_0_0(op_I1_0_0_0),
    .I1_1_0_0(op_I1_1_0_0),
    .I1_2_0_0(op_I1_2_0_0),
    .I1_3_0_0(op_I1_3_0_0),
    .I1_4_0_0(op_I1_4_0_0),
    .I1_5_0_0(op_I1_5_0_0),
    .I1_6_0_0(op_I1_6_0_0),
    .I1_7_0_0(op_I1_7_0_0),
    .I1_8_0_0(op_I1_8_0_0),
    .I1_9_0_0(op_I1_9_0_0),
    .I1_10_0_0(op_I1_10_0_0),
    .I1_11_0_0(op_I1_11_0_0),
    .I1_12_0_0(op_I1_12_0_0),
    .I1_13_0_0(op_I1_13_0_0),
    .I1_14_0_0(op_I1_14_0_0),
    .I1_15_0_0(op_I1_15_0_0),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_0_0_0_2(op_O_0_0_0_2),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_1_0_0_2(op_O_1_0_0_2),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_2_0_0_2(op_O_2_0_0_2),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_3_0_0_2(op_O_3_0_0_2),
    .O_4_0_0_0(op_O_4_0_0_0),
    .O_4_0_0_1(op_O_4_0_0_1),
    .O_4_0_0_2(op_O_4_0_0_2),
    .O_5_0_0_0(op_O_5_0_0_0),
    .O_5_0_0_1(op_O_5_0_0_1),
    .O_5_0_0_2(op_O_5_0_0_2),
    .O_6_0_0_0(op_O_6_0_0_0),
    .O_6_0_0_1(op_O_6_0_0_1),
    .O_6_0_0_2(op_O_6_0_0_2),
    .O_7_0_0_0(op_O_7_0_0_0),
    .O_7_0_0_1(op_O_7_0_0_1),
    .O_7_0_0_2(op_O_7_0_0_2),
    .O_8_0_0_0(op_O_8_0_0_0),
    .O_8_0_0_1(op_O_8_0_0_1),
    .O_8_0_0_2(op_O_8_0_0_2),
    .O_9_0_0_0(op_O_9_0_0_0),
    .O_9_0_0_1(op_O_9_0_0_1),
    .O_9_0_0_2(op_O_9_0_0_2),
    .O_10_0_0_0(op_O_10_0_0_0),
    .O_10_0_0_1(op_O_10_0_0_1),
    .O_10_0_0_2(op_O_10_0_0_2),
    .O_11_0_0_0(op_O_11_0_0_0),
    .O_11_0_0_1(op_O_11_0_0_1),
    .O_11_0_0_2(op_O_11_0_0_2),
    .O_12_0_0_0(op_O_12_0_0_0),
    .O_12_0_0_1(op_O_12_0_0_1),
    .O_12_0_0_2(op_O_12_0_0_2),
    .O_13_0_0_0(op_O_13_0_0_0),
    .O_13_0_0_1(op_O_13_0_0_1),
    .O_13_0_0_2(op_O_13_0_0_2),
    .O_14_0_0_0(op_O_14_0_0_0),
    .O_14_0_0_1(op_O_14_0_0_1),
    .O_14_0_0_2(op_O_14_0_0_2),
    .O_15_0_0_0(op_O_15_0_0_0),
    .O_15_0_0_1(op_O_15_0_0_1),
    .O_15_0_0_2(op_O_15_0_0_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_0_2 = op_O_0_0_0_2; // @[Map2T.scala 17:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_0_2 = op_O_1_0_0_2; // @[Map2T.scala 17:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_0_2 = op_O_2_0_0_2; // @[Map2T.scala 17:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_0_2 = op_O_3_0_0_2; // @[Map2T.scala 17:7]
  assign O_4_0_0_0 = op_O_4_0_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_0_1 = op_O_4_0_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_0_2 = op_O_4_0_0_2; // @[Map2T.scala 17:7]
  assign O_5_0_0_0 = op_O_5_0_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_0_1 = op_O_5_0_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_0_2 = op_O_5_0_0_2; // @[Map2T.scala 17:7]
  assign O_6_0_0_0 = op_O_6_0_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_0_1 = op_O_6_0_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_0_2 = op_O_6_0_0_2; // @[Map2T.scala 17:7]
  assign O_7_0_0_0 = op_O_7_0_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_0_1 = op_O_7_0_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_0_2 = op_O_7_0_0_2; // @[Map2T.scala 17:7]
  assign O_8_0_0_0 = op_O_8_0_0_0; // @[Map2T.scala 17:7]
  assign O_8_0_0_1 = op_O_8_0_0_1; // @[Map2T.scala 17:7]
  assign O_8_0_0_2 = op_O_8_0_0_2; // @[Map2T.scala 17:7]
  assign O_9_0_0_0 = op_O_9_0_0_0; // @[Map2T.scala 17:7]
  assign O_9_0_0_1 = op_O_9_0_0_1; // @[Map2T.scala 17:7]
  assign O_9_0_0_2 = op_O_9_0_0_2; // @[Map2T.scala 17:7]
  assign O_10_0_0_0 = op_O_10_0_0_0; // @[Map2T.scala 17:7]
  assign O_10_0_0_1 = op_O_10_0_0_1; // @[Map2T.scala 17:7]
  assign O_10_0_0_2 = op_O_10_0_0_2; // @[Map2T.scala 17:7]
  assign O_11_0_0_0 = op_O_11_0_0_0; // @[Map2T.scala 17:7]
  assign O_11_0_0_1 = op_O_11_0_0_1; // @[Map2T.scala 17:7]
  assign O_11_0_0_2 = op_O_11_0_0_2; // @[Map2T.scala 17:7]
  assign O_12_0_0_0 = op_O_12_0_0_0; // @[Map2T.scala 17:7]
  assign O_12_0_0_1 = op_O_12_0_0_1; // @[Map2T.scala 17:7]
  assign O_12_0_0_2 = op_O_12_0_0_2; // @[Map2T.scala 17:7]
  assign O_13_0_0_0 = op_O_13_0_0_0; // @[Map2T.scala 17:7]
  assign O_13_0_0_1 = op_O_13_0_0_1; // @[Map2T.scala 17:7]
  assign O_13_0_0_2 = op_O_13_0_0_2; // @[Map2T.scala 17:7]
  assign O_14_0_0_0 = op_O_14_0_0_0; // @[Map2T.scala 17:7]
  assign O_14_0_0_1 = op_O_14_0_0_1; // @[Map2T.scala 17:7]
  assign O_14_0_0_2 = op_O_14_0_0_2; // @[Map2T.scala 17:7]
  assign O_15_0_0_0 = op_O_15_0_0_0; // @[Map2T.scala 17:7]
  assign O_15_0_0_1 = op_O_15_0_0_1; // @[Map2T.scala 17:7]
  assign O_15_0_0_2 = op_O_15_0_0_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0_0 = I0_0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_0_1 = I0_0_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0_0 = I0_1_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0_1 = I0_1_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0_0 = I0_2_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0_1 = I0_2_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0_0 = I0_3_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0_1 = I0_3_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0_0 = I0_4_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0_1 = I0_4_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0_0 = I0_5_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0_1 = I0_5_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0_0 = I0_6_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0_1 = I0_6_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0_0 = I0_7_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0_1 = I0_7_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_8_0_0_0 = I0_8_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_8_0_0_1 = I0_8_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_9_0_0_0 = I0_9_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_9_0_0_1 = I0_9_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_10_0_0_0 = I0_10_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_10_0_0_1 = I0_10_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_11_0_0_0 = I0_11_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_11_0_0_1 = I0_11_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_12_0_0_0 = I0_12_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_12_0_0_1 = I0_12_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_13_0_0_0 = I0_13_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_13_0_0_1 = I0_13_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_14_0_0_0 = I0_14_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_14_0_0_1 = I0_14_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_15_0_0_0 = I0_15_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_15_0_0_1 = I0_15_0_0_1; // @[Map2T.scala 15:11]
  assign op_I1_0_0_0 = I1_0_0_0; // @[Map2T.scala 16:11]
  assign op_I1_1_0_0 = I1_1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_2_0_0 = I1_2_0_0; // @[Map2T.scala 16:11]
  assign op_I1_3_0_0 = I1_3_0_0; // @[Map2T.scala 16:11]
  assign op_I1_4_0_0 = I1_4_0_0; // @[Map2T.scala 16:11]
  assign op_I1_5_0_0 = I1_5_0_0; // @[Map2T.scala 16:11]
  assign op_I1_6_0_0 = I1_6_0_0; // @[Map2T.scala 16:11]
  assign op_I1_7_0_0 = I1_7_0_0; // @[Map2T.scala 16:11]
  assign op_I1_8_0_0 = I1_8_0_0; // @[Map2T.scala 16:11]
  assign op_I1_9_0_0 = I1_9_0_0; // @[Map2T.scala 16:11]
  assign op_I1_10_0_0 = I1_10_0_0; // @[Map2T.scala 16:11]
  assign op_I1_11_0_0 = I1_11_0_0; // @[Map2T.scala 16:11]
  assign op_I1_12_0_0 = I1_12_0_0; // @[Map2T.scala 16:11]
  assign op_I1_13_0_0 = I1_13_0_0; // @[Map2T.scala 16:11]
  assign op_I1_14_0_0 = I1_14_0_0; // @[Map2T.scala 16:11]
  assign op_I1_15_0_0 = I1_15_0_0; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleToSSeq(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0 = I_0; // @[Tuple.scala 41:5]
  assign O_1 = I_1; // @[Tuple.scala 41:5]
  assign O_2 = I_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0(op_inst_I_0),
    .I_1(op_inst_I_1),
    .I_2(op_inst_I_2),
    .O_0(op_inst_O_0),
    .O_1(op_inst_O_1),
    .O_2(op_inst_O_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0 = op_inst_O_0; // @[Remove1S.scala 14:5]
  assign O_1 = op_inst_O_1; // @[Remove1S.scala 14:5]
  assign O_2 = op_inst_O_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0 = I_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1 = I_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2 = I_0_2; // @[Remove1S.scala 13:13]
endmodule
module MapS(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2; // @[MapS.scala 9:22]
  Remove1S fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
endmodule
module MapS_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0_0,
  input  [7:0] I_0_0_0_1,
  input  [7:0] I_0_0_0_2,
  input  [7:0] I_1_0_0_0,
  input  [7:0] I_1_0_0_1,
  input  [7:0] I_1_0_0_2,
  input  [7:0] I_2_0_0_0,
  input  [7:0] I_2_0_0_1,
  input  [7:0] I_2_0_0_2,
  input  [7:0] I_3_0_0_0,
  input  [7:0] I_3_0_0_1,
  input  [7:0] I_3_0_0_2,
  input  [7:0] I_4_0_0_0,
  input  [7:0] I_4_0_0_1,
  input  [7:0] I_4_0_0_2,
  input  [7:0] I_5_0_0_0,
  input  [7:0] I_5_0_0_1,
  input  [7:0] I_5_0_0_2,
  input  [7:0] I_6_0_0_0,
  input  [7:0] I_6_0_0_1,
  input  [7:0] I_6_0_0_2,
  input  [7:0] I_7_0_0_0,
  input  [7:0] I_7_0_0_1,
  input  [7:0] I_7_0_0_2,
  input  [7:0] I_8_0_0_0,
  input  [7:0] I_8_0_0_1,
  input  [7:0] I_8_0_0_2,
  input  [7:0] I_9_0_0_0,
  input  [7:0] I_9_0_0_1,
  input  [7:0] I_9_0_0_2,
  input  [7:0] I_10_0_0_0,
  input  [7:0] I_10_0_0_1,
  input  [7:0] I_10_0_0_2,
  input  [7:0] I_11_0_0_0,
  input  [7:0] I_11_0_0_1,
  input  [7:0] I_11_0_0_2,
  input  [7:0] I_12_0_0_0,
  input  [7:0] I_12_0_0_1,
  input  [7:0] I_12_0_0_2,
  input  [7:0] I_13_0_0_0,
  input  [7:0] I_13_0_0_1,
  input  [7:0] I_13_0_0_2,
  input  [7:0] I_14_0_0_0,
  input  [7:0] I_14_0_0_1,
  input  [7:0] I_14_0_0_2,
  input  [7:0] I_15_0_0_0,
  input  [7:0] I_15_0_0_1,
  input  [7:0] I_15_0_0_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_2; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  MapS fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0_0(fst_op_I_0_0_0),
    .I_0_0_1(fst_op_I_0_0_1),
    .I_0_0_2(fst_op_I_0_0_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2)
  );
  MapS other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0_0(other_ops_0_I_0_0_0),
    .I_0_0_1(other_ops_0_I_0_0_1),
    .I_0_0_2(other_ops_0_I_0_0_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2)
  );
  MapS other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0_0(other_ops_1_I_0_0_0),
    .I_0_0_1(other_ops_1_I_0_0_1),
    .I_0_0_2(other_ops_1_I_0_0_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2)
  );
  MapS other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0_0(other_ops_2_I_0_0_0),
    .I_0_0_1(other_ops_2_I_0_0_1),
    .I_0_0_2(other_ops_2_I_0_0_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2)
  );
  MapS other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0_0(other_ops_3_I_0_0_0),
    .I_0_0_1(other_ops_3_I_0_0_1),
    .I_0_0_2(other_ops_3_I_0_0_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2)
  );
  MapS other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0_0(other_ops_4_I_0_0_0),
    .I_0_0_1(other_ops_4_I_0_0_1),
    .I_0_0_2(other_ops_4_I_0_0_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2)
  );
  MapS other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0_0(other_ops_5_I_0_0_0),
    .I_0_0_1(other_ops_5_I_0_0_1),
    .I_0_0_2(other_ops_5_I_0_0_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2)
  );
  MapS other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0_0(other_ops_6_I_0_0_0),
    .I_0_0_1(other_ops_6_I_0_0_1),
    .I_0_0_2(other_ops_6_I_0_0_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2)
  );
  MapS other_ops_7 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0_0(other_ops_7_I_0_0_0),
    .I_0_0_1(other_ops_7_I_0_0_1),
    .I_0_0_2(other_ops_7_I_0_0_2),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_0_2(other_ops_7_O_0_2)
  );
  MapS other_ops_8 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0_0(other_ops_8_I_0_0_0),
    .I_0_0_1(other_ops_8_I_0_0_1),
    .I_0_0_2(other_ops_8_I_0_0_2),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_0_2(other_ops_8_O_0_2)
  );
  MapS other_ops_9 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0_0(other_ops_9_I_0_0_0),
    .I_0_0_1(other_ops_9_I_0_0_1),
    .I_0_0_2(other_ops_9_I_0_0_2),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_0_2(other_ops_9_O_0_2)
  );
  MapS other_ops_10 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0_0(other_ops_10_I_0_0_0),
    .I_0_0_1(other_ops_10_I_0_0_1),
    .I_0_0_2(other_ops_10_I_0_0_2),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_0_2(other_ops_10_O_0_2)
  );
  MapS other_ops_11 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0_0(other_ops_11_I_0_0_0),
    .I_0_0_1(other_ops_11_I_0_0_1),
    .I_0_0_2(other_ops_11_I_0_0_2),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_0_2(other_ops_11_O_0_2)
  );
  MapS other_ops_12 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0_0(other_ops_12_I_0_0_0),
    .I_0_0_1(other_ops_12_I_0_0_1),
    .I_0_0_2(other_ops_12_I_0_0_2),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_0_2(other_ops_12_O_0_2)
  );
  MapS other_ops_13 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0_0(other_ops_13_I_0_0_0),
    .I_0_0_1(other_ops_13_I_0_0_1),
    .I_0_0_2(other_ops_13_I_0_0_2),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_0_2(other_ops_13_O_0_2)
  );
  MapS other_ops_14 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0_0(other_ops_14_I_0_0_0),
    .I_0_0_1(other_ops_14_I_0_0_1),
    .I_0_0_2(other_ops_14_I_0_0_2),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_0_2(other_ops_14_O_0_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[MapS.scala 17:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[MapS.scala 21:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[MapS.scala 21:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[MapS.scala 21:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[MapS.scala 21:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[MapS.scala 21:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[MapS.scala 21:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[MapS.scala 21:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[MapS.scala 21:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[MapS.scala 21:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[MapS.scala 21:12]
  assign O_8_0_2 = other_ops_7_O_0_2; // @[MapS.scala 21:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[MapS.scala 21:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[MapS.scala 21:12]
  assign O_9_0_2 = other_ops_8_O_0_2; // @[MapS.scala 21:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[MapS.scala 21:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[MapS.scala 21:12]
  assign O_10_0_2 = other_ops_9_O_0_2; // @[MapS.scala 21:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[MapS.scala 21:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[MapS.scala 21:12]
  assign O_11_0_2 = other_ops_10_O_0_2; // @[MapS.scala 21:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[MapS.scala 21:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[MapS.scala 21:12]
  assign O_12_0_2 = other_ops_11_O_0_2; // @[MapS.scala 21:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[MapS.scala 21:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[MapS.scala 21:12]
  assign O_13_0_2 = other_ops_12_O_0_2; // @[MapS.scala 21:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[MapS.scala 21:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[MapS.scala 21:12]
  assign O_14_0_2 = other_ops_13_O_0_2; // @[MapS.scala 21:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[MapS.scala 21:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[MapS.scala 21:12]
  assign O_15_0_2 = other_ops_14_O_0_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0_0 = I_0_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_1 = I_0_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_2 = I_0_0_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0_0 = I_1_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_1 = I_1_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_2 = I_1_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0_0 = I_2_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_1 = I_2_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_2 = I_2_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0_0 = I_3_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_1 = I_3_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_2 = I_3_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0_0 = I_4_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_1 = I_4_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_2 = I_4_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0_0 = I_5_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_1 = I_5_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_2 = I_5_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0_0 = I_6_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_1 = I_6_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_2 = I_6_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0_0 = I_7_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_1 = I_7_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_2 = I_7_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0_0 = I_8_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_0_1 = I_8_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_0_2 = I_8_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0_0 = I_9_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_0_1 = I_9_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_0_2 = I_9_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0_0 = I_10_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_0_1 = I_10_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_0_2 = I_10_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0_0 = I_11_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_0_1 = I_11_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_0_2 = I_11_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0_0 = I_12_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_0_1 = I_12_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_0_2 = I_12_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0_0 = I_13_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_0_1 = I_13_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_0_2 = I_13_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0_0 = I_14_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_0_1 = I_14_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_0_2 = I_14_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0_0 = I_15_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_0_1 = I_15_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_0_2 = I_15_0_0_2; // @[MapS.scala 20:41]
endmodule
module MapT(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0_0,
  input  [7:0] I_0_0_0_1,
  input  [7:0] I_0_0_0_2,
  input  [7:0] I_1_0_0_0,
  input  [7:0] I_1_0_0_1,
  input  [7:0] I_1_0_0_2,
  input  [7:0] I_2_0_0_0,
  input  [7:0] I_2_0_0_1,
  input  [7:0] I_2_0_0_2,
  input  [7:0] I_3_0_0_0,
  input  [7:0] I_3_0_0_1,
  input  [7:0] I_3_0_0_2,
  input  [7:0] I_4_0_0_0,
  input  [7:0] I_4_0_0_1,
  input  [7:0] I_4_0_0_2,
  input  [7:0] I_5_0_0_0,
  input  [7:0] I_5_0_0_1,
  input  [7:0] I_5_0_0_2,
  input  [7:0] I_6_0_0_0,
  input  [7:0] I_6_0_0_1,
  input  [7:0] I_6_0_0_2,
  input  [7:0] I_7_0_0_0,
  input  [7:0] I_7_0_0_1,
  input  [7:0] I_7_0_0_2,
  input  [7:0] I_8_0_0_0,
  input  [7:0] I_8_0_0_1,
  input  [7:0] I_8_0_0_2,
  input  [7:0] I_9_0_0_0,
  input  [7:0] I_9_0_0_1,
  input  [7:0] I_9_0_0_2,
  input  [7:0] I_10_0_0_0,
  input  [7:0] I_10_0_0_1,
  input  [7:0] I_10_0_0_2,
  input  [7:0] I_11_0_0_0,
  input  [7:0] I_11_0_0_1,
  input  [7:0] I_11_0_0_2,
  input  [7:0] I_12_0_0_0,
  input  [7:0] I_12_0_0_1,
  input  [7:0] I_12_0_0_2,
  input  [7:0] I_13_0_0_0,
  input  [7:0] I_13_0_0_1,
  input  [7:0] I_13_0_0_2,
  input  [7:0] I_14_0_0_0,
  input  [7:0] I_14_0_0_1,
  input  [7:0] I_14_0_0_2,
  input  [7:0] I_15_0_0_0,
  input  [7:0] I_15_0_0_1,
  input  [7:0] I_15_0_0_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_2; // @[MapT.scala 8:20]
  MapS_1 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0_0(op_I_0_0_0_0),
    .I_0_0_0_1(op_I_0_0_0_1),
    .I_0_0_0_2(op_I_0_0_0_2),
    .I_1_0_0_0(op_I_1_0_0_0),
    .I_1_0_0_1(op_I_1_0_0_1),
    .I_1_0_0_2(op_I_1_0_0_2),
    .I_2_0_0_0(op_I_2_0_0_0),
    .I_2_0_0_1(op_I_2_0_0_1),
    .I_2_0_0_2(op_I_2_0_0_2),
    .I_3_0_0_0(op_I_3_0_0_0),
    .I_3_0_0_1(op_I_3_0_0_1),
    .I_3_0_0_2(op_I_3_0_0_2),
    .I_4_0_0_0(op_I_4_0_0_0),
    .I_4_0_0_1(op_I_4_0_0_1),
    .I_4_0_0_2(op_I_4_0_0_2),
    .I_5_0_0_0(op_I_5_0_0_0),
    .I_5_0_0_1(op_I_5_0_0_1),
    .I_5_0_0_2(op_I_5_0_0_2),
    .I_6_0_0_0(op_I_6_0_0_0),
    .I_6_0_0_1(op_I_6_0_0_1),
    .I_6_0_0_2(op_I_6_0_0_2),
    .I_7_0_0_0(op_I_7_0_0_0),
    .I_7_0_0_1(op_I_7_0_0_1),
    .I_7_0_0_2(op_I_7_0_0_2),
    .I_8_0_0_0(op_I_8_0_0_0),
    .I_8_0_0_1(op_I_8_0_0_1),
    .I_8_0_0_2(op_I_8_0_0_2),
    .I_9_0_0_0(op_I_9_0_0_0),
    .I_9_0_0_1(op_I_9_0_0_1),
    .I_9_0_0_2(op_I_9_0_0_2),
    .I_10_0_0_0(op_I_10_0_0_0),
    .I_10_0_0_1(op_I_10_0_0_1),
    .I_10_0_0_2(op_I_10_0_0_2),
    .I_11_0_0_0(op_I_11_0_0_0),
    .I_11_0_0_1(op_I_11_0_0_1),
    .I_11_0_0_2(op_I_11_0_0_2),
    .I_12_0_0_0(op_I_12_0_0_0),
    .I_12_0_0_1(op_I_12_0_0_1),
    .I_12_0_0_2(op_I_12_0_0_2),
    .I_13_0_0_0(op_I_13_0_0_0),
    .I_13_0_0_1(op_I_13_0_0_1),
    .I_13_0_0_2(op_I_13_0_0_2),
    .I_14_0_0_0(op_I_14_0_0_0),
    .I_14_0_0_1(op_I_14_0_0_1),
    .I_14_0_0_2(op_I_14_0_0_2),
    .I_15_0_0_0(op_I_15_0_0_0),
    .I_15_0_0_1(op_I_15_0_0_1),
    .I_15_0_0_2(op_I_15_0_0_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_0_2(op_O_8_0_2),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_0_2(op_O_9_0_2),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_0_2(op_O_10_0_2),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_0_2(op_O_11_0_2),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_0_2(op_O_12_0_2),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_0_2(op_O_13_0_2),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_0_2(op_O_14_0_2),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_0_2(op_O_15_0_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_4_0_2 = op_O_4_0_2; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_5_0_2 = op_O_5_0_2; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_6_0_2 = op_O_6_0_2; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_7_0_2 = op_O_7_0_2; // @[MapT.scala 15:7]
  assign O_8_0_0 = op_O_8_0_0; // @[MapT.scala 15:7]
  assign O_8_0_1 = op_O_8_0_1; // @[MapT.scala 15:7]
  assign O_8_0_2 = op_O_8_0_2; // @[MapT.scala 15:7]
  assign O_9_0_0 = op_O_9_0_0; // @[MapT.scala 15:7]
  assign O_9_0_1 = op_O_9_0_1; // @[MapT.scala 15:7]
  assign O_9_0_2 = op_O_9_0_2; // @[MapT.scala 15:7]
  assign O_10_0_0 = op_O_10_0_0; // @[MapT.scala 15:7]
  assign O_10_0_1 = op_O_10_0_1; // @[MapT.scala 15:7]
  assign O_10_0_2 = op_O_10_0_2; // @[MapT.scala 15:7]
  assign O_11_0_0 = op_O_11_0_0; // @[MapT.scala 15:7]
  assign O_11_0_1 = op_O_11_0_1; // @[MapT.scala 15:7]
  assign O_11_0_2 = op_O_11_0_2; // @[MapT.scala 15:7]
  assign O_12_0_0 = op_O_12_0_0; // @[MapT.scala 15:7]
  assign O_12_0_1 = op_O_12_0_1; // @[MapT.scala 15:7]
  assign O_12_0_2 = op_O_12_0_2; // @[MapT.scala 15:7]
  assign O_13_0_0 = op_O_13_0_0; // @[MapT.scala 15:7]
  assign O_13_0_1 = op_O_13_0_1; // @[MapT.scala 15:7]
  assign O_13_0_2 = op_O_13_0_2; // @[MapT.scala 15:7]
  assign O_14_0_0 = op_O_14_0_0; // @[MapT.scala 15:7]
  assign O_14_0_1 = op_O_14_0_1; // @[MapT.scala 15:7]
  assign O_14_0_2 = op_O_14_0_2; // @[MapT.scala 15:7]
  assign O_15_0_0 = op_O_15_0_0; // @[MapT.scala 15:7]
  assign O_15_0_1 = op_O_15_0_1; // @[MapT.scala 15:7]
  assign O_15_0_2 = op_O_15_0_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0_0 = I_0_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_0_1 = I_0_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_0_2 = I_0_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0_0 = I_1_0_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_0_1 = I_1_0_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0_2 = I_1_0_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0_0 = I_2_0_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_0_1 = I_2_0_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0_2 = I_2_0_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0_0 = I_3_0_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_0_1 = I_3_0_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0_2 = I_3_0_0_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0_0 = I_4_0_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_0_1 = I_4_0_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_0_2 = I_4_0_0_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0_0 = I_5_0_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_0_1 = I_5_0_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_0_2 = I_5_0_0_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0_0 = I_6_0_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_0_1 = I_6_0_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_0_2 = I_6_0_0_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0_0 = I_7_0_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_0_1 = I_7_0_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_0_2 = I_7_0_0_2; // @[MapT.scala 14:10]
  assign op_I_8_0_0_0 = I_8_0_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_0_1 = I_8_0_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_0_2 = I_8_0_0_2; // @[MapT.scala 14:10]
  assign op_I_9_0_0_0 = I_9_0_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_0_1 = I_9_0_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_0_2 = I_9_0_0_2; // @[MapT.scala 14:10]
  assign op_I_10_0_0_0 = I_10_0_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_0_1 = I_10_0_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_0_2 = I_10_0_0_2; // @[MapT.scala 14:10]
  assign op_I_11_0_0_0 = I_11_0_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_0_1 = I_11_0_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_0_2 = I_11_0_0_2; // @[MapT.scala 14:10]
  assign op_I_12_0_0_0 = I_12_0_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_0_1 = I_12_0_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_0_2 = I_12_0_0_2; // @[MapT.scala 14:10]
  assign op_I_13_0_0_0 = I_13_0_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_0_1 = I_13_0_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_0_2 = I_13_0_0_2; // @[MapT.scala 14:10]
  assign op_I_14_0_0_0 = I_14_0_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_0_1 = I_14_0_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_0_2 = I_14_0_0_2; // @[MapT.scala 14:10]
  assign op_I_15_0_0_0 = I_15_0_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_0_1 = I_15_0_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_0_2 = I_15_0_0_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleCreator_2(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0_0 = I0_0; // @[Tuple.scala 12:32]
  assign O_0_1 = I0_1; // @[Tuple.scala 12:32]
  assign O_0_2 = I0_2; // @[Tuple.scala 12:32]
  assign O_1_0 = I1_0; // @[Tuple.scala 13:32]
  assign O_1_1 = I1_1; // @[Tuple.scala 13:32]
  assign O_1_2 = I1_2; // @[Tuple.scala 13:32]
endmodule
module Map2S_12(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_0_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  SSeqTupleCreator_2 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
endmodule
module Map2S_13(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_0_0_1,
  input  [7:0] I0_0_0_2,
  input  [7:0] I0_1_0_0,
  input  [7:0] I0_1_0_1,
  input  [7:0] I0_1_0_2,
  input  [7:0] I0_2_0_0,
  input  [7:0] I0_2_0_1,
  input  [7:0] I0_2_0_2,
  input  [7:0] I0_3_0_0,
  input  [7:0] I0_3_0_1,
  input  [7:0] I0_3_0_2,
  input  [7:0] I0_4_0_0,
  input  [7:0] I0_4_0_1,
  input  [7:0] I0_4_0_2,
  input  [7:0] I0_5_0_0,
  input  [7:0] I0_5_0_1,
  input  [7:0] I0_5_0_2,
  input  [7:0] I0_6_0_0,
  input  [7:0] I0_6_0_1,
  input  [7:0] I0_6_0_2,
  input  [7:0] I0_7_0_0,
  input  [7:0] I0_7_0_1,
  input  [7:0] I0_7_0_2,
  input  [7:0] I0_8_0_0,
  input  [7:0] I0_8_0_1,
  input  [7:0] I0_8_0_2,
  input  [7:0] I0_9_0_0,
  input  [7:0] I0_9_0_1,
  input  [7:0] I0_9_0_2,
  input  [7:0] I0_10_0_0,
  input  [7:0] I0_10_0_1,
  input  [7:0] I0_10_0_2,
  input  [7:0] I0_11_0_0,
  input  [7:0] I0_11_0_1,
  input  [7:0] I0_11_0_2,
  input  [7:0] I0_12_0_0,
  input  [7:0] I0_12_0_1,
  input  [7:0] I0_12_0_2,
  input  [7:0] I0_13_0_0,
  input  [7:0] I0_13_0_1,
  input  [7:0] I0_13_0_2,
  input  [7:0] I0_14_0_0,
  input  [7:0] I0_14_0_1,
  input  [7:0] I0_14_0_2,
  input  [7:0] I0_15_0_0,
  input  [7:0] I0_15_0_1,
  input  [7:0] I0_15_0_2,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_0_0_1,
  input  [7:0] I1_0_0_2,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_1_0_1,
  input  [7:0] I1_1_0_2,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_2_0_1,
  input  [7:0] I1_2_0_2,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_3_0_1,
  input  [7:0] I1_3_0_2,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_4_0_1,
  input  [7:0] I1_4_0_2,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_5_0_1,
  input  [7:0] I1_5_0_2,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_6_0_1,
  input  [7:0] I1_6_0_2,
  input  [7:0] I1_7_0_0,
  input  [7:0] I1_7_0_1,
  input  [7:0] I1_7_0_2,
  input  [7:0] I1_8_0_0,
  input  [7:0] I1_8_0_1,
  input  [7:0] I1_8_0_2,
  input  [7:0] I1_9_0_0,
  input  [7:0] I1_9_0_1,
  input  [7:0] I1_9_0_2,
  input  [7:0] I1_10_0_0,
  input  [7:0] I1_10_0_1,
  input  [7:0] I1_10_0_2,
  input  [7:0] I1_11_0_0,
  input  [7:0] I1_11_0_1,
  input  [7:0] I1_11_0_2,
  input  [7:0] I1_12_0_0,
  input  [7:0] I1_12_0_1,
  input  [7:0] I1_12_0_2,
  input  [7:0] I1_13_0_0,
  input  [7:0] I1_13_0_1,
  input  [7:0] I1_13_0_2,
  input  [7:0] I1_14_0_0,
  input  [7:0] I1_14_0_1,
  input  [7:0] I1_14_0_2,
  input  [7:0] I1_15_0_0,
  input  [7:0] I1_15_0_1,
  input  [7:0] I1_15_0_2,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_0_0_1_0,
  output [7:0] O_0_0_1_1,
  output [7:0] O_0_0_1_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_1_0_1_0,
  output [7:0] O_1_0_1_1,
  output [7:0] O_1_0_1_2,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_0_2,
  output [7:0] O_2_0_1_0,
  output [7:0] O_2_0_1_1,
  output [7:0] O_2_0_1_2,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_0_2,
  output [7:0] O_3_0_1_0,
  output [7:0] O_3_0_1_1,
  output [7:0] O_3_0_1_2,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_0_2,
  output [7:0] O_4_0_1_0,
  output [7:0] O_4_0_1_1,
  output [7:0] O_4_0_1_2,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_0_2,
  output [7:0] O_5_0_1_0,
  output [7:0] O_5_0_1_1,
  output [7:0] O_5_0_1_2,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_0_2,
  output [7:0] O_6_0_1_0,
  output [7:0] O_6_0_1_1,
  output [7:0] O_6_0_1_2,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_0_2,
  output [7:0] O_7_0_1_0,
  output [7:0] O_7_0_1_1,
  output [7:0] O_7_0_1_2,
  output [7:0] O_8_0_0_0,
  output [7:0] O_8_0_0_1,
  output [7:0] O_8_0_0_2,
  output [7:0] O_8_0_1_0,
  output [7:0] O_8_0_1_1,
  output [7:0] O_8_0_1_2,
  output [7:0] O_9_0_0_0,
  output [7:0] O_9_0_0_1,
  output [7:0] O_9_0_0_2,
  output [7:0] O_9_0_1_0,
  output [7:0] O_9_0_1_1,
  output [7:0] O_9_0_1_2,
  output [7:0] O_10_0_0_0,
  output [7:0] O_10_0_0_1,
  output [7:0] O_10_0_0_2,
  output [7:0] O_10_0_1_0,
  output [7:0] O_10_0_1_1,
  output [7:0] O_10_0_1_2,
  output [7:0] O_11_0_0_0,
  output [7:0] O_11_0_0_1,
  output [7:0] O_11_0_0_2,
  output [7:0] O_11_0_1_0,
  output [7:0] O_11_0_1_1,
  output [7:0] O_11_0_1_2,
  output [7:0] O_12_0_0_0,
  output [7:0] O_12_0_0_1,
  output [7:0] O_12_0_0_2,
  output [7:0] O_12_0_1_0,
  output [7:0] O_12_0_1_1,
  output [7:0] O_12_0_1_2,
  output [7:0] O_13_0_0_0,
  output [7:0] O_13_0_0_1,
  output [7:0] O_13_0_0_2,
  output [7:0] O_13_0_1_0,
  output [7:0] O_13_0_1_1,
  output [7:0] O_13_0_1_2,
  output [7:0] O_14_0_0_0,
  output [7:0] O_14_0_0_1,
  output [7:0] O_14_0_0_2,
  output [7:0] O_14_0_1_0,
  output [7:0] O_14_0_1_1,
  output [7:0] O_14_0_1_2,
  output [7:0] O_15_0_0_0,
  output [7:0] O_15_0_0_1,
  output [7:0] O_15_0_0_2,
  output [7:0] O_15_0_1_0,
  output [7:0] O_15_0_1_1,
  output [7:0] O_15_0_1_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_1_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  Map2S_12 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I1_0_0(fst_op_I1_0_0),
    .I1_0_1(fst_op_I1_0_1),
    .I1_0_2(fst_op_I1_0_2),
    .O_0_0_0(fst_op_O_0_0_0),
    .O_0_0_1(fst_op_O_0_0_1),
    .O_0_0_2(fst_op_O_0_0_2),
    .O_0_1_0(fst_op_O_0_1_0),
    .O_0_1_1(fst_op_O_0_1_1),
    .O_0_1_2(fst_op_O_0_1_2)
  );
  Map2S_12 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0(other_ops_0_I0_0_0),
    .I0_0_1(other_ops_0_I0_0_1),
    .I0_0_2(other_ops_0_I0_0_2),
    .I1_0_0(other_ops_0_I1_0_0),
    .I1_0_1(other_ops_0_I1_0_1),
    .I1_0_2(other_ops_0_I1_0_2),
    .O_0_0_0(other_ops_0_O_0_0_0),
    .O_0_0_1(other_ops_0_O_0_0_1),
    .O_0_0_2(other_ops_0_O_0_0_2),
    .O_0_1_0(other_ops_0_O_0_1_0),
    .O_0_1_1(other_ops_0_O_0_1_1),
    .O_0_1_2(other_ops_0_O_0_1_2)
  );
  Map2S_12 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0(other_ops_1_I0_0_0),
    .I0_0_1(other_ops_1_I0_0_1),
    .I0_0_2(other_ops_1_I0_0_2),
    .I1_0_0(other_ops_1_I1_0_0),
    .I1_0_1(other_ops_1_I1_0_1),
    .I1_0_2(other_ops_1_I1_0_2),
    .O_0_0_0(other_ops_1_O_0_0_0),
    .O_0_0_1(other_ops_1_O_0_0_1),
    .O_0_0_2(other_ops_1_O_0_0_2),
    .O_0_1_0(other_ops_1_O_0_1_0),
    .O_0_1_1(other_ops_1_O_0_1_1),
    .O_0_1_2(other_ops_1_O_0_1_2)
  );
  Map2S_12 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0(other_ops_2_I0_0_0),
    .I0_0_1(other_ops_2_I0_0_1),
    .I0_0_2(other_ops_2_I0_0_2),
    .I1_0_0(other_ops_2_I1_0_0),
    .I1_0_1(other_ops_2_I1_0_1),
    .I1_0_2(other_ops_2_I1_0_2),
    .O_0_0_0(other_ops_2_O_0_0_0),
    .O_0_0_1(other_ops_2_O_0_0_1),
    .O_0_0_2(other_ops_2_O_0_0_2),
    .O_0_1_0(other_ops_2_O_0_1_0),
    .O_0_1_1(other_ops_2_O_0_1_1),
    .O_0_1_2(other_ops_2_O_0_1_2)
  );
  Map2S_12 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0(other_ops_3_I0_0_0),
    .I0_0_1(other_ops_3_I0_0_1),
    .I0_0_2(other_ops_3_I0_0_2),
    .I1_0_0(other_ops_3_I1_0_0),
    .I1_0_1(other_ops_3_I1_0_1),
    .I1_0_2(other_ops_3_I1_0_2),
    .O_0_0_0(other_ops_3_O_0_0_0),
    .O_0_0_1(other_ops_3_O_0_0_1),
    .O_0_0_2(other_ops_3_O_0_0_2),
    .O_0_1_0(other_ops_3_O_0_1_0),
    .O_0_1_1(other_ops_3_O_0_1_1),
    .O_0_1_2(other_ops_3_O_0_1_2)
  );
  Map2S_12 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0(other_ops_4_I0_0_0),
    .I0_0_1(other_ops_4_I0_0_1),
    .I0_0_2(other_ops_4_I0_0_2),
    .I1_0_0(other_ops_4_I1_0_0),
    .I1_0_1(other_ops_4_I1_0_1),
    .I1_0_2(other_ops_4_I1_0_2),
    .O_0_0_0(other_ops_4_O_0_0_0),
    .O_0_0_1(other_ops_4_O_0_0_1),
    .O_0_0_2(other_ops_4_O_0_0_2),
    .O_0_1_0(other_ops_4_O_0_1_0),
    .O_0_1_1(other_ops_4_O_0_1_1),
    .O_0_1_2(other_ops_4_O_0_1_2)
  );
  Map2S_12 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0(other_ops_5_I0_0_0),
    .I0_0_1(other_ops_5_I0_0_1),
    .I0_0_2(other_ops_5_I0_0_2),
    .I1_0_0(other_ops_5_I1_0_0),
    .I1_0_1(other_ops_5_I1_0_1),
    .I1_0_2(other_ops_5_I1_0_2),
    .O_0_0_0(other_ops_5_O_0_0_0),
    .O_0_0_1(other_ops_5_O_0_0_1),
    .O_0_0_2(other_ops_5_O_0_0_2),
    .O_0_1_0(other_ops_5_O_0_1_0),
    .O_0_1_1(other_ops_5_O_0_1_1),
    .O_0_1_2(other_ops_5_O_0_1_2)
  );
  Map2S_12 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0(other_ops_6_I0_0_0),
    .I0_0_1(other_ops_6_I0_0_1),
    .I0_0_2(other_ops_6_I0_0_2),
    .I1_0_0(other_ops_6_I1_0_0),
    .I1_0_1(other_ops_6_I1_0_1),
    .I1_0_2(other_ops_6_I1_0_2),
    .O_0_0_0(other_ops_6_O_0_0_0),
    .O_0_0_1(other_ops_6_O_0_0_1),
    .O_0_0_2(other_ops_6_O_0_0_2),
    .O_0_1_0(other_ops_6_O_0_1_0),
    .O_0_1_1(other_ops_6_O_0_1_1),
    .O_0_1_2(other_ops_6_O_0_1_2)
  );
  Map2S_12 other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0_0(other_ops_7_I0_0_0),
    .I0_0_1(other_ops_7_I0_0_1),
    .I0_0_2(other_ops_7_I0_0_2),
    .I1_0_0(other_ops_7_I1_0_0),
    .I1_0_1(other_ops_7_I1_0_1),
    .I1_0_2(other_ops_7_I1_0_2),
    .O_0_0_0(other_ops_7_O_0_0_0),
    .O_0_0_1(other_ops_7_O_0_0_1),
    .O_0_0_2(other_ops_7_O_0_0_2),
    .O_0_1_0(other_ops_7_O_0_1_0),
    .O_0_1_1(other_ops_7_O_0_1_1),
    .O_0_1_2(other_ops_7_O_0_1_2)
  );
  Map2S_12 other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0_0(other_ops_8_I0_0_0),
    .I0_0_1(other_ops_8_I0_0_1),
    .I0_0_2(other_ops_8_I0_0_2),
    .I1_0_0(other_ops_8_I1_0_0),
    .I1_0_1(other_ops_8_I1_0_1),
    .I1_0_2(other_ops_8_I1_0_2),
    .O_0_0_0(other_ops_8_O_0_0_0),
    .O_0_0_1(other_ops_8_O_0_0_1),
    .O_0_0_2(other_ops_8_O_0_0_2),
    .O_0_1_0(other_ops_8_O_0_1_0),
    .O_0_1_1(other_ops_8_O_0_1_1),
    .O_0_1_2(other_ops_8_O_0_1_2)
  );
  Map2S_12 other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0_0(other_ops_9_I0_0_0),
    .I0_0_1(other_ops_9_I0_0_1),
    .I0_0_2(other_ops_9_I0_0_2),
    .I1_0_0(other_ops_9_I1_0_0),
    .I1_0_1(other_ops_9_I1_0_1),
    .I1_0_2(other_ops_9_I1_0_2),
    .O_0_0_0(other_ops_9_O_0_0_0),
    .O_0_0_1(other_ops_9_O_0_0_1),
    .O_0_0_2(other_ops_9_O_0_0_2),
    .O_0_1_0(other_ops_9_O_0_1_0),
    .O_0_1_1(other_ops_9_O_0_1_1),
    .O_0_1_2(other_ops_9_O_0_1_2)
  );
  Map2S_12 other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0_0(other_ops_10_I0_0_0),
    .I0_0_1(other_ops_10_I0_0_1),
    .I0_0_2(other_ops_10_I0_0_2),
    .I1_0_0(other_ops_10_I1_0_0),
    .I1_0_1(other_ops_10_I1_0_1),
    .I1_0_2(other_ops_10_I1_0_2),
    .O_0_0_0(other_ops_10_O_0_0_0),
    .O_0_0_1(other_ops_10_O_0_0_1),
    .O_0_0_2(other_ops_10_O_0_0_2),
    .O_0_1_0(other_ops_10_O_0_1_0),
    .O_0_1_1(other_ops_10_O_0_1_1),
    .O_0_1_2(other_ops_10_O_0_1_2)
  );
  Map2S_12 other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0_0(other_ops_11_I0_0_0),
    .I0_0_1(other_ops_11_I0_0_1),
    .I0_0_2(other_ops_11_I0_0_2),
    .I1_0_0(other_ops_11_I1_0_0),
    .I1_0_1(other_ops_11_I1_0_1),
    .I1_0_2(other_ops_11_I1_0_2),
    .O_0_0_0(other_ops_11_O_0_0_0),
    .O_0_0_1(other_ops_11_O_0_0_1),
    .O_0_0_2(other_ops_11_O_0_0_2),
    .O_0_1_0(other_ops_11_O_0_1_0),
    .O_0_1_1(other_ops_11_O_0_1_1),
    .O_0_1_2(other_ops_11_O_0_1_2)
  );
  Map2S_12 other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0_0(other_ops_12_I0_0_0),
    .I0_0_1(other_ops_12_I0_0_1),
    .I0_0_2(other_ops_12_I0_0_2),
    .I1_0_0(other_ops_12_I1_0_0),
    .I1_0_1(other_ops_12_I1_0_1),
    .I1_0_2(other_ops_12_I1_0_2),
    .O_0_0_0(other_ops_12_O_0_0_0),
    .O_0_0_1(other_ops_12_O_0_0_1),
    .O_0_0_2(other_ops_12_O_0_0_2),
    .O_0_1_0(other_ops_12_O_0_1_0),
    .O_0_1_1(other_ops_12_O_0_1_1),
    .O_0_1_2(other_ops_12_O_0_1_2)
  );
  Map2S_12 other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0_0(other_ops_13_I0_0_0),
    .I0_0_1(other_ops_13_I0_0_1),
    .I0_0_2(other_ops_13_I0_0_2),
    .I1_0_0(other_ops_13_I1_0_0),
    .I1_0_1(other_ops_13_I1_0_1),
    .I1_0_2(other_ops_13_I1_0_2),
    .O_0_0_0(other_ops_13_O_0_0_0),
    .O_0_0_1(other_ops_13_O_0_0_1),
    .O_0_0_2(other_ops_13_O_0_0_2),
    .O_0_1_0(other_ops_13_O_0_1_0),
    .O_0_1_1(other_ops_13_O_0_1_1),
    .O_0_1_2(other_ops_13_O_0_1_2)
  );
  Map2S_12 other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0_0(other_ops_14_I0_0_0),
    .I0_0_1(other_ops_14_I0_0_1),
    .I0_0_2(other_ops_14_I0_0_2),
    .I1_0_0(other_ops_14_I1_0_0),
    .I1_0_1(other_ops_14_I1_0_1),
    .I1_0_2(other_ops_14_I1_0_2),
    .O_0_0_0(other_ops_14_O_0_0_0),
    .O_0_0_1(other_ops_14_O_0_0_1),
    .O_0_0_2(other_ops_14_O_0_0_2),
    .O_0_1_0(other_ops_14_O_0_1_0),
    .O_0_1_1(other_ops_14_O_0_1_1),
    .O_0_1_2(other_ops_14_O_0_1_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0_0 = fst_op_O_0_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_0_1 = fst_op_O_0_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_0_2 = fst_op_O_0_0_2; // @[Map2S.scala 19:8]
  assign O_0_0_1_0 = fst_op_O_0_1_0; // @[Map2S.scala 19:8]
  assign O_0_0_1_1 = fst_op_O_0_1_1; // @[Map2S.scala 19:8]
  assign O_0_0_1_2 = fst_op_O_0_1_2; // @[Map2S.scala 19:8]
  assign O_1_0_0_0 = other_ops_0_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_0_1 = other_ops_0_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_0_2 = other_ops_0_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_1_0_1_0 = other_ops_0_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_1_0_1_1 = other_ops_0_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_1_0_1_2 = other_ops_0_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_2_0_0_0 = other_ops_1_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_0_1 = other_ops_1_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_0_2 = other_ops_1_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_2_0_1_0 = other_ops_1_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_2_0_1_1 = other_ops_1_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_2_0_1_2 = other_ops_1_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_3_0_0_0 = other_ops_2_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_0_1 = other_ops_2_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_0_2 = other_ops_2_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_3_0_1_0 = other_ops_2_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_3_0_1_1 = other_ops_2_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_3_0_1_2 = other_ops_2_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_4_0_0_0 = other_ops_3_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_0_1 = other_ops_3_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_0_2 = other_ops_3_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_4_0_1_0 = other_ops_3_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_4_0_1_1 = other_ops_3_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_4_0_1_2 = other_ops_3_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_5_0_0_0 = other_ops_4_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_0_1 = other_ops_4_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_0_2 = other_ops_4_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_5_0_1_0 = other_ops_4_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_5_0_1_1 = other_ops_4_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_5_0_1_2 = other_ops_4_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_6_0_0_0 = other_ops_5_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_0_1 = other_ops_5_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_0_2 = other_ops_5_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_6_0_1_0 = other_ops_5_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_6_0_1_1 = other_ops_5_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_6_0_1_2 = other_ops_5_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_7_0_0_0 = other_ops_6_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_0_1 = other_ops_6_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_0_2 = other_ops_6_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_7_0_1_0 = other_ops_6_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_7_0_1_1 = other_ops_6_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_7_0_1_2 = other_ops_6_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_8_0_0_0 = other_ops_7_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_8_0_0_1 = other_ops_7_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_8_0_0_2 = other_ops_7_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_8_0_1_0 = other_ops_7_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_8_0_1_1 = other_ops_7_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_8_0_1_2 = other_ops_7_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_9_0_0_0 = other_ops_8_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_9_0_0_1 = other_ops_8_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_9_0_0_2 = other_ops_8_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_9_0_1_0 = other_ops_8_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_9_0_1_1 = other_ops_8_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_9_0_1_2 = other_ops_8_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_10_0_0_0 = other_ops_9_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_10_0_0_1 = other_ops_9_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_10_0_0_2 = other_ops_9_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_10_0_1_0 = other_ops_9_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_10_0_1_1 = other_ops_9_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_10_0_1_2 = other_ops_9_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_11_0_0_0 = other_ops_10_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_11_0_0_1 = other_ops_10_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_11_0_0_2 = other_ops_10_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_11_0_1_0 = other_ops_10_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_11_0_1_1 = other_ops_10_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_11_0_1_2 = other_ops_10_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_12_0_0_0 = other_ops_11_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_12_0_0_1 = other_ops_11_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_12_0_0_2 = other_ops_11_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_12_0_1_0 = other_ops_11_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_12_0_1_1 = other_ops_11_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_12_0_1_2 = other_ops_11_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_13_0_0_0 = other_ops_12_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_13_0_0_1 = other_ops_12_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_13_0_0_2 = other_ops_12_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_13_0_1_0 = other_ops_12_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_13_0_1_1 = other_ops_12_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_13_0_1_2 = other_ops_12_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_14_0_0_0 = other_ops_13_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_14_0_0_1 = other_ops_13_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_14_0_0_2 = other_ops_13_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_14_0_1_0 = other_ops_13_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_14_0_1_1 = other_ops_13_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_14_0_1_2 = other_ops_13_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_15_0_0_0 = other_ops_14_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_15_0_0_1 = other_ops_14_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_15_0_0_2 = other_ops_14_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_15_0_1_0 = other_ops_14_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_15_0_1_1 = other_ops_14_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_15_0_1_2 = other_ops_14_O_0_1_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_0 = I1_0_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_1 = I1_0_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_2 = I1_0_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0 = I0_1_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1 = I0_1_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_2 = I0_1_0_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0_0 = I1_1_0_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_0_1 = I1_1_0_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_0_2 = I1_1_0_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0 = I0_2_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1 = I0_2_0_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_2 = I0_2_0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0_0 = I1_2_0_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_0_1 = I1_2_0_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_0_2 = I1_2_0_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0 = I0_3_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1 = I0_3_0_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_2 = I0_3_0_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0_0 = I1_3_0_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_0_1 = I1_3_0_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_0_2 = I1_3_0_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0 = I0_4_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1 = I0_4_0_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_2 = I0_4_0_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0_0 = I1_4_0_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_0_1 = I1_4_0_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_0_2 = I1_4_0_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0 = I0_5_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1 = I0_5_0_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_2 = I0_5_0_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0_0 = I1_5_0_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_0_1 = I1_5_0_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_0_2 = I1_5_0_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0 = I0_6_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1 = I0_6_0_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_2 = I0_6_0_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0_0 = I1_6_0_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_0_1 = I1_6_0_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_0_2 = I1_6_0_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0 = I0_7_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1 = I0_7_0_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_2 = I0_7_0_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0_0 = I1_7_0_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_0_1 = I1_7_0_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_0_2 = I1_7_0_2; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0_0 = I0_8_0_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_1 = I0_8_0_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_2 = I0_8_0_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I1_0_0 = I1_8_0_0; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_0_1 = I1_8_0_1; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_0_2 = I1_8_0_2; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0_0 = I0_9_0_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_1 = I0_9_0_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_2 = I0_9_0_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I1_0_0 = I1_9_0_0; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_0_1 = I1_9_0_1; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_0_2 = I1_9_0_2; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0_0 = I0_10_0_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_1 = I0_10_0_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_2 = I0_10_0_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I1_0_0 = I1_10_0_0; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_0_1 = I1_10_0_1; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_0_2 = I1_10_0_2; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0_0 = I0_11_0_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_1 = I0_11_0_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_2 = I0_11_0_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I1_0_0 = I1_11_0_0; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_0_1 = I1_11_0_1; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_0_2 = I1_11_0_2; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0_0 = I0_12_0_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_1 = I0_12_0_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_2 = I0_12_0_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I1_0_0 = I1_12_0_0; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_0_1 = I1_12_0_1; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_0_2 = I1_12_0_2; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0_0 = I0_13_0_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_1 = I0_13_0_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_2 = I0_13_0_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I1_0_0 = I1_13_0_0; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_0_1 = I1_13_0_1; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_0_2 = I1_13_0_2; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0_0 = I0_14_0_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_1 = I0_14_0_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_2 = I0_14_0_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I1_0_0 = I1_14_0_0; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_0_1 = I1_14_0_1; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_0_2 = I1_14_0_2; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0_0 = I0_15_0_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_1 = I0_15_0_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_2 = I0_15_0_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I1_0_0 = I1_15_0_0; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_0_1 = I1_15_0_1; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_0_2 = I1_15_0_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_0_0_1,
  input  [7:0] I0_0_0_2,
  input  [7:0] I0_1_0_0,
  input  [7:0] I0_1_0_1,
  input  [7:0] I0_1_0_2,
  input  [7:0] I0_2_0_0,
  input  [7:0] I0_2_0_1,
  input  [7:0] I0_2_0_2,
  input  [7:0] I0_3_0_0,
  input  [7:0] I0_3_0_1,
  input  [7:0] I0_3_0_2,
  input  [7:0] I0_4_0_0,
  input  [7:0] I0_4_0_1,
  input  [7:0] I0_4_0_2,
  input  [7:0] I0_5_0_0,
  input  [7:0] I0_5_0_1,
  input  [7:0] I0_5_0_2,
  input  [7:0] I0_6_0_0,
  input  [7:0] I0_6_0_1,
  input  [7:0] I0_6_0_2,
  input  [7:0] I0_7_0_0,
  input  [7:0] I0_7_0_1,
  input  [7:0] I0_7_0_2,
  input  [7:0] I0_8_0_0,
  input  [7:0] I0_8_0_1,
  input  [7:0] I0_8_0_2,
  input  [7:0] I0_9_0_0,
  input  [7:0] I0_9_0_1,
  input  [7:0] I0_9_0_2,
  input  [7:0] I0_10_0_0,
  input  [7:0] I0_10_0_1,
  input  [7:0] I0_10_0_2,
  input  [7:0] I0_11_0_0,
  input  [7:0] I0_11_0_1,
  input  [7:0] I0_11_0_2,
  input  [7:0] I0_12_0_0,
  input  [7:0] I0_12_0_1,
  input  [7:0] I0_12_0_2,
  input  [7:0] I0_13_0_0,
  input  [7:0] I0_13_0_1,
  input  [7:0] I0_13_0_2,
  input  [7:0] I0_14_0_0,
  input  [7:0] I0_14_0_1,
  input  [7:0] I0_14_0_2,
  input  [7:0] I0_15_0_0,
  input  [7:0] I0_15_0_1,
  input  [7:0] I0_15_0_2,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_0_0_1,
  input  [7:0] I1_0_0_2,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_1_0_1,
  input  [7:0] I1_1_0_2,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_2_0_1,
  input  [7:0] I1_2_0_2,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_3_0_1,
  input  [7:0] I1_3_0_2,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_4_0_1,
  input  [7:0] I1_4_0_2,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_5_0_1,
  input  [7:0] I1_5_0_2,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_6_0_1,
  input  [7:0] I1_6_0_2,
  input  [7:0] I1_7_0_0,
  input  [7:0] I1_7_0_1,
  input  [7:0] I1_7_0_2,
  input  [7:0] I1_8_0_0,
  input  [7:0] I1_8_0_1,
  input  [7:0] I1_8_0_2,
  input  [7:0] I1_9_0_0,
  input  [7:0] I1_9_0_1,
  input  [7:0] I1_9_0_2,
  input  [7:0] I1_10_0_0,
  input  [7:0] I1_10_0_1,
  input  [7:0] I1_10_0_2,
  input  [7:0] I1_11_0_0,
  input  [7:0] I1_11_0_1,
  input  [7:0] I1_11_0_2,
  input  [7:0] I1_12_0_0,
  input  [7:0] I1_12_0_1,
  input  [7:0] I1_12_0_2,
  input  [7:0] I1_13_0_0,
  input  [7:0] I1_13_0_1,
  input  [7:0] I1_13_0_2,
  input  [7:0] I1_14_0_0,
  input  [7:0] I1_14_0_1,
  input  [7:0] I1_14_0_2,
  input  [7:0] I1_15_0_0,
  input  [7:0] I1_15_0_1,
  input  [7:0] I1_15_0_2,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_0_0_1_0,
  output [7:0] O_0_0_1_1,
  output [7:0] O_0_0_1_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_1_0_1_0,
  output [7:0] O_1_0_1_1,
  output [7:0] O_1_0_1_2,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_0_2,
  output [7:0] O_2_0_1_0,
  output [7:0] O_2_0_1_1,
  output [7:0] O_2_0_1_2,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_0_2,
  output [7:0] O_3_0_1_0,
  output [7:0] O_3_0_1_1,
  output [7:0] O_3_0_1_2,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_0_2,
  output [7:0] O_4_0_1_0,
  output [7:0] O_4_0_1_1,
  output [7:0] O_4_0_1_2,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_0_2,
  output [7:0] O_5_0_1_0,
  output [7:0] O_5_0_1_1,
  output [7:0] O_5_0_1_2,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_0_2,
  output [7:0] O_6_0_1_0,
  output [7:0] O_6_0_1_1,
  output [7:0] O_6_0_1_2,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_0_2,
  output [7:0] O_7_0_1_0,
  output [7:0] O_7_0_1_1,
  output [7:0] O_7_0_1_2,
  output [7:0] O_8_0_0_0,
  output [7:0] O_8_0_0_1,
  output [7:0] O_8_0_0_2,
  output [7:0] O_8_0_1_0,
  output [7:0] O_8_0_1_1,
  output [7:0] O_8_0_1_2,
  output [7:0] O_9_0_0_0,
  output [7:0] O_9_0_0_1,
  output [7:0] O_9_0_0_2,
  output [7:0] O_9_0_1_0,
  output [7:0] O_9_0_1_1,
  output [7:0] O_9_0_1_2,
  output [7:0] O_10_0_0_0,
  output [7:0] O_10_0_0_1,
  output [7:0] O_10_0_0_2,
  output [7:0] O_10_0_1_0,
  output [7:0] O_10_0_1_1,
  output [7:0] O_10_0_1_2,
  output [7:0] O_11_0_0_0,
  output [7:0] O_11_0_0_1,
  output [7:0] O_11_0_0_2,
  output [7:0] O_11_0_1_0,
  output [7:0] O_11_0_1_1,
  output [7:0] O_11_0_1_2,
  output [7:0] O_12_0_0_0,
  output [7:0] O_12_0_0_1,
  output [7:0] O_12_0_0_2,
  output [7:0] O_12_0_1_0,
  output [7:0] O_12_0_1_1,
  output [7:0] O_12_0_1_2,
  output [7:0] O_13_0_0_0,
  output [7:0] O_13_0_0_1,
  output [7:0] O_13_0_0_2,
  output [7:0] O_13_0_1_0,
  output [7:0] O_13_0_1_1,
  output [7:0] O_13_0_1_2,
  output [7:0] O_14_0_0_0,
  output [7:0] O_14_0_0_1,
  output [7:0] O_14_0_0_2,
  output [7:0] O_14_0_1_0,
  output [7:0] O_14_0_1_1,
  output [7:0] O_14_0_1_2,
  output [7:0] O_15_0_0_0,
  output [7:0] O_15_0_0_1,
  output [7:0] O_15_0_0_2,
  output [7:0] O_15_0_1_0,
  output [7:0] O_15_0_1_1,
  output [7:0] O_15_0_1_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_1_2; // @[Map2T.scala 8:20]
  Map2S_13 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0(op_I0_0_0_0),
    .I0_0_0_1(op_I0_0_0_1),
    .I0_0_0_2(op_I0_0_0_2),
    .I0_1_0_0(op_I0_1_0_0),
    .I0_1_0_1(op_I0_1_0_1),
    .I0_1_0_2(op_I0_1_0_2),
    .I0_2_0_0(op_I0_2_0_0),
    .I0_2_0_1(op_I0_2_0_1),
    .I0_2_0_2(op_I0_2_0_2),
    .I0_3_0_0(op_I0_3_0_0),
    .I0_3_0_1(op_I0_3_0_1),
    .I0_3_0_2(op_I0_3_0_2),
    .I0_4_0_0(op_I0_4_0_0),
    .I0_4_0_1(op_I0_4_0_1),
    .I0_4_0_2(op_I0_4_0_2),
    .I0_5_0_0(op_I0_5_0_0),
    .I0_5_0_1(op_I0_5_0_1),
    .I0_5_0_2(op_I0_5_0_2),
    .I0_6_0_0(op_I0_6_0_0),
    .I0_6_0_1(op_I0_6_0_1),
    .I0_6_0_2(op_I0_6_0_2),
    .I0_7_0_0(op_I0_7_0_0),
    .I0_7_0_1(op_I0_7_0_1),
    .I0_7_0_2(op_I0_7_0_2),
    .I0_8_0_0(op_I0_8_0_0),
    .I0_8_0_1(op_I0_8_0_1),
    .I0_8_0_2(op_I0_8_0_2),
    .I0_9_0_0(op_I0_9_0_0),
    .I0_9_0_1(op_I0_9_0_1),
    .I0_9_0_2(op_I0_9_0_2),
    .I0_10_0_0(op_I0_10_0_0),
    .I0_10_0_1(op_I0_10_0_1),
    .I0_10_0_2(op_I0_10_0_2),
    .I0_11_0_0(op_I0_11_0_0),
    .I0_11_0_1(op_I0_11_0_1),
    .I0_11_0_2(op_I0_11_0_2),
    .I0_12_0_0(op_I0_12_0_0),
    .I0_12_0_1(op_I0_12_0_1),
    .I0_12_0_2(op_I0_12_0_2),
    .I0_13_0_0(op_I0_13_0_0),
    .I0_13_0_1(op_I0_13_0_1),
    .I0_13_0_2(op_I0_13_0_2),
    .I0_14_0_0(op_I0_14_0_0),
    .I0_14_0_1(op_I0_14_0_1),
    .I0_14_0_2(op_I0_14_0_2),
    .I0_15_0_0(op_I0_15_0_0),
    .I0_15_0_1(op_I0_15_0_1),
    .I0_15_0_2(op_I0_15_0_2),
    .I1_0_0_0(op_I1_0_0_0),
    .I1_0_0_1(op_I1_0_0_1),
    .I1_0_0_2(op_I1_0_0_2),
    .I1_1_0_0(op_I1_1_0_0),
    .I1_1_0_1(op_I1_1_0_1),
    .I1_1_0_2(op_I1_1_0_2),
    .I1_2_0_0(op_I1_2_0_0),
    .I1_2_0_1(op_I1_2_0_1),
    .I1_2_0_2(op_I1_2_0_2),
    .I1_3_0_0(op_I1_3_0_0),
    .I1_3_0_1(op_I1_3_0_1),
    .I1_3_0_2(op_I1_3_0_2),
    .I1_4_0_0(op_I1_4_0_0),
    .I1_4_0_1(op_I1_4_0_1),
    .I1_4_0_2(op_I1_4_0_2),
    .I1_5_0_0(op_I1_5_0_0),
    .I1_5_0_1(op_I1_5_0_1),
    .I1_5_0_2(op_I1_5_0_2),
    .I1_6_0_0(op_I1_6_0_0),
    .I1_6_0_1(op_I1_6_0_1),
    .I1_6_0_2(op_I1_6_0_2),
    .I1_7_0_0(op_I1_7_0_0),
    .I1_7_0_1(op_I1_7_0_1),
    .I1_7_0_2(op_I1_7_0_2),
    .I1_8_0_0(op_I1_8_0_0),
    .I1_8_0_1(op_I1_8_0_1),
    .I1_8_0_2(op_I1_8_0_2),
    .I1_9_0_0(op_I1_9_0_0),
    .I1_9_0_1(op_I1_9_0_1),
    .I1_9_0_2(op_I1_9_0_2),
    .I1_10_0_0(op_I1_10_0_0),
    .I1_10_0_1(op_I1_10_0_1),
    .I1_10_0_2(op_I1_10_0_2),
    .I1_11_0_0(op_I1_11_0_0),
    .I1_11_0_1(op_I1_11_0_1),
    .I1_11_0_2(op_I1_11_0_2),
    .I1_12_0_0(op_I1_12_0_0),
    .I1_12_0_1(op_I1_12_0_1),
    .I1_12_0_2(op_I1_12_0_2),
    .I1_13_0_0(op_I1_13_0_0),
    .I1_13_0_1(op_I1_13_0_1),
    .I1_13_0_2(op_I1_13_0_2),
    .I1_14_0_0(op_I1_14_0_0),
    .I1_14_0_1(op_I1_14_0_1),
    .I1_14_0_2(op_I1_14_0_2),
    .I1_15_0_0(op_I1_15_0_0),
    .I1_15_0_1(op_I1_15_0_1),
    .I1_15_0_2(op_I1_15_0_2),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_0_0_0_2(op_O_0_0_0_2),
    .O_0_0_1_0(op_O_0_0_1_0),
    .O_0_0_1_1(op_O_0_0_1_1),
    .O_0_0_1_2(op_O_0_0_1_2),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_1_0_0_2(op_O_1_0_0_2),
    .O_1_0_1_0(op_O_1_0_1_0),
    .O_1_0_1_1(op_O_1_0_1_1),
    .O_1_0_1_2(op_O_1_0_1_2),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_2_0_0_2(op_O_2_0_0_2),
    .O_2_0_1_0(op_O_2_0_1_0),
    .O_2_0_1_1(op_O_2_0_1_1),
    .O_2_0_1_2(op_O_2_0_1_2),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_3_0_0_2(op_O_3_0_0_2),
    .O_3_0_1_0(op_O_3_0_1_0),
    .O_3_0_1_1(op_O_3_0_1_1),
    .O_3_0_1_2(op_O_3_0_1_2),
    .O_4_0_0_0(op_O_4_0_0_0),
    .O_4_0_0_1(op_O_4_0_0_1),
    .O_4_0_0_2(op_O_4_0_0_2),
    .O_4_0_1_0(op_O_4_0_1_0),
    .O_4_0_1_1(op_O_4_0_1_1),
    .O_4_0_1_2(op_O_4_0_1_2),
    .O_5_0_0_0(op_O_5_0_0_0),
    .O_5_0_0_1(op_O_5_0_0_1),
    .O_5_0_0_2(op_O_5_0_0_2),
    .O_5_0_1_0(op_O_5_0_1_0),
    .O_5_0_1_1(op_O_5_0_1_1),
    .O_5_0_1_2(op_O_5_0_1_2),
    .O_6_0_0_0(op_O_6_0_0_0),
    .O_6_0_0_1(op_O_6_0_0_1),
    .O_6_0_0_2(op_O_6_0_0_2),
    .O_6_0_1_0(op_O_6_0_1_0),
    .O_6_0_1_1(op_O_6_0_1_1),
    .O_6_0_1_2(op_O_6_0_1_2),
    .O_7_0_0_0(op_O_7_0_0_0),
    .O_7_0_0_1(op_O_7_0_0_1),
    .O_7_0_0_2(op_O_7_0_0_2),
    .O_7_0_1_0(op_O_7_0_1_0),
    .O_7_0_1_1(op_O_7_0_1_1),
    .O_7_0_1_2(op_O_7_0_1_2),
    .O_8_0_0_0(op_O_8_0_0_0),
    .O_8_0_0_1(op_O_8_0_0_1),
    .O_8_0_0_2(op_O_8_0_0_2),
    .O_8_0_1_0(op_O_8_0_1_0),
    .O_8_0_1_1(op_O_8_0_1_1),
    .O_8_0_1_2(op_O_8_0_1_2),
    .O_9_0_0_0(op_O_9_0_0_0),
    .O_9_0_0_1(op_O_9_0_0_1),
    .O_9_0_0_2(op_O_9_0_0_2),
    .O_9_0_1_0(op_O_9_0_1_0),
    .O_9_0_1_1(op_O_9_0_1_1),
    .O_9_0_1_2(op_O_9_0_1_2),
    .O_10_0_0_0(op_O_10_0_0_0),
    .O_10_0_0_1(op_O_10_0_0_1),
    .O_10_0_0_2(op_O_10_0_0_2),
    .O_10_0_1_0(op_O_10_0_1_0),
    .O_10_0_1_1(op_O_10_0_1_1),
    .O_10_0_1_2(op_O_10_0_1_2),
    .O_11_0_0_0(op_O_11_0_0_0),
    .O_11_0_0_1(op_O_11_0_0_1),
    .O_11_0_0_2(op_O_11_0_0_2),
    .O_11_0_1_0(op_O_11_0_1_0),
    .O_11_0_1_1(op_O_11_0_1_1),
    .O_11_0_1_2(op_O_11_0_1_2),
    .O_12_0_0_0(op_O_12_0_0_0),
    .O_12_0_0_1(op_O_12_0_0_1),
    .O_12_0_0_2(op_O_12_0_0_2),
    .O_12_0_1_0(op_O_12_0_1_0),
    .O_12_0_1_1(op_O_12_0_1_1),
    .O_12_0_1_2(op_O_12_0_1_2),
    .O_13_0_0_0(op_O_13_0_0_0),
    .O_13_0_0_1(op_O_13_0_0_1),
    .O_13_0_0_2(op_O_13_0_0_2),
    .O_13_0_1_0(op_O_13_0_1_0),
    .O_13_0_1_1(op_O_13_0_1_1),
    .O_13_0_1_2(op_O_13_0_1_2),
    .O_14_0_0_0(op_O_14_0_0_0),
    .O_14_0_0_1(op_O_14_0_0_1),
    .O_14_0_0_2(op_O_14_0_0_2),
    .O_14_0_1_0(op_O_14_0_1_0),
    .O_14_0_1_1(op_O_14_0_1_1),
    .O_14_0_1_2(op_O_14_0_1_2),
    .O_15_0_0_0(op_O_15_0_0_0),
    .O_15_0_0_1(op_O_15_0_0_1),
    .O_15_0_0_2(op_O_15_0_0_2),
    .O_15_0_1_0(op_O_15_0_1_0),
    .O_15_0_1_1(op_O_15_0_1_1),
    .O_15_0_1_2(op_O_15_0_1_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_0_2 = op_O_0_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_0_1_0 = op_O_0_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_0_1_1 = op_O_0_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_0_1_2 = op_O_0_0_1_2; // @[Map2T.scala 17:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_0_2 = op_O_1_0_0_2; // @[Map2T.scala 17:7]
  assign O_1_0_1_0 = op_O_1_0_1_0; // @[Map2T.scala 17:7]
  assign O_1_0_1_1 = op_O_1_0_1_1; // @[Map2T.scala 17:7]
  assign O_1_0_1_2 = op_O_1_0_1_2; // @[Map2T.scala 17:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_0_2 = op_O_2_0_0_2; // @[Map2T.scala 17:7]
  assign O_2_0_1_0 = op_O_2_0_1_0; // @[Map2T.scala 17:7]
  assign O_2_0_1_1 = op_O_2_0_1_1; // @[Map2T.scala 17:7]
  assign O_2_0_1_2 = op_O_2_0_1_2; // @[Map2T.scala 17:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_0_2 = op_O_3_0_0_2; // @[Map2T.scala 17:7]
  assign O_3_0_1_0 = op_O_3_0_1_0; // @[Map2T.scala 17:7]
  assign O_3_0_1_1 = op_O_3_0_1_1; // @[Map2T.scala 17:7]
  assign O_3_0_1_2 = op_O_3_0_1_2; // @[Map2T.scala 17:7]
  assign O_4_0_0_0 = op_O_4_0_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_0_1 = op_O_4_0_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_0_2 = op_O_4_0_0_2; // @[Map2T.scala 17:7]
  assign O_4_0_1_0 = op_O_4_0_1_0; // @[Map2T.scala 17:7]
  assign O_4_0_1_1 = op_O_4_0_1_1; // @[Map2T.scala 17:7]
  assign O_4_0_1_2 = op_O_4_0_1_2; // @[Map2T.scala 17:7]
  assign O_5_0_0_0 = op_O_5_0_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_0_1 = op_O_5_0_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_0_2 = op_O_5_0_0_2; // @[Map2T.scala 17:7]
  assign O_5_0_1_0 = op_O_5_0_1_0; // @[Map2T.scala 17:7]
  assign O_5_0_1_1 = op_O_5_0_1_1; // @[Map2T.scala 17:7]
  assign O_5_0_1_2 = op_O_5_0_1_2; // @[Map2T.scala 17:7]
  assign O_6_0_0_0 = op_O_6_0_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_0_1 = op_O_6_0_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_0_2 = op_O_6_0_0_2; // @[Map2T.scala 17:7]
  assign O_6_0_1_0 = op_O_6_0_1_0; // @[Map2T.scala 17:7]
  assign O_6_0_1_1 = op_O_6_0_1_1; // @[Map2T.scala 17:7]
  assign O_6_0_1_2 = op_O_6_0_1_2; // @[Map2T.scala 17:7]
  assign O_7_0_0_0 = op_O_7_0_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_0_1 = op_O_7_0_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_0_2 = op_O_7_0_0_2; // @[Map2T.scala 17:7]
  assign O_7_0_1_0 = op_O_7_0_1_0; // @[Map2T.scala 17:7]
  assign O_7_0_1_1 = op_O_7_0_1_1; // @[Map2T.scala 17:7]
  assign O_7_0_1_2 = op_O_7_0_1_2; // @[Map2T.scala 17:7]
  assign O_8_0_0_0 = op_O_8_0_0_0; // @[Map2T.scala 17:7]
  assign O_8_0_0_1 = op_O_8_0_0_1; // @[Map2T.scala 17:7]
  assign O_8_0_0_2 = op_O_8_0_0_2; // @[Map2T.scala 17:7]
  assign O_8_0_1_0 = op_O_8_0_1_0; // @[Map2T.scala 17:7]
  assign O_8_0_1_1 = op_O_8_0_1_1; // @[Map2T.scala 17:7]
  assign O_8_0_1_2 = op_O_8_0_1_2; // @[Map2T.scala 17:7]
  assign O_9_0_0_0 = op_O_9_0_0_0; // @[Map2T.scala 17:7]
  assign O_9_0_0_1 = op_O_9_0_0_1; // @[Map2T.scala 17:7]
  assign O_9_0_0_2 = op_O_9_0_0_2; // @[Map2T.scala 17:7]
  assign O_9_0_1_0 = op_O_9_0_1_0; // @[Map2T.scala 17:7]
  assign O_9_0_1_1 = op_O_9_0_1_1; // @[Map2T.scala 17:7]
  assign O_9_0_1_2 = op_O_9_0_1_2; // @[Map2T.scala 17:7]
  assign O_10_0_0_0 = op_O_10_0_0_0; // @[Map2T.scala 17:7]
  assign O_10_0_0_1 = op_O_10_0_0_1; // @[Map2T.scala 17:7]
  assign O_10_0_0_2 = op_O_10_0_0_2; // @[Map2T.scala 17:7]
  assign O_10_0_1_0 = op_O_10_0_1_0; // @[Map2T.scala 17:7]
  assign O_10_0_1_1 = op_O_10_0_1_1; // @[Map2T.scala 17:7]
  assign O_10_0_1_2 = op_O_10_0_1_2; // @[Map2T.scala 17:7]
  assign O_11_0_0_0 = op_O_11_0_0_0; // @[Map2T.scala 17:7]
  assign O_11_0_0_1 = op_O_11_0_0_1; // @[Map2T.scala 17:7]
  assign O_11_0_0_2 = op_O_11_0_0_2; // @[Map2T.scala 17:7]
  assign O_11_0_1_0 = op_O_11_0_1_0; // @[Map2T.scala 17:7]
  assign O_11_0_1_1 = op_O_11_0_1_1; // @[Map2T.scala 17:7]
  assign O_11_0_1_2 = op_O_11_0_1_2; // @[Map2T.scala 17:7]
  assign O_12_0_0_0 = op_O_12_0_0_0; // @[Map2T.scala 17:7]
  assign O_12_0_0_1 = op_O_12_0_0_1; // @[Map2T.scala 17:7]
  assign O_12_0_0_2 = op_O_12_0_0_2; // @[Map2T.scala 17:7]
  assign O_12_0_1_0 = op_O_12_0_1_0; // @[Map2T.scala 17:7]
  assign O_12_0_1_1 = op_O_12_0_1_1; // @[Map2T.scala 17:7]
  assign O_12_0_1_2 = op_O_12_0_1_2; // @[Map2T.scala 17:7]
  assign O_13_0_0_0 = op_O_13_0_0_0; // @[Map2T.scala 17:7]
  assign O_13_0_0_1 = op_O_13_0_0_1; // @[Map2T.scala 17:7]
  assign O_13_0_0_2 = op_O_13_0_0_2; // @[Map2T.scala 17:7]
  assign O_13_0_1_0 = op_O_13_0_1_0; // @[Map2T.scala 17:7]
  assign O_13_0_1_1 = op_O_13_0_1_1; // @[Map2T.scala 17:7]
  assign O_13_0_1_2 = op_O_13_0_1_2; // @[Map2T.scala 17:7]
  assign O_14_0_0_0 = op_O_14_0_0_0; // @[Map2T.scala 17:7]
  assign O_14_0_0_1 = op_O_14_0_0_1; // @[Map2T.scala 17:7]
  assign O_14_0_0_2 = op_O_14_0_0_2; // @[Map2T.scala 17:7]
  assign O_14_0_1_0 = op_O_14_0_1_0; // @[Map2T.scala 17:7]
  assign O_14_0_1_1 = op_O_14_0_1_1; // @[Map2T.scala 17:7]
  assign O_14_0_1_2 = op_O_14_0_1_2; // @[Map2T.scala 17:7]
  assign O_15_0_0_0 = op_O_15_0_0_0; // @[Map2T.scala 17:7]
  assign O_15_0_0_1 = op_O_15_0_0_1; // @[Map2T.scala 17:7]
  assign O_15_0_0_2 = op_O_15_0_0_2; // @[Map2T.scala 17:7]
  assign O_15_0_1_0 = op_O_15_0_1_0; // @[Map2T.scala 17:7]
  assign O_15_0_1_1 = op_O_15_0_1_1; // @[Map2T.scala 17:7]
  assign O_15_0_1_2 = op_O_15_0_1_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0 = I0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1 = I0_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_0_2 = I0_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0 = I0_1_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1 = I0_1_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_2 = I0_1_0_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0 = I0_2_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1 = I0_2_0_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_2 = I0_2_0_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0 = I0_3_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1 = I0_3_0_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_2 = I0_3_0_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0 = I0_4_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_1 = I0_4_0_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0_2 = I0_4_0_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0 = I0_5_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_1 = I0_5_0_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0_2 = I0_5_0_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0 = I0_6_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_1 = I0_6_0_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0_2 = I0_6_0_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0 = I0_7_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_1 = I0_7_0_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0_2 = I0_7_0_2; // @[Map2T.scala 15:11]
  assign op_I0_8_0_0 = I0_8_0_0; // @[Map2T.scala 15:11]
  assign op_I0_8_0_1 = I0_8_0_1; // @[Map2T.scala 15:11]
  assign op_I0_8_0_2 = I0_8_0_2; // @[Map2T.scala 15:11]
  assign op_I0_9_0_0 = I0_9_0_0; // @[Map2T.scala 15:11]
  assign op_I0_9_0_1 = I0_9_0_1; // @[Map2T.scala 15:11]
  assign op_I0_9_0_2 = I0_9_0_2; // @[Map2T.scala 15:11]
  assign op_I0_10_0_0 = I0_10_0_0; // @[Map2T.scala 15:11]
  assign op_I0_10_0_1 = I0_10_0_1; // @[Map2T.scala 15:11]
  assign op_I0_10_0_2 = I0_10_0_2; // @[Map2T.scala 15:11]
  assign op_I0_11_0_0 = I0_11_0_0; // @[Map2T.scala 15:11]
  assign op_I0_11_0_1 = I0_11_0_1; // @[Map2T.scala 15:11]
  assign op_I0_11_0_2 = I0_11_0_2; // @[Map2T.scala 15:11]
  assign op_I0_12_0_0 = I0_12_0_0; // @[Map2T.scala 15:11]
  assign op_I0_12_0_1 = I0_12_0_1; // @[Map2T.scala 15:11]
  assign op_I0_12_0_2 = I0_12_0_2; // @[Map2T.scala 15:11]
  assign op_I0_13_0_0 = I0_13_0_0; // @[Map2T.scala 15:11]
  assign op_I0_13_0_1 = I0_13_0_1; // @[Map2T.scala 15:11]
  assign op_I0_13_0_2 = I0_13_0_2; // @[Map2T.scala 15:11]
  assign op_I0_14_0_0 = I0_14_0_0; // @[Map2T.scala 15:11]
  assign op_I0_14_0_1 = I0_14_0_1; // @[Map2T.scala 15:11]
  assign op_I0_14_0_2 = I0_14_0_2; // @[Map2T.scala 15:11]
  assign op_I0_15_0_0 = I0_15_0_0; // @[Map2T.scala 15:11]
  assign op_I0_15_0_1 = I0_15_0_1; // @[Map2T.scala 15:11]
  assign op_I0_15_0_2 = I0_15_0_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0_0 = I1_0_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_0_1 = I1_0_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_0_2 = I1_0_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0_0 = I1_1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_1_0_1 = I1_1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_1_0_2 = I1_1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0_0 = I1_2_0_0; // @[Map2T.scala 16:11]
  assign op_I1_2_0_1 = I1_2_0_1; // @[Map2T.scala 16:11]
  assign op_I1_2_0_2 = I1_2_0_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0_0 = I1_3_0_0; // @[Map2T.scala 16:11]
  assign op_I1_3_0_1 = I1_3_0_1; // @[Map2T.scala 16:11]
  assign op_I1_3_0_2 = I1_3_0_2; // @[Map2T.scala 16:11]
  assign op_I1_4_0_0 = I1_4_0_0; // @[Map2T.scala 16:11]
  assign op_I1_4_0_1 = I1_4_0_1; // @[Map2T.scala 16:11]
  assign op_I1_4_0_2 = I1_4_0_2; // @[Map2T.scala 16:11]
  assign op_I1_5_0_0 = I1_5_0_0; // @[Map2T.scala 16:11]
  assign op_I1_5_0_1 = I1_5_0_1; // @[Map2T.scala 16:11]
  assign op_I1_5_0_2 = I1_5_0_2; // @[Map2T.scala 16:11]
  assign op_I1_6_0_0 = I1_6_0_0; // @[Map2T.scala 16:11]
  assign op_I1_6_0_1 = I1_6_0_1; // @[Map2T.scala 16:11]
  assign op_I1_6_0_2 = I1_6_0_2; // @[Map2T.scala 16:11]
  assign op_I1_7_0_0 = I1_7_0_0; // @[Map2T.scala 16:11]
  assign op_I1_7_0_1 = I1_7_0_1; // @[Map2T.scala 16:11]
  assign op_I1_7_0_2 = I1_7_0_2; // @[Map2T.scala 16:11]
  assign op_I1_8_0_0 = I1_8_0_0; // @[Map2T.scala 16:11]
  assign op_I1_8_0_1 = I1_8_0_1; // @[Map2T.scala 16:11]
  assign op_I1_8_0_2 = I1_8_0_2; // @[Map2T.scala 16:11]
  assign op_I1_9_0_0 = I1_9_0_0; // @[Map2T.scala 16:11]
  assign op_I1_9_0_1 = I1_9_0_1; // @[Map2T.scala 16:11]
  assign op_I1_9_0_2 = I1_9_0_2; // @[Map2T.scala 16:11]
  assign op_I1_10_0_0 = I1_10_0_0; // @[Map2T.scala 16:11]
  assign op_I1_10_0_1 = I1_10_0_1; // @[Map2T.scala 16:11]
  assign op_I1_10_0_2 = I1_10_0_2; // @[Map2T.scala 16:11]
  assign op_I1_11_0_0 = I1_11_0_0; // @[Map2T.scala 16:11]
  assign op_I1_11_0_1 = I1_11_0_1; // @[Map2T.scala 16:11]
  assign op_I1_11_0_2 = I1_11_0_2; // @[Map2T.scala 16:11]
  assign op_I1_12_0_0 = I1_12_0_0; // @[Map2T.scala 16:11]
  assign op_I1_12_0_1 = I1_12_0_1; // @[Map2T.scala 16:11]
  assign op_I1_12_0_2 = I1_12_0_2; // @[Map2T.scala 16:11]
  assign op_I1_13_0_0 = I1_13_0_0; // @[Map2T.scala 16:11]
  assign op_I1_13_0_1 = I1_13_0_1; // @[Map2T.scala 16:11]
  assign op_I1_13_0_2 = I1_13_0_2; // @[Map2T.scala 16:11]
  assign op_I1_14_0_0 = I1_14_0_0; // @[Map2T.scala 16:11]
  assign op_I1_14_0_1 = I1_14_0_1; // @[Map2T.scala 16:11]
  assign op_I1_14_0_2 = I1_14_0_2; // @[Map2T.scala 16:11]
  assign op_I1_15_0_0 = I1_15_0_0; // @[Map2T.scala 16:11]
  assign op_I1_15_0_1 = I1_15_0_1; // @[Map2T.scala 16:11]
  assign op_I1_15_0_2 = I1_15_0_2; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_1_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0_0 = I0_0_0; // @[Tuple.scala 24:34]
  assign O_0_1 = I0_0_1; // @[Tuple.scala 24:34]
  assign O_0_2 = I0_0_2; // @[Tuple.scala 24:34]
  assign O_1_0 = I0_1_0; // @[Tuple.scala 24:34]
  assign O_1_1 = I0_1_1; // @[Tuple.scala 24:34]
  assign O_1_2 = I0_1_2; // @[Tuple.scala 24:34]
  assign O_2_0 = I1_0; // @[Tuple.scala 26:32]
  assign O_2_1 = I1_1; // @[Tuple.scala 26:32]
  assign O_2_2 = I1_2; // @[Tuple.scala 26:32]
endmodule
module Map2S_20(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_0_0_1,
  input  [7:0] I0_0_0_2,
  input  [7:0] I0_0_1_0,
  input  [7:0] I0_0_1_1,
  input  [7:0] I0_0_1_2,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_0_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_2; // @[Map2S.scala 9:22]
  SSeqTupleAppender_3 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I0_1_0(fst_op_I0_1_0),
    .I0_1_1(fst_op_I0_1_1),
    .I0_1_2(fst_op_I0_1_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[Map2S.scala 19:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[Map2S.scala 19:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_0 = I0_0_1_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_1 = I0_0_1_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_2 = I0_0_1_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
endmodule
module Map2S_21(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0_0,
  input  [7:0] I0_0_0_0_1,
  input  [7:0] I0_0_0_0_2,
  input  [7:0] I0_0_0_1_0,
  input  [7:0] I0_0_0_1_1,
  input  [7:0] I0_0_0_1_2,
  input  [7:0] I0_1_0_0_0,
  input  [7:0] I0_1_0_0_1,
  input  [7:0] I0_1_0_0_2,
  input  [7:0] I0_1_0_1_0,
  input  [7:0] I0_1_0_1_1,
  input  [7:0] I0_1_0_1_2,
  input  [7:0] I0_2_0_0_0,
  input  [7:0] I0_2_0_0_1,
  input  [7:0] I0_2_0_0_2,
  input  [7:0] I0_2_0_1_0,
  input  [7:0] I0_2_0_1_1,
  input  [7:0] I0_2_0_1_2,
  input  [7:0] I0_3_0_0_0,
  input  [7:0] I0_3_0_0_1,
  input  [7:0] I0_3_0_0_2,
  input  [7:0] I0_3_0_1_0,
  input  [7:0] I0_3_0_1_1,
  input  [7:0] I0_3_0_1_2,
  input  [7:0] I0_4_0_0_0,
  input  [7:0] I0_4_0_0_1,
  input  [7:0] I0_4_0_0_2,
  input  [7:0] I0_4_0_1_0,
  input  [7:0] I0_4_0_1_1,
  input  [7:0] I0_4_0_1_2,
  input  [7:0] I0_5_0_0_0,
  input  [7:0] I0_5_0_0_1,
  input  [7:0] I0_5_0_0_2,
  input  [7:0] I0_5_0_1_0,
  input  [7:0] I0_5_0_1_1,
  input  [7:0] I0_5_0_1_2,
  input  [7:0] I0_6_0_0_0,
  input  [7:0] I0_6_0_0_1,
  input  [7:0] I0_6_0_0_2,
  input  [7:0] I0_6_0_1_0,
  input  [7:0] I0_6_0_1_1,
  input  [7:0] I0_6_0_1_2,
  input  [7:0] I0_7_0_0_0,
  input  [7:0] I0_7_0_0_1,
  input  [7:0] I0_7_0_0_2,
  input  [7:0] I0_7_0_1_0,
  input  [7:0] I0_7_0_1_1,
  input  [7:0] I0_7_0_1_2,
  input  [7:0] I0_8_0_0_0,
  input  [7:0] I0_8_0_0_1,
  input  [7:0] I0_8_0_0_2,
  input  [7:0] I0_8_0_1_0,
  input  [7:0] I0_8_0_1_1,
  input  [7:0] I0_8_0_1_2,
  input  [7:0] I0_9_0_0_0,
  input  [7:0] I0_9_0_0_1,
  input  [7:0] I0_9_0_0_2,
  input  [7:0] I0_9_0_1_0,
  input  [7:0] I0_9_0_1_1,
  input  [7:0] I0_9_0_1_2,
  input  [7:0] I0_10_0_0_0,
  input  [7:0] I0_10_0_0_1,
  input  [7:0] I0_10_0_0_2,
  input  [7:0] I0_10_0_1_0,
  input  [7:0] I0_10_0_1_1,
  input  [7:0] I0_10_0_1_2,
  input  [7:0] I0_11_0_0_0,
  input  [7:0] I0_11_0_0_1,
  input  [7:0] I0_11_0_0_2,
  input  [7:0] I0_11_0_1_0,
  input  [7:0] I0_11_0_1_1,
  input  [7:0] I0_11_0_1_2,
  input  [7:0] I0_12_0_0_0,
  input  [7:0] I0_12_0_0_1,
  input  [7:0] I0_12_0_0_2,
  input  [7:0] I0_12_0_1_0,
  input  [7:0] I0_12_0_1_1,
  input  [7:0] I0_12_0_1_2,
  input  [7:0] I0_13_0_0_0,
  input  [7:0] I0_13_0_0_1,
  input  [7:0] I0_13_0_0_2,
  input  [7:0] I0_13_0_1_0,
  input  [7:0] I0_13_0_1_1,
  input  [7:0] I0_13_0_1_2,
  input  [7:0] I0_14_0_0_0,
  input  [7:0] I0_14_0_0_1,
  input  [7:0] I0_14_0_0_2,
  input  [7:0] I0_14_0_1_0,
  input  [7:0] I0_14_0_1_1,
  input  [7:0] I0_14_0_1_2,
  input  [7:0] I0_15_0_0_0,
  input  [7:0] I0_15_0_0_1,
  input  [7:0] I0_15_0_0_2,
  input  [7:0] I0_15_0_1_0,
  input  [7:0] I0_15_0_1_1,
  input  [7:0] I0_15_0_1_2,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_0_0_1,
  input  [7:0] I1_0_0_2,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_1_0_1,
  input  [7:0] I1_1_0_2,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_2_0_1,
  input  [7:0] I1_2_0_2,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_3_0_1,
  input  [7:0] I1_3_0_2,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_4_0_1,
  input  [7:0] I1_4_0_2,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_5_0_1,
  input  [7:0] I1_5_0_2,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_6_0_1,
  input  [7:0] I1_6_0_2,
  input  [7:0] I1_7_0_0,
  input  [7:0] I1_7_0_1,
  input  [7:0] I1_7_0_2,
  input  [7:0] I1_8_0_0,
  input  [7:0] I1_8_0_1,
  input  [7:0] I1_8_0_2,
  input  [7:0] I1_9_0_0,
  input  [7:0] I1_9_0_1,
  input  [7:0] I1_9_0_2,
  input  [7:0] I1_10_0_0,
  input  [7:0] I1_10_0_1,
  input  [7:0] I1_10_0_2,
  input  [7:0] I1_11_0_0,
  input  [7:0] I1_11_0_1,
  input  [7:0] I1_11_0_2,
  input  [7:0] I1_12_0_0,
  input  [7:0] I1_12_0_1,
  input  [7:0] I1_12_0_2,
  input  [7:0] I1_13_0_0,
  input  [7:0] I1_13_0_1,
  input  [7:0] I1_13_0_2,
  input  [7:0] I1_14_0_0,
  input  [7:0] I1_14_0_1,
  input  [7:0] I1_14_0_2,
  input  [7:0] I1_15_0_0,
  input  [7:0] I1_15_0_1,
  input  [7:0] I1_15_0_2,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_0_0_1_0,
  output [7:0] O_0_0_1_1,
  output [7:0] O_0_0_1_2,
  output [7:0] O_0_0_2_0,
  output [7:0] O_0_0_2_1,
  output [7:0] O_0_0_2_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_1_0_1_0,
  output [7:0] O_1_0_1_1,
  output [7:0] O_1_0_1_2,
  output [7:0] O_1_0_2_0,
  output [7:0] O_1_0_2_1,
  output [7:0] O_1_0_2_2,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_0_2,
  output [7:0] O_2_0_1_0,
  output [7:0] O_2_0_1_1,
  output [7:0] O_2_0_1_2,
  output [7:0] O_2_0_2_0,
  output [7:0] O_2_0_2_1,
  output [7:0] O_2_0_2_2,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_0_2,
  output [7:0] O_3_0_1_0,
  output [7:0] O_3_0_1_1,
  output [7:0] O_3_0_1_2,
  output [7:0] O_3_0_2_0,
  output [7:0] O_3_0_2_1,
  output [7:0] O_3_0_2_2,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_0_2,
  output [7:0] O_4_0_1_0,
  output [7:0] O_4_0_1_1,
  output [7:0] O_4_0_1_2,
  output [7:0] O_4_0_2_0,
  output [7:0] O_4_0_2_1,
  output [7:0] O_4_0_2_2,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_0_2,
  output [7:0] O_5_0_1_0,
  output [7:0] O_5_0_1_1,
  output [7:0] O_5_0_1_2,
  output [7:0] O_5_0_2_0,
  output [7:0] O_5_0_2_1,
  output [7:0] O_5_0_2_2,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_0_2,
  output [7:0] O_6_0_1_0,
  output [7:0] O_6_0_1_1,
  output [7:0] O_6_0_1_2,
  output [7:0] O_6_0_2_0,
  output [7:0] O_6_0_2_1,
  output [7:0] O_6_0_2_2,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_0_2,
  output [7:0] O_7_0_1_0,
  output [7:0] O_7_0_1_1,
  output [7:0] O_7_0_1_2,
  output [7:0] O_7_0_2_0,
  output [7:0] O_7_0_2_1,
  output [7:0] O_7_0_2_2,
  output [7:0] O_8_0_0_0,
  output [7:0] O_8_0_0_1,
  output [7:0] O_8_0_0_2,
  output [7:0] O_8_0_1_0,
  output [7:0] O_8_0_1_1,
  output [7:0] O_8_0_1_2,
  output [7:0] O_8_0_2_0,
  output [7:0] O_8_0_2_1,
  output [7:0] O_8_0_2_2,
  output [7:0] O_9_0_0_0,
  output [7:0] O_9_0_0_1,
  output [7:0] O_9_0_0_2,
  output [7:0] O_9_0_1_0,
  output [7:0] O_9_0_1_1,
  output [7:0] O_9_0_1_2,
  output [7:0] O_9_0_2_0,
  output [7:0] O_9_0_2_1,
  output [7:0] O_9_0_2_2,
  output [7:0] O_10_0_0_0,
  output [7:0] O_10_0_0_1,
  output [7:0] O_10_0_0_2,
  output [7:0] O_10_0_1_0,
  output [7:0] O_10_0_1_1,
  output [7:0] O_10_0_1_2,
  output [7:0] O_10_0_2_0,
  output [7:0] O_10_0_2_1,
  output [7:0] O_10_0_2_2,
  output [7:0] O_11_0_0_0,
  output [7:0] O_11_0_0_1,
  output [7:0] O_11_0_0_2,
  output [7:0] O_11_0_1_0,
  output [7:0] O_11_0_1_1,
  output [7:0] O_11_0_1_2,
  output [7:0] O_11_0_2_0,
  output [7:0] O_11_0_2_1,
  output [7:0] O_11_0_2_2,
  output [7:0] O_12_0_0_0,
  output [7:0] O_12_0_0_1,
  output [7:0] O_12_0_0_2,
  output [7:0] O_12_0_1_0,
  output [7:0] O_12_0_1_1,
  output [7:0] O_12_0_1_2,
  output [7:0] O_12_0_2_0,
  output [7:0] O_12_0_2_1,
  output [7:0] O_12_0_2_2,
  output [7:0] O_13_0_0_0,
  output [7:0] O_13_0_0_1,
  output [7:0] O_13_0_0_2,
  output [7:0] O_13_0_1_0,
  output [7:0] O_13_0_1_1,
  output [7:0] O_13_0_1_2,
  output [7:0] O_13_0_2_0,
  output [7:0] O_13_0_2_1,
  output [7:0] O_13_0_2_2,
  output [7:0] O_14_0_0_0,
  output [7:0] O_14_0_0_1,
  output [7:0] O_14_0_0_2,
  output [7:0] O_14_0_1_0,
  output [7:0] O_14_0_1_1,
  output [7:0] O_14_0_1_2,
  output [7:0] O_14_0_2_0,
  output [7:0] O_14_0_2_1,
  output [7:0] O_14_0_2_2,
  output [7:0] O_15_0_0_0,
  output [7:0] O_15_0_0_1,
  output [7:0] O_15_0_0_2,
  output [7:0] O_15_0_1_0,
  output [7:0] O_15_0_1_1,
  output [7:0] O_15_0_1_2,
  output [7:0] O_15_0_2_0,
  output [7:0] O_15_0_2_1,
  output [7:0] O_15_0_2_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_2_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  Map2S_20 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0_0(fst_op_I0_0_0_0),
    .I0_0_0_1(fst_op_I0_0_0_1),
    .I0_0_0_2(fst_op_I0_0_0_2),
    .I0_0_1_0(fst_op_I0_0_1_0),
    .I0_0_1_1(fst_op_I0_0_1_1),
    .I0_0_1_2(fst_op_I0_0_1_2),
    .I1_0_0(fst_op_I1_0_0),
    .I1_0_1(fst_op_I1_0_1),
    .I1_0_2(fst_op_I1_0_2),
    .O_0_0_0(fst_op_O_0_0_0),
    .O_0_0_1(fst_op_O_0_0_1),
    .O_0_0_2(fst_op_O_0_0_2),
    .O_0_1_0(fst_op_O_0_1_0),
    .O_0_1_1(fst_op_O_0_1_1),
    .O_0_1_2(fst_op_O_0_1_2),
    .O_0_2_0(fst_op_O_0_2_0),
    .O_0_2_1(fst_op_O_0_2_1),
    .O_0_2_2(fst_op_O_0_2_2)
  );
  Map2S_20 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0_0(other_ops_0_I0_0_0_0),
    .I0_0_0_1(other_ops_0_I0_0_0_1),
    .I0_0_0_2(other_ops_0_I0_0_0_2),
    .I0_0_1_0(other_ops_0_I0_0_1_0),
    .I0_0_1_1(other_ops_0_I0_0_1_1),
    .I0_0_1_2(other_ops_0_I0_0_1_2),
    .I1_0_0(other_ops_0_I1_0_0),
    .I1_0_1(other_ops_0_I1_0_1),
    .I1_0_2(other_ops_0_I1_0_2),
    .O_0_0_0(other_ops_0_O_0_0_0),
    .O_0_0_1(other_ops_0_O_0_0_1),
    .O_0_0_2(other_ops_0_O_0_0_2),
    .O_0_1_0(other_ops_0_O_0_1_0),
    .O_0_1_1(other_ops_0_O_0_1_1),
    .O_0_1_2(other_ops_0_O_0_1_2),
    .O_0_2_0(other_ops_0_O_0_2_0),
    .O_0_2_1(other_ops_0_O_0_2_1),
    .O_0_2_2(other_ops_0_O_0_2_2)
  );
  Map2S_20 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0_0(other_ops_1_I0_0_0_0),
    .I0_0_0_1(other_ops_1_I0_0_0_1),
    .I0_0_0_2(other_ops_1_I0_0_0_2),
    .I0_0_1_0(other_ops_1_I0_0_1_0),
    .I0_0_1_1(other_ops_1_I0_0_1_1),
    .I0_0_1_2(other_ops_1_I0_0_1_2),
    .I1_0_0(other_ops_1_I1_0_0),
    .I1_0_1(other_ops_1_I1_0_1),
    .I1_0_2(other_ops_1_I1_0_2),
    .O_0_0_0(other_ops_1_O_0_0_0),
    .O_0_0_1(other_ops_1_O_0_0_1),
    .O_0_0_2(other_ops_1_O_0_0_2),
    .O_0_1_0(other_ops_1_O_0_1_0),
    .O_0_1_1(other_ops_1_O_0_1_1),
    .O_0_1_2(other_ops_1_O_0_1_2),
    .O_0_2_0(other_ops_1_O_0_2_0),
    .O_0_2_1(other_ops_1_O_0_2_1),
    .O_0_2_2(other_ops_1_O_0_2_2)
  );
  Map2S_20 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0_0(other_ops_2_I0_0_0_0),
    .I0_0_0_1(other_ops_2_I0_0_0_1),
    .I0_0_0_2(other_ops_2_I0_0_0_2),
    .I0_0_1_0(other_ops_2_I0_0_1_0),
    .I0_0_1_1(other_ops_2_I0_0_1_1),
    .I0_0_1_2(other_ops_2_I0_0_1_2),
    .I1_0_0(other_ops_2_I1_0_0),
    .I1_0_1(other_ops_2_I1_0_1),
    .I1_0_2(other_ops_2_I1_0_2),
    .O_0_0_0(other_ops_2_O_0_0_0),
    .O_0_0_1(other_ops_2_O_0_0_1),
    .O_0_0_2(other_ops_2_O_0_0_2),
    .O_0_1_0(other_ops_2_O_0_1_0),
    .O_0_1_1(other_ops_2_O_0_1_1),
    .O_0_1_2(other_ops_2_O_0_1_2),
    .O_0_2_0(other_ops_2_O_0_2_0),
    .O_0_2_1(other_ops_2_O_0_2_1),
    .O_0_2_2(other_ops_2_O_0_2_2)
  );
  Map2S_20 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0_0(other_ops_3_I0_0_0_0),
    .I0_0_0_1(other_ops_3_I0_0_0_1),
    .I0_0_0_2(other_ops_3_I0_0_0_2),
    .I0_0_1_0(other_ops_3_I0_0_1_0),
    .I0_0_1_1(other_ops_3_I0_0_1_1),
    .I0_0_1_2(other_ops_3_I0_0_1_2),
    .I1_0_0(other_ops_3_I1_0_0),
    .I1_0_1(other_ops_3_I1_0_1),
    .I1_0_2(other_ops_3_I1_0_2),
    .O_0_0_0(other_ops_3_O_0_0_0),
    .O_0_0_1(other_ops_3_O_0_0_1),
    .O_0_0_2(other_ops_3_O_0_0_2),
    .O_0_1_0(other_ops_3_O_0_1_0),
    .O_0_1_1(other_ops_3_O_0_1_1),
    .O_0_1_2(other_ops_3_O_0_1_2),
    .O_0_2_0(other_ops_3_O_0_2_0),
    .O_0_2_1(other_ops_3_O_0_2_1),
    .O_0_2_2(other_ops_3_O_0_2_2)
  );
  Map2S_20 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0_0(other_ops_4_I0_0_0_0),
    .I0_0_0_1(other_ops_4_I0_0_0_1),
    .I0_0_0_2(other_ops_4_I0_0_0_2),
    .I0_0_1_0(other_ops_4_I0_0_1_0),
    .I0_0_1_1(other_ops_4_I0_0_1_1),
    .I0_0_1_2(other_ops_4_I0_0_1_2),
    .I1_0_0(other_ops_4_I1_0_0),
    .I1_0_1(other_ops_4_I1_0_1),
    .I1_0_2(other_ops_4_I1_0_2),
    .O_0_0_0(other_ops_4_O_0_0_0),
    .O_0_0_1(other_ops_4_O_0_0_1),
    .O_0_0_2(other_ops_4_O_0_0_2),
    .O_0_1_0(other_ops_4_O_0_1_0),
    .O_0_1_1(other_ops_4_O_0_1_1),
    .O_0_1_2(other_ops_4_O_0_1_2),
    .O_0_2_0(other_ops_4_O_0_2_0),
    .O_0_2_1(other_ops_4_O_0_2_1),
    .O_0_2_2(other_ops_4_O_0_2_2)
  );
  Map2S_20 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0_0(other_ops_5_I0_0_0_0),
    .I0_0_0_1(other_ops_5_I0_0_0_1),
    .I0_0_0_2(other_ops_5_I0_0_0_2),
    .I0_0_1_0(other_ops_5_I0_0_1_0),
    .I0_0_1_1(other_ops_5_I0_0_1_1),
    .I0_0_1_2(other_ops_5_I0_0_1_2),
    .I1_0_0(other_ops_5_I1_0_0),
    .I1_0_1(other_ops_5_I1_0_1),
    .I1_0_2(other_ops_5_I1_0_2),
    .O_0_0_0(other_ops_5_O_0_0_0),
    .O_0_0_1(other_ops_5_O_0_0_1),
    .O_0_0_2(other_ops_5_O_0_0_2),
    .O_0_1_0(other_ops_5_O_0_1_0),
    .O_0_1_1(other_ops_5_O_0_1_1),
    .O_0_1_2(other_ops_5_O_0_1_2),
    .O_0_2_0(other_ops_5_O_0_2_0),
    .O_0_2_1(other_ops_5_O_0_2_1),
    .O_0_2_2(other_ops_5_O_0_2_2)
  );
  Map2S_20 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0_0(other_ops_6_I0_0_0_0),
    .I0_0_0_1(other_ops_6_I0_0_0_1),
    .I0_0_0_2(other_ops_6_I0_0_0_2),
    .I0_0_1_0(other_ops_6_I0_0_1_0),
    .I0_0_1_1(other_ops_6_I0_0_1_1),
    .I0_0_1_2(other_ops_6_I0_0_1_2),
    .I1_0_0(other_ops_6_I1_0_0),
    .I1_0_1(other_ops_6_I1_0_1),
    .I1_0_2(other_ops_6_I1_0_2),
    .O_0_0_0(other_ops_6_O_0_0_0),
    .O_0_0_1(other_ops_6_O_0_0_1),
    .O_0_0_2(other_ops_6_O_0_0_2),
    .O_0_1_0(other_ops_6_O_0_1_0),
    .O_0_1_1(other_ops_6_O_0_1_1),
    .O_0_1_2(other_ops_6_O_0_1_2),
    .O_0_2_0(other_ops_6_O_0_2_0),
    .O_0_2_1(other_ops_6_O_0_2_1),
    .O_0_2_2(other_ops_6_O_0_2_2)
  );
  Map2S_20 other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0_0_0(other_ops_7_I0_0_0_0),
    .I0_0_0_1(other_ops_7_I0_0_0_1),
    .I0_0_0_2(other_ops_7_I0_0_0_2),
    .I0_0_1_0(other_ops_7_I0_0_1_0),
    .I0_0_1_1(other_ops_7_I0_0_1_1),
    .I0_0_1_2(other_ops_7_I0_0_1_2),
    .I1_0_0(other_ops_7_I1_0_0),
    .I1_0_1(other_ops_7_I1_0_1),
    .I1_0_2(other_ops_7_I1_0_2),
    .O_0_0_0(other_ops_7_O_0_0_0),
    .O_0_0_1(other_ops_7_O_0_0_1),
    .O_0_0_2(other_ops_7_O_0_0_2),
    .O_0_1_0(other_ops_7_O_0_1_0),
    .O_0_1_1(other_ops_7_O_0_1_1),
    .O_0_1_2(other_ops_7_O_0_1_2),
    .O_0_2_0(other_ops_7_O_0_2_0),
    .O_0_2_1(other_ops_7_O_0_2_1),
    .O_0_2_2(other_ops_7_O_0_2_2)
  );
  Map2S_20 other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0_0_0(other_ops_8_I0_0_0_0),
    .I0_0_0_1(other_ops_8_I0_0_0_1),
    .I0_0_0_2(other_ops_8_I0_0_0_2),
    .I0_0_1_0(other_ops_8_I0_0_1_0),
    .I0_0_1_1(other_ops_8_I0_0_1_1),
    .I0_0_1_2(other_ops_8_I0_0_1_2),
    .I1_0_0(other_ops_8_I1_0_0),
    .I1_0_1(other_ops_8_I1_0_1),
    .I1_0_2(other_ops_8_I1_0_2),
    .O_0_0_0(other_ops_8_O_0_0_0),
    .O_0_0_1(other_ops_8_O_0_0_1),
    .O_0_0_2(other_ops_8_O_0_0_2),
    .O_0_1_0(other_ops_8_O_0_1_0),
    .O_0_1_1(other_ops_8_O_0_1_1),
    .O_0_1_2(other_ops_8_O_0_1_2),
    .O_0_2_0(other_ops_8_O_0_2_0),
    .O_0_2_1(other_ops_8_O_0_2_1),
    .O_0_2_2(other_ops_8_O_0_2_2)
  );
  Map2S_20 other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0_0_0(other_ops_9_I0_0_0_0),
    .I0_0_0_1(other_ops_9_I0_0_0_1),
    .I0_0_0_2(other_ops_9_I0_0_0_2),
    .I0_0_1_0(other_ops_9_I0_0_1_0),
    .I0_0_1_1(other_ops_9_I0_0_1_1),
    .I0_0_1_2(other_ops_9_I0_0_1_2),
    .I1_0_0(other_ops_9_I1_0_0),
    .I1_0_1(other_ops_9_I1_0_1),
    .I1_0_2(other_ops_9_I1_0_2),
    .O_0_0_0(other_ops_9_O_0_0_0),
    .O_0_0_1(other_ops_9_O_0_0_1),
    .O_0_0_2(other_ops_9_O_0_0_2),
    .O_0_1_0(other_ops_9_O_0_1_0),
    .O_0_1_1(other_ops_9_O_0_1_1),
    .O_0_1_2(other_ops_9_O_0_1_2),
    .O_0_2_0(other_ops_9_O_0_2_0),
    .O_0_2_1(other_ops_9_O_0_2_1),
    .O_0_2_2(other_ops_9_O_0_2_2)
  );
  Map2S_20 other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0_0_0(other_ops_10_I0_0_0_0),
    .I0_0_0_1(other_ops_10_I0_0_0_1),
    .I0_0_0_2(other_ops_10_I0_0_0_2),
    .I0_0_1_0(other_ops_10_I0_0_1_0),
    .I0_0_1_1(other_ops_10_I0_0_1_1),
    .I0_0_1_2(other_ops_10_I0_0_1_2),
    .I1_0_0(other_ops_10_I1_0_0),
    .I1_0_1(other_ops_10_I1_0_1),
    .I1_0_2(other_ops_10_I1_0_2),
    .O_0_0_0(other_ops_10_O_0_0_0),
    .O_0_0_1(other_ops_10_O_0_0_1),
    .O_0_0_2(other_ops_10_O_0_0_2),
    .O_0_1_0(other_ops_10_O_0_1_0),
    .O_0_1_1(other_ops_10_O_0_1_1),
    .O_0_1_2(other_ops_10_O_0_1_2),
    .O_0_2_0(other_ops_10_O_0_2_0),
    .O_0_2_1(other_ops_10_O_0_2_1),
    .O_0_2_2(other_ops_10_O_0_2_2)
  );
  Map2S_20 other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0_0_0(other_ops_11_I0_0_0_0),
    .I0_0_0_1(other_ops_11_I0_0_0_1),
    .I0_0_0_2(other_ops_11_I0_0_0_2),
    .I0_0_1_0(other_ops_11_I0_0_1_0),
    .I0_0_1_1(other_ops_11_I0_0_1_1),
    .I0_0_1_2(other_ops_11_I0_0_1_2),
    .I1_0_0(other_ops_11_I1_0_0),
    .I1_0_1(other_ops_11_I1_0_1),
    .I1_0_2(other_ops_11_I1_0_2),
    .O_0_0_0(other_ops_11_O_0_0_0),
    .O_0_0_1(other_ops_11_O_0_0_1),
    .O_0_0_2(other_ops_11_O_0_0_2),
    .O_0_1_0(other_ops_11_O_0_1_0),
    .O_0_1_1(other_ops_11_O_0_1_1),
    .O_0_1_2(other_ops_11_O_0_1_2),
    .O_0_2_0(other_ops_11_O_0_2_0),
    .O_0_2_1(other_ops_11_O_0_2_1),
    .O_0_2_2(other_ops_11_O_0_2_2)
  );
  Map2S_20 other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0_0_0(other_ops_12_I0_0_0_0),
    .I0_0_0_1(other_ops_12_I0_0_0_1),
    .I0_0_0_2(other_ops_12_I0_0_0_2),
    .I0_0_1_0(other_ops_12_I0_0_1_0),
    .I0_0_1_1(other_ops_12_I0_0_1_1),
    .I0_0_1_2(other_ops_12_I0_0_1_2),
    .I1_0_0(other_ops_12_I1_0_0),
    .I1_0_1(other_ops_12_I1_0_1),
    .I1_0_2(other_ops_12_I1_0_2),
    .O_0_0_0(other_ops_12_O_0_0_0),
    .O_0_0_1(other_ops_12_O_0_0_1),
    .O_0_0_2(other_ops_12_O_0_0_2),
    .O_0_1_0(other_ops_12_O_0_1_0),
    .O_0_1_1(other_ops_12_O_0_1_1),
    .O_0_1_2(other_ops_12_O_0_1_2),
    .O_0_2_0(other_ops_12_O_0_2_0),
    .O_0_2_1(other_ops_12_O_0_2_1),
    .O_0_2_2(other_ops_12_O_0_2_2)
  );
  Map2S_20 other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0_0_0(other_ops_13_I0_0_0_0),
    .I0_0_0_1(other_ops_13_I0_0_0_1),
    .I0_0_0_2(other_ops_13_I0_0_0_2),
    .I0_0_1_0(other_ops_13_I0_0_1_0),
    .I0_0_1_1(other_ops_13_I0_0_1_1),
    .I0_0_1_2(other_ops_13_I0_0_1_2),
    .I1_0_0(other_ops_13_I1_0_0),
    .I1_0_1(other_ops_13_I1_0_1),
    .I1_0_2(other_ops_13_I1_0_2),
    .O_0_0_0(other_ops_13_O_0_0_0),
    .O_0_0_1(other_ops_13_O_0_0_1),
    .O_0_0_2(other_ops_13_O_0_0_2),
    .O_0_1_0(other_ops_13_O_0_1_0),
    .O_0_1_1(other_ops_13_O_0_1_1),
    .O_0_1_2(other_ops_13_O_0_1_2),
    .O_0_2_0(other_ops_13_O_0_2_0),
    .O_0_2_1(other_ops_13_O_0_2_1),
    .O_0_2_2(other_ops_13_O_0_2_2)
  );
  Map2S_20 other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0_0_0(other_ops_14_I0_0_0_0),
    .I0_0_0_1(other_ops_14_I0_0_0_1),
    .I0_0_0_2(other_ops_14_I0_0_0_2),
    .I0_0_1_0(other_ops_14_I0_0_1_0),
    .I0_0_1_1(other_ops_14_I0_0_1_1),
    .I0_0_1_2(other_ops_14_I0_0_1_2),
    .I1_0_0(other_ops_14_I1_0_0),
    .I1_0_1(other_ops_14_I1_0_1),
    .I1_0_2(other_ops_14_I1_0_2),
    .O_0_0_0(other_ops_14_O_0_0_0),
    .O_0_0_1(other_ops_14_O_0_0_1),
    .O_0_0_2(other_ops_14_O_0_0_2),
    .O_0_1_0(other_ops_14_O_0_1_0),
    .O_0_1_1(other_ops_14_O_0_1_1),
    .O_0_1_2(other_ops_14_O_0_1_2),
    .O_0_2_0(other_ops_14_O_0_2_0),
    .O_0_2_1(other_ops_14_O_0_2_1),
    .O_0_2_2(other_ops_14_O_0_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0_0 = fst_op_O_0_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_0_1 = fst_op_O_0_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_0_2 = fst_op_O_0_0_2; // @[Map2S.scala 19:8]
  assign O_0_0_1_0 = fst_op_O_0_1_0; // @[Map2S.scala 19:8]
  assign O_0_0_1_1 = fst_op_O_0_1_1; // @[Map2S.scala 19:8]
  assign O_0_0_1_2 = fst_op_O_0_1_2; // @[Map2S.scala 19:8]
  assign O_0_0_2_0 = fst_op_O_0_2_0; // @[Map2S.scala 19:8]
  assign O_0_0_2_1 = fst_op_O_0_2_1; // @[Map2S.scala 19:8]
  assign O_0_0_2_2 = fst_op_O_0_2_2; // @[Map2S.scala 19:8]
  assign O_1_0_0_0 = other_ops_0_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_0_1 = other_ops_0_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_0_2 = other_ops_0_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_1_0_1_0 = other_ops_0_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_1_0_1_1 = other_ops_0_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_1_0_1_2 = other_ops_0_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_1_0_2_0 = other_ops_0_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_1_0_2_1 = other_ops_0_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_1_0_2_2 = other_ops_0_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_2_0_0_0 = other_ops_1_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_0_1 = other_ops_1_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_0_2 = other_ops_1_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_2_0_1_0 = other_ops_1_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_2_0_1_1 = other_ops_1_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_2_0_1_2 = other_ops_1_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_2_0_2_0 = other_ops_1_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_2_0_2_1 = other_ops_1_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_2_0_2_2 = other_ops_1_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_3_0_0_0 = other_ops_2_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_0_1 = other_ops_2_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_0_2 = other_ops_2_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_3_0_1_0 = other_ops_2_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_3_0_1_1 = other_ops_2_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_3_0_1_2 = other_ops_2_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_3_0_2_0 = other_ops_2_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_3_0_2_1 = other_ops_2_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_3_0_2_2 = other_ops_2_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_4_0_0_0 = other_ops_3_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_0_1 = other_ops_3_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_0_2 = other_ops_3_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_4_0_1_0 = other_ops_3_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_4_0_1_1 = other_ops_3_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_4_0_1_2 = other_ops_3_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_4_0_2_0 = other_ops_3_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_4_0_2_1 = other_ops_3_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_4_0_2_2 = other_ops_3_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_5_0_0_0 = other_ops_4_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_0_1 = other_ops_4_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_0_2 = other_ops_4_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_5_0_1_0 = other_ops_4_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_5_0_1_1 = other_ops_4_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_5_0_1_2 = other_ops_4_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_5_0_2_0 = other_ops_4_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_5_0_2_1 = other_ops_4_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_5_0_2_2 = other_ops_4_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_6_0_0_0 = other_ops_5_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_0_1 = other_ops_5_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_0_2 = other_ops_5_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_6_0_1_0 = other_ops_5_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_6_0_1_1 = other_ops_5_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_6_0_1_2 = other_ops_5_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_6_0_2_0 = other_ops_5_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_6_0_2_1 = other_ops_5_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_6_0_2_2 = other_ops_5_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_7_0_0_0 = other_ops_6_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_0_1 = other_ops_6_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_0_2 = other_ops_6_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_7_0_1_0 = other_ops_6_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_7_0_1_1 = other_ops_6_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_7_0_1_2 = other_ops_6_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_7_0_2_0 = other_ops_6_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_7_0_2_1 = other_ops_6_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_7_0_2_2 = other_ops_6_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_8_0_0_0 = other_ops_7_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_8_0_0_1 = other_ops_7_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_8_0_0_2 = other_ops_7_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_8_0_1_0 = other_ops_7_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_8_0_1_1 = other_ops_7_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_8_0_1_2 = other_ops_7_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_8_0_2_0 = other_ops_7_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_8_0_2_1 = other_ops_7_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_8_0_2_2 = other_ops_7_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_9_0_0_0 = other_ops_8_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_9_0_0_1 = other_ops_8_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_9_0_0_2 = other_ops_8_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_9_0_1_0 = other_ops_8_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_9_0_1_1 = other_ops_8_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_9_0_1_2 = other_ops_8_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_9_0_2_0 = other_ops_8_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_9_0_2_1 = other_ops_8_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_9_0_2_2 = other_ops_8_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_10_0_0_0 = other_ops_9_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_10_0_0_1 = other_ops_9_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_10_0_0_2 = other_ops_9_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_10_0_1_0 = other_ops_9_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_10_0_1_1 = other_ops_9_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_10_0_1_2 = other_ops_9_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_10_0_2_0 = other_ops_9_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_10_0_2_1 = other_ops_9_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_10_0_2_2 = other_ops_9_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_11_0_0_0 = other_ops_10_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_11_0_0_1 = other_ops_10_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_11_0_0_2 = other_ops_10_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_11_0_1_0 = other_ops_10_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_11_0_1_1 = other_ops_10_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_11_0_1_2 = other_ops_10_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_11_0_2_0 = other_ops_10_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_11_0_2_1 = other_ops_10_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_11_0_2_2 = other_ops_10_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_12_0_0_0 = other_ops_11_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_12_0_0_1 = other_ops_11_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_12_0_0_2 = other_ops_11_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_12_0_1_0 = other_ops_11_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_12_0_1_1 = other_ops_11_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_12_0_1_2 = other_ops_11_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_12_0_2_0 = other_ops_11_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_12_0_2_1 = other_ops_11_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_12_0_2_2 = other_ops_11_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_13_0_0_0 = other_ops_12_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_13_0_0_1 = other_ops_12_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_13_0_0_2 = other_ops_12_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_13_0_1_0 = other_ops_12_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_13_0_1_1 = other_ops_12_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_13_0_1_2 = other_ops_12_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_13_0_2_0 = other_ops_12_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_13_0_2_1 = other_ops_12_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_13_0_2_2 = other_ops_12_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_14_0_0_0 = other_ops_13_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_14_0_0_1 = other_ops_13_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_14_0_0_2 = other_ops_13_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_14_0_1_0 = other_ops_13_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_14_0_1_1 = other_ops_13_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_14_0_1_2 = other_ops_13_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_14_0_2_0 = other_ops_13_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_14_0_2_1 = other_ops_13_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_14_0_2_2 = other_ops_13_O_0_2_2; // @[Map2S.scala 24:12]
  assign O_15_0_0_0 = other_ops_14_O_0_0_0; // @[Map2S.scala 24:12]
  assign O_15_0_0_1 = other_ops_14_O_0_0_1; // @[Map2S.scala 24:12]
  assign O_15_0_0_2 = other_ops_14_O_0_0_2; // @[Map2S.scala 24:12]
  assign O_15_0_1_0 = other_ops_14_O_0_1_0; // @[Map2S.scala 24:12]
  assign O_15_0_1_1 = other_ops_14_O_0_1_1; // @[Map2S.scala 24:12]
  assign O_15_0_1_2 = other_ops_14_O_0_1_2; // @[Map2S.scala 24:12]
  assign O_15_0_2_0 = other_ops_14_O_0_2_0; // @[Map2S.scala 24:12]
  assign O_15_0_2_1 = other_ops_14_O_0_2_1; // @[Map2S.scala 24:12]
  assign O_15_0_2_2 = other_ops_14_O_0_2_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0_0 = I0_0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_0_1 = I0_0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_0_2 = I0_0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1_0 = I0_0_0_1_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1_1 = I0_0_0_1_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1_2 = I0_0_0_1_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_0 = I1_0_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_1 = I1_0_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_2 = I1_0_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0_0 = I0_1_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_0_1 = I0_1_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_0_2 = I0_1_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1_0 = I0_1_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1_1 = I0_1_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1_2 = I0_1_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0_0 = I1_1_0_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_0_1 = I1_1_0_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_0_2 = I1_1_0_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0_0 = I0_2_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_0_1 = I0_2_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_0_2 = I0_2_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1_0 = I0_2_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1_1 = I0_2_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1_2 = I0_2_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0_0 = I1_2_0_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_0_1 = I1_2_0_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_0_2 = I1_2_0_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0_0 = I0_3_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_0_1 = I0_3_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_0_2 = I0_3_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1_0 = I0_3_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1_1 = I0_3_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1_2 = I0_3_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0_0 = I1_3_0_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_0_1 = I1_3_0_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_0_2 = I1_3_0_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0_0 = I0_4_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_0_1 = I0_4_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_0_2 = I0_4_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1_0 = I0_4_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1_1 = I0_4_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1_2 = I0_4_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0_0 = I1_4_0_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_0_1 = I1_4_0_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_0_2 = I1_4_0_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0_0 = I0_5_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_0_1 = I0_5_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_0_2 = I0_5_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1_0 = I0_5_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1_1 = I0_5_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1_2 = I0_5_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0_0 = I1_5_0_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_0_1 = I1_5_0_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_0_2 = I1_5_0_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0_0 = I0_6_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_0_1 = I0_6_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_0_2 = I0_6_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1_0 = I0_6_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1_1 = I0_6_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1_2 = I0_6_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0_0 = I1_6_0_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_0_1 = I1_6_0_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_0_2 = I1_6_0_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0_0 = I0_7_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_0_1 = I0_7_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_0_2 = I0_7_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1_0 = I0_7_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1_1 = I0_7_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1_2 = I0_7_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0_0 = I1_7_0_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_0_1 = I1_7_0_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_0_2 = I1_7_0_2; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0_0_0 = I0_8_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_0_1 = I0_8_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_0_2 = I0_8_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_1_0 = I0_8_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_1_1 = I0_8_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_1_2 = I0_8_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I1_0_0 = I1_8_0_0; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_0_1 = I1_8_0_1; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_0_2 = I1_8_0_2; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0_0_0 = I0_9_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_0_1 = I0_9_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_0_2 = I0_9_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_1_0 = I0_9_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_1_1 = I0_9_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_1_2 = I0_9_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I1_0_0 = I1_9_0_0; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_0_1 = I1_9_0_1; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_0_2 = I1_9_0_2; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0_0_0 = I0_10_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_0_1 = I0_10_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_0_2 = I0_10_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_1_0 = I0_10_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_1_1 = I0_10_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_1_2 = I0_10_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I1_0_0 = I1_10_0_0; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_0_1 = I1_10_0_1; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_0_2 = I1_10_0_2; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0_0_0 = I0_11_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_0_1 = I0_11_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_0_2 = I0_11_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_1_0 = I0_11_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_1_1 = I0_11_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_1_2 = I0_11_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I1_0_0 = I1_11_0_0; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_0_1 = I1_11_0_1; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_0_2 = I1_11_0_2; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0_0_0 = I0_12_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_0_1 = I0_12_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_0_2 = I0_12_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_1_0 = I0_12_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_1_1 = I0_12_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_1_2 = I0_12_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I1_0_0 = I1_12_0_0; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_0_1 = I1_12_0_1; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_0_2 = I1_12_0_2; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0_0_0 = I0_13_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_0_1 = I0_13_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_0_2 = I0_13_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_1_0 = I0_13_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_1_1 = I0_13_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_1_2 = I0_13_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I1_0_0 = I1_13_0_0; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_0_1 = I1_13_0_1; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_0_2 = I1_13_0_2; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0_0_0 = I0_14_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_0_1 = I0_14_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_0_2 = I0_14_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_1_0 = I0_14_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_1_1 = I0_14_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_1_2 = I0_14_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I1_0_0 = I1_14_0_0; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_0_1 = I1_14_0_1; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_0_2 = I1_14_0_2; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0_0_0 = I0_15_0_0_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_0_1 = I0_15_0_0_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_0_2 = I0_15_0_0_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_1_0 = I0_15_0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_1_1 = I0_15_0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_1_2 = I0_15_0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I1_0_0 = I1_15_0_0; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_0_1 = I1_15_0_1; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_0_2 = I1_15_0_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_7(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0_0,
  input  [7:0] I0_0_0_0_1,
  input  [7:0] I0_0_0_0_2,
  input  [7:0] I0_0_0_1_0,
  input  [7:0] I0_0_0_1_1,
  input  [7:0] I0_0_0_1_2,
  input  [7:0] I0_1_0_0_0,
  input  [7:0] I0_1_0_0_1,
  input  [7:0] I0_1_0_0_2,
  input  [7:0] I0_1_0_1_0,
  input  [7:0] I0_1_0_1_1,
  input  [7:0] I0_1_0_1_2,
  input  [7:0] I0_2_0_0_0,
  input  [7:0] I0_2_0_0_1,
  input  [7:0] I0_2_0_0_2,
  input  [7:0] I0_2_0_1_0,
  input  [7:0] I0_2_0_1_1,
  input  [7:0] I0_2_0_1_2,
  input  [7:0] I0_3_0_0_0,
  input  [7:0] I0_3_0_0_1,
  input  [7:0] I0_3_0_0_2,
  input  [7:0] I0_3_0_1_0,
  input  [7:0] I0_3_0_1_1,
  input  [7:0] I0_3_0_1_2,
  input  [7:0] I0_4_0_0_0,
  input  [7:0] I0_4_0_0_1,
  input  [7:0] I0_4_0_0_2,
  input  [7:0] I0_4_0_1_0,
  input  [7:0] I0_4_0_1_1,
  input  [7:0] I0_4_0_1_2,
  input  [7:0] I0_5_0_0_0,
  input  [7:0] I0_5_0_0_1,
  input  [7:0] I0_5_0_0_2,
  input  [7:0] I0_5_0_1_0,
  input  [7:0] I0_5_0_1_1,
  input  [7:0] I0_5_0_1_2,
  input  [7:0] I0_6_0_0_0,
  input  [7:0] I0_6_0_0_1,
  input  [7:0] I0_6_0_0_2,
  input  [7:0] I0_6_0_1_0,
  input  [7:0] I0_6_0_1_1,
  input  [7:0] I0_6_0_1_2,
  input  [7:0] I0_7_0_0_0,
  input  [7:0] I0_7_0_0_1,
  input  [7:0] I0_7_0_0_2,
  input  [7:0] I0_7_0_1_0,
  input  [7:0] I0_7_0_1_1,
  input  [7:0] I0_7_0_1_2,
  input  [7:0] I0_8_0_0_0,
  input  [7:0] I0_8_0_0_1,
  input  [7:0] I0_8_0_0_2,
  input  [7:0] I0_8_0_1_0,
  input  [7:0] I0_8_0_1_1,
  input  [7:0] I0_8_0_1_2,
  input  [7:0] I0_9_0_0_0,
  input  [7:0] I0_9_0_0_1,
  input  [7:0] I0_9_0_0_2,
  input  [7:0] I0_9_0_1_0,
  input  [7:0] I0_9_0_1_1,
  input  [7:0] I0_9_0_1_2,
  input  [7:0] I0_10_0_0_0,
  input  [7:0] I0_10_0_0_1,
  input  [7:0] I0_10_0_0_2,
  input  [7:0] I0_10_0_1_0,
  input  [7:0] I0_10_0_1_1,
  input  [7:0] I0_10_0_1_2,
  input  [7:0] I0_11_0_0_0,
  input  [7:0] I0_11_0_0_1,
  input  [7:0] I0_11_0_0_2,
  input  [7:0] I0_11_0_1_0,
  input  [7:0] I0_11_0_1_1,
  input  [7:0] I0_11_0_1_2,
  input  [7:0] I0_12_0_0_0,
  input  [7:0] I0_12_0_0_1,
  input  [7:0] I0_12_0_0_2,
  input  [7:0] I0_12_0_1_0,
  input  [7:0] I0_12_0_1_1,
  input  [7:0] I0_12_0_1_2,
  input  [7:0] I0_13_0_0_0,
  input  [7:0] I0_13_0_0_1,
  input  [7:0] I0_13_0_0_2,
  input  [7:0] I0_13_0_1_0,
  input  [7:0] I0_13_0_1_1,
  input  [7:0] I0_13_0_1_2,
  input  [7:0] I0_14_0_0_0,
  input  [7:0] I0_14_0_0_1,
  input  [7:0] I0_14_0_0_2,
  input  [7:0] I0_14_0_1_0,
  input  [7:0] I0_14_0_1_1,
  input  [7:0] I0_14_0_1_2,
  input  [7:0] I0_15_0_0_0,
  input  [7:0] I0_15_0_0_1,
  input  [7:0] I0_15_0_0_2,
  input  [7:0] I0_15_0_1_0,
  input  [7:0] I0_15_0_1_1,
  input  [7:0] I0_15_0_1_2,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_0_0_1,
  input  [7:0] I1_0_0_2,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_1_0_1,
  input  [7:0] I1_1_0_2,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_2_0_1,
  input  [7:0] I1_2_0_2,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_3_0_1,
  input  [7:0] I1_3_0_2,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_4_0_1,
  input  [7:0] I1_4_0_2,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_5_0_1,
  input  [7:0] I1_5_0_2,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_6_0_1,
  input  [7:0] I1_6_0_2,
  input  [7:0] I1_7_0_0,
  input  [7:0] I1_7_0_1,
  input  [7:0] I1_7_0_2,
  input  [7:0] I1_8_0_0,
  input  [7:0] I1_8_0_1,
  input  [7:0] I1_8_0_2,
  input  [7:0] I1_9_0_0,
  input  [7:0] I1_9_0_1,
  input  [7:0] I1_9_0_2,
  input  [7:0] I1_10_0_0,
  input  [7:0] I1_10_0_1,
  input  [7:0] I1_10_0_2,
  input  [7:0] I1_11_0_0,
  input  [7:0] I1_11_0_1,
  input  [7:0] I1_11_0_2,
  input  [7:0] I1_12_0_0,
  input  [7:0] I1_12_0_1,
  input  [7:0] I1_12_0_2,
  input  [7:0] I1_13_0_0,
  input  [7:0] I1_13_0_1,
  input  [7:0] I1_13_0_2,
  input  [7:0] I1_14_0_0,
  input  [7:0] I1_14_0_1,
  input  [7:0] I1_14_0_2,
  input  [7:0] I1_15_0_0,
  input  [7:0] I1_15_0_1,
  input  [7:0] I1_15_0_2,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_0_0_1_0,
  output [7:0] O_0_0_1_1,
  output [7:0] O_0_0_1_2,
  output [7:0] O_0_0_2_0,
  output [7:0] O_0_0_2_1,
  output [7:0] O_0_0_2_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_1_0_1_0,
  output [7:0] O_1_0_1_1,
  output [7:0] O_1_0_1_2,
  output [7:0] O_1_0_2_0,
  output [7:0] O_1_0_2_1,
  output [7:0] O_1_0_2_2,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_0_2,
  output [7:0] O_2_0_1_0,
  output [7:0] O_2_0_1_1,
  output [7:0] O_2_0_1_2,
  output [7:0] O_2_0_2_0,
  output [7:0] O_2_0_2_1,
  output [7:0] O_2_0_2_2,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_0_2,
  output [7:0] O_3_0_1_0,
  output [7:0] O_3_0_1_1,
  output [7:0] O_3_0_1_2,
  output [7:0] O_3_0_2_0,
  output [7:0] O_3_0_2_1,
  output [7:0] O_3_0_2_2,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_0_2,
  output [7:0] O_4_0_1_0,
  output [7:0] O_4_0_1_1,
  output [7:0] O_4_0_1_2,
  output [7:0] O_4_0_2_0,
  output [7:0] O_4_0_2_1,
  output [7:0] O_4_0_2_2,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_0_2,
  output [7:0] O_5_0_1_0,
  output [7:0] O_5_0_1_1,
  output [7:0] O_5_0_1_2,
  output [7:0] O_5_0_2_0,
  output [7:0] O_5_0_2_1,
  output [7:0] O_5_0_2_2,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_0_2,
  output [7:0] O_6_0_1_0,
  output [7:0] O_6_0_1_1,
  output [7:0] O_6_0_1_2,
  output [7:0] O_6_0_2_0,
  output [7:0] O_6_0_2_1,
  output [7:0] O_6_0_2_2,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_0_2,
  output [7:0] O_7_0_1_0,
  output [7:0] O_7_0_1_1,
  output [7:0] O_7_0_1_2,
  output [7:0] O_7_0_2_0,
  output [7:0] O_7_0_2_1,
  output [7:0] O_7_0_2_2,
  output [7:0] O_8_0_0_0,
  output [7:0] O_8_0_0_1,
  output [7:0] O_8_0_0_2,
  output [7:0] O_8_0_1_0,
  output [7:0] O_8_0_1_1,
  output [7:0] O_8_0_1_2,
  output [7:0] O_8_0_2_0,
  output [7:0] O_8_0_2_1,
  output [7:0] O_8_0_2_2,
  output [7:0] O_9_0_0_0,
  output [7:0] O_9_0_0_1,
  output [7:0] O_9_0_0_2,
  output [7:0] O_9_0_1_0,
  output [7:0] O_9_0_1_1,
  output [7:0] O_9_0_1_2,
  output [7:0] O_9_0_2_0,
  output [7:0] O_9_0_2_1,
  output [7:0] O_9_0_2_2,
  output [7:0] O_10_0_0_0,
  output [7:0] O_10_0_0_1,
  output [7:0] O_10_0_0_2,
  output [7:0] O_10_0_1_0,
  output [7:0] O_10_0_1_1,
  output [7:0] O_10_0_1_2,
  output [7:0] O_10_0_2_0,
  output [7:0] O_10_0_2_1,
  output [7:0] O_10_0_2_2,
  output [7:0] O_11_0_0_0,
  output [7:0] O_11_0_0_1,
  output [7:0] O_11_0_0_2,
  output [7:0] O_11_0_1_0,
  output [7:0] O_11_0_1_1,
  output [7:0] O_11_0_1_2,
  output [7:0] O_11_0_2_0,
  output [7:0] O_11_0_2_1,
  output [7:0] O_11_0_2_2,
  output [7:0] O_12_0_0_0,
  output [7:0] O_12_0_0_1,
  output [7:0] O_12_0_0_2,
  output [7:0] O_12_0_1_0,
  output [7:0] O_12_0_1_1,
  output [7:0] O_12_0_1_2,
  output [7:0] O_12_0_2_0,
  output [7:0] O_12_0_2_1,
  output [7:0] O_12_0_2_2,
  output [7:0] O_13_0_0_0,
  output [7:0] O_13_0_0_1,
  output [7:0] O_13_0_0_2,
  output [7:0] O_13_0_1_0,
  output [7:0] O_13_0_1_1,
  output [7:0] O_13_0_1_2,
  output [7:0] O_13_0_2_0,
  output [7:0] O_13_0_2_1,
  output [7:0] O_13_0_2_2,
  output [7:0] O_14_0_0_0,
  output [7:0] O_14_0_0_1,
  output [7:0] O_14_0_0_2,
  output [7:0] O_14_0_1_0,
  output [7:0] O_14_0_1_1,
  output [7:0] O_14_0_1_2,
  output [7:0] O_14_0_2_0,
  output [7:0] O_14_0_2_1,
  output [7:0] O_14_0_2_2,
  output [7:0] O_15_0_0_0,
  output [7:0] O_15_0_0_1,
  output [7:0] O_15_0_0_2,
  output [7:0] O_15_0_1_0,
  output [7:0] O_15_0_1_1,
  output [7:0] O_15_0_1_2,
  output [7:0] O_15_0_2_0,
  output [7:0] O_15_0_2_1,
  output [7:0] O_15_0_2_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_2_2; // @[Map2T.scala 8:20]
  Map2S_21 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0_0(op_I0_0_0_0_0),
    .I0_0_0_0_1(op_I0_0_0_0_1),
    .I0_0_0_0_2(op_I0_0_0_0_2),
    .I0_0_0_1_0(op_I0_0_0_1_0),
    .I0_0_0_1_1(op_I0_0_0_1_1),
    .I0_0_0_1_2(op_I0_0_0_1_2),
    .I0_1_0_0_0(op_I0_1_0_0_0),
    .I0_1_0_0_1(op_I0_1_0_0_1),
    .I0_1_0_0_2(op_I0_1_0_0_2),
    .I0_1_0_1_0(op_I0_1_0_1_0),
    .I0_1_0_1_1(op_I0_1_0_1_1),
    .I0_1_0_1_2(op_I0_1_0_1_2),
    .I0_2_0_0_0(op_I0_2_0_0_0),
    .I0_2_0_0_1(op_I0_2_0_0_1),
    .I0_2_0_0_2(op_I0_2_0_0_2),
    .I0_2_0_1_0(op_I0_2_0_1_0),
    .I0_2_0_1_1(op_I0_2_0_1_1),
    .I0_2_0_1_2(op_I0_2_0_1_2),
    .I0_3_0_0_0(op_I0_3_0_0_0),
    .I0_3_0_0_1(op_I0_3_0_0_1),
    .I0_3_0_0_2(op_I0_3_0_0_2),
    .I0_3_0_1_0(op_I0_3_0_1_0),
    .I0_3_0_1_1(op_I0_3_0_1_1),
    .I0_3_0_1_2(op_I0_3_0_1_2),
    .I0_4_0_0_0(op_I0_4_0_0_0),
    .I0_4_0_0_1(op_I0_4_0_0_1),
    .I0_4_0_0_2(op_I0_4_0_0_2),
    .I0_4_0_1_0(op_I0_4_0_1_0),
    .I0_4_0_1_1(op_I0_4_0_1_1),
    .I0_4_0_1_2(op_I0_4_0_1_2),
    .I0_5_0_0_0(op_I0_5_0_0_0),
    .I0_5_0_0_1(op_I0_5_0_0_1),
    .I0_5_0_0_2(op_I0_5_0_0_2),
    .I0_5_0_1_0(op_I0_5_0_1_0),
    .I0_5_0_1_1(op_I0_5_0_1_1),
    .I0_5_0_1_2(op_I0_5_0_1_2),
    .I0_6_0_0_0(op_I0_6_0_0_0),
    .I0_6_0_0_1(op_I0_6_0_0_1),
    .I0_6_0_0_2(op_I0_6_0_0_2),
    .I0_6_0_1_0(op_I0_6_0_1_0),
    .I0_6_0_1_1(op_I0_6_0_1_1),
    .I0_6_0_1_2(op_I0_6_0_1_2),
    .I0_7_0_0_0(op_I0_7_0_0_0),
    .I0_7_0_0_1(op_I0_7_0_0_1),
    .I0_7_0_0_2(op_I0_7_0_0_2),
    .I0_7_0_1_0(op_I0_7_0_1_0),
    .I0_7_0_1_1(op_I0_7_0_1_1),
    .I0_7_0_1_2(op_I0_7_0_1_2),
    .I0_8_0_0_0(op_I0_8_0_0_0),
    .I0_8_0_0_1(op_I0_8_0_0_1),
    .I0_8_0_0_2(op_I0_8_0_0_2),
    .I0_8_0_1_0(op_I0_8_0_1_0),
    .I0_8_0_1_1(op_I0_8_0_1_1),
    .I0_8_0_1_2(op_I0_8_0_1_2),
    .I0_9_0_0_0(op_I0_9_0_0_0),
    .I0_9_0_0_1(op_I0_9_0_0_1),
    .I0_9_0_0_2(op_I0_9_0_0_2),
    .I0_9_0_1_0(op_I0_9_0_1_0),
    .I0_9_0_1_1(op_I0_9_0_1_1),
    .I0_9_0_1_2(op_I0_9_0_1_2),
    .I0_10_0_0_0(op_I0_10_0_0_0),
    .I0_10_0_0_1(op_I0_10_0_0_1),
    .I0_10_0_0_2(op_I0_10_0_0_2),
    .I0_10_0_1_0(op_I0_10_0_1_0),
    .I0_10_0_1_1(op_I0_10_0_1_1),
    .I0_10_0_1_2(op_I0_10_0_1_2),
    .I0_11_0_0_0(op_I0_11_0_0_0),
    .I0_11_0_0_1(op_I0_11_0_0_1),
    .I0_11_0_0_2(op_I0_11_0_0_2),
    .I0_11_0_1_0(op_I0_11_0_1_0),
    .I0_11_0_1_1(op_I0_11_0_1_1),
    .I0_11_0_1_2(op_I0_11_0_1_2),
    .I0_12_0_0_0(op_I0_12_0_0_0),
    .I0_12_0_0_1(op_I0_12_0_0_1),
    .I0_12_0_0_2(op_I0_12_0_0_2),
    .I0_12_0_1_0(op_I0_12_0_1_0),
    .I0_12_0_1_1(op_I0_12_0_1_1),
    .I0_12_0_1_2(op_I0_12_0_1_2),
    .I0_13_0_0_0(op_I0_13_0_0_0),
    .I0_13_0_0_1(op_I0_13_0_0_1),
    .I0_13_0_0_2(op_I0_13_0_0_2),
    .I0_13_0_1_0(op_I0_13_0_1_0),
    .I0_13_0_1_1(op_I0_13_0_1_1),
    .I0_13_0_1_2(op_I0_13_0_1_2),
    .I0_14_0_0_0(op_I0_14_0_0_0),
    .I0_14_0_0_1(op_I0_14_0_0_1),
    .I0_14_0_0_2(op_I0_14_0_0_2),
    .I0_14_0_1_0(op_I0_14_0_1_0),
    .I0_14_0_1_1(op_I0_14_0_1_1),
    .I0_14_0_1_2(op_I0_14_0_1_2),
    .I0_15_0_0_0(op_I0_15_0_0_0),
    .I0_15_0_0_1(op_I0_15_0_0_1),
    .I0_15_0_0_2(op_I0_15_0_0_2),
    .I0_15_0_1_0(op_I0_15_0_1_0),
    .I0_15_0_1_1(op_I0_15_0_1_1),
    .I0_15_0_1_2(op_I0_15_0_1_2),
    .I1_0_0_0(op_I1_0_0_0),
    .I1_0_0_1(op_I1_0_0_1),
    .I1_0_0_2(op_I1_0_0_2),
    .I1_1_0_0(op_I1_1_0_0),
    .I1_1_0_1(op_I1_1_0_1),
    .I1_1_0_2(op_I1_1_0_2),
    .I1_2_0_0(op_I1_2_0_0),
    .I1_2_0_1(op_I1_2_0_1),
    .I1_2_0_2(op_I1_2_0_2),
    .I1_3_0_0(op_I1_3_0_0),
    .I1_3_0_1(op_I1_3_0_1),
    .I1_3_0_2(op_I1_3_0_2),
    .I1_4_0_0(op_I1_4_0_0),
    .I1_4_0_1(op_I1_4_0_1),
    .I1_4_0_2(op_I1_4_0_2),
    .I1_5_0_0(op_I1_5_0_0),
    .I1_5_0_1(op_I1_5_0_1),
    .I1_5_0_2(op_I1_5_0_2),
    .I1_6_0_0(op_I1_6_0_0),
    .I1_6_0_1(op_I1_6_0_1),
    .I1_6_0_2(op_I1_6_0_2),
    .I1_7_0_0(op_I1_7_0_0),
    .I1_7_0_1(op_I1_7_0_1),
    .I1_7_0_2(op_I1_7_0_2),
    .I1_8_0_0(op_I1_8_0_0),
    .I1_8_0_1(op_I1_8_0_1),
    .I1_8_0_2(op_I1_8_0_2),
    .I1_9_0_0(op_I1_9_0_0),
    .I1_9_0_1(op_I1_9_0_1),
    .I1_9_0_2(op_I1_9_0_2),
    .I1_10_0_0(op_I1_10_0_0),
    .I1_10_0_1(op_I1_10_0_1),
    .I1_10_0_2(op_I1_10_0_2),
    .I1_11_0_0(op_I1_11_0_0),
    .I1_11_0_1(op_I1_11_0_1),
    .I1_11_0_2(op_I1_11_0_2),
    .I1_12_0_0(op_I1_12_0_0),
    .I1_12_0_1(op_I1_12_0_1),
    .I1_12_0_2(op_I1_12_0_2),
    .I1_13_0_0(op_I1_13_0_0),
    .I1_13_0_1(op_I1_13_0_1),
    .I1_13_0_2(op_I1_13_0_2),
    .I1_14_0_0(op_I1_14_0_0),
    .I1_14_0_1(op_I1_14_0_1),
    .I1_14_0_2(op_I1_14_0_2),
    .I1_15_0_0(op_I1_15_0_0),
    .I1_15_0_1(op_I1_15_0_1),
    .I1_15_0_2(op_I1_15_0_2),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_0_0_0_2(op_O_0_0_0_2),
    .O_0_0_1_0(op_O_0_0_1_0),
    .O_0_0_1_1(op_O_0_0_1_1),
    .O_0_0_1_2(op_O_0_0_1_2),
    .O_0_0_2_0(op_O_0_0_2_0),
    .O_0_0_2_1(op_O_0_0_2_1),
    .O_0_0_2_2(op_O_0_0_2_2),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_1_0_0_2(op_O_1_0_0_2),
    .O_1_0_1_0(op_O_1_0_1_0),
    .O_1_0_1_1(op_O_1_0_1_1),
    .O_1_0_1_2(op_O_1_0_1_2),
    .O_1_0_2_0(op_O_1_0_2_0),
    .O_1_0_2_1(op_O_1_0_2_1),
    .O_1_0_2_2(op_O_1_0_2_2),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_2_0_0_2(op_O_2_0_0_2),
    .O_2_0_1_0(op_O_2_0_1_0),
    .O_2_0_1_1(op_O_2_0_1_1),
    .O_2_0_1_2(op_O_2_0_1_2),
    .O_2_0_2_0(op_O_2_0_2_0),
    .O_2_0_2_1(op_O_2_0_2_1),
    .O_2_0_2_2(op_O_2_0_2_2),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_3_0_0_2(op_O_3_0_0_2),
    .O_3_0_1_0(op_O_3_0_1_0),
    .O_3_0_1_1(op_O_3_0_1_1),
    .O_3_0_1_2(op_O_3_0_1_2),
    .O_3_0_2_0(op_O_3_0_2_0),
    .O_3_0_2_1(op_O_3_0_2_1),
    .O_3_0_2_2(op_O_3_0_2_2),
    .O_4_0_0_0(op_O_4_0_0_0),
    .O_4_0_0_1(op_O_4_0_0_1),
    .O_4_0_0_2(op_O_4_0_0_2),
    .O_4_0_1_0(op_O_4_0_1_0),
    .O_4_0_1_1(op_O_4_0_1_1),
    .O_4_0_1_2(op_O_4_0_1_2),
    .O_4_0_2_0(op_O_4_0_2_0),
    .O_4_0_2_1(op_O_4_0_2_1),
    .O_4_0_2_2(op_O_4_0_2_2),
    .O_5_0_0_0(op_O_5_0_0_0),
    .O_5_0_0_1(op_O_5_0_0_1),
    .O_5_0_0_2(op_O_5_0_0_2),
    .O_5_0_1_0(op_O_5_0_1_0),
    .O_5_0_1_1(op_O_5_0_1_1),
    .O_5_0_1_2(op_O_5_0_1_2),
    .O_5_0_2_0(op_O_5_0_2_0),
    .O_5_0_2_1(op_O_5_0_2_1),
    .O_5_0_2_2(op_O_5_0_2_2),
    .O_6_0_0_0(op_O_6_0_0_0),
    .O_6_0_0_1(op_O_6_0_0_1),
    .O_6_0_0_2(op_O_6_0_0_2),
    .O_6_0_1_0(op_O_6_0_1_0),
    .O_6_0_1_1(op_O_6_0_1_1),
    .O_6_0_1_2(op_O_6_0_1_2),
    .O_6_0_2_0(op_O_6_0_2_0),
    .O_6_0_2_1(op_O_6_0_2_1),
    .O_6_0_2_2(op_O_6_0_2_2),
    .O_7_0_0_0(op_O_7_0_0_0),
    .O_7_0_0_1(op_O_7_0_0_1),
    .O_7_0_0_2(op_O_7_0_0_2),
    .O_7_0_1_0(op_O_7_0_1_0),
    .O_7_0_1_1(op_O_7_0_1_1),
    .O_7_0_1_2(op_O_7_0_1_2),
    .O_7_0_2_0(op_O_7_0_2_0),
    .O_7_0_2_1(op_O_7_0_2_1),
    .O_7_0_2_2(op_O_7_0_2_2),
    .O_8_0_0_0(op_O_8_0_0_0),
    .O_8_0_0_1(op_O_8_0_0_1),
    .O_8_0_0_2(op_O_8_0_0_2),
    .O_8_0_1_0(op_O_8_0_1_0),
    .O_8_0_1_1(op_O_8_0_1_1),
    .O_8_0_1_2(op_O_8_0_1_2),
    .O_8_0_2_0(op_O_8_0_2_0),
    .O_8_0_2_1(op_O_8_0_2_1),
    .O_8_0_2_2(op_O_8_0_2_2),
    .O_9_0_0_0(op_O_9_0_0_0),
    .O_9_0_0_1(op_O_9_0_0_1),
    .O_9_0_0_2(op_O_9_0_0_2),
    .O_9_0_1_0(op_O_9_0_1_0),
    .O_9_0_1_1(op_O_9_0_1_1),
    .O_9_0_1_2(op_O_9_0_1_2),
    .O_9_0_2_0(op_O_9_0_2_0),
    .O_9_0_2_1(op_O_9_0_2_1),
    .O_9_0_2_2(op_O_9_0_2_2),
    .O_10_0_0_0(op_O_10_0_0_0),
    .O_10_0_0_1(op_O_10_0_0_1),
    .O_10_0_0_2(op_O_10_0_0_2),
    .O_10_0_1_0(op_O_10_0_1_0),
    .O_10_0_1_1(op_O_10_0_1_1),
    .O_10_0_1_2(op_O_10_0_1_2),
    .O_10_0_2_0(op_O_10_0_2_0),
    .O_10_0_2_1(op_O_10_0_2_1),
    .O_10_0_2_2(op_O_10_0_2_2),
    .O_11_0_0_0(op_O_11_0_0_0),
    .O_11_0_0_1(op_O_11_0_0_1),
    .O_11_0_0_2(op_O_11_0_0_2),
    .O_11_0_1_0(op_O_11_0_1_0),
    .O_11_0_1_1(op_O_11_0_1_1),
    .O_11_0_1_2(op_O_11_0_1_2),
    .O_11_0_2_0(op_O_11_0_2_0),
    .O_11_0_2_1(op_O_11_0_2_1),
    .O_11_0_2_2(op_O_11_0_2_2),
    .O_12_0_0_0(op_O_12_0_0_0),
    .O_12_0_0_1(op_O_12_0_0_1),
    .O_12_0_0_2(op_O_12_0_0_2),
    .O_12_0_1_0(op_O_12_0_1_0),
    .O_12_0_1_1(op_O_12_0_1_1),
    .O_12_0_1_2(op_O_12_0_1_2),
    .O_12_0_2_0(op_O_12_0_2_0),
    .O_12_0_2_1(op_O_12_0_2_1),
    .O_12_0_2_2(op_O_12_0_2_2),
    .O_13_0_0_0(op_O_13_0_0_0),
    .O_13_0_0_1(op_O_13_0_0_1),
    .O_13_0_0_2(op_O_13_0_0_2),
    .O_13_0_1_0(op_O_13_0_1_0),
    .O_13_0_1_1(op_O_13_0_1_1),
    .O_13_0_1_2(op_O_13_0_1_2),
    .O_13_0_2_0(op_O_13_0_2_0),
    .O_13_0_2_1(op_O_13_0_2_1),
    .O_13_0_2_2(op_O_13_0_2_2),
    .O_14_0_0_0(op_O_14_0_0_0),
    .O_14_0_0_1(op_O_14_0_0_1),
    .O_14_0_0_2(op_O_14_0_0_2),
    .O_14_0_1_0(op_O_14_0_1_0),
    .O_14_0_1_1(op_O_14_0_1_1),
    .O_14_0_1_2(op_O_14_0_1_2),
    .O_14_0_2_0(op_O_14_0_2_0),
    .O_14_0_2_1(op_O_14_0_2_1),
    .O_14_0_2_2(op_O_14_0_2_2),
    .O_15_0_0_0(op_O_15_0_0_0),
    .O_15_0_0_1(op_O_15_0_0_1),
    .O_15_0_0_2(op_O_15_0_0_2),
    .O_15_0_1_0(op_O_15_0_1_0),
    .O_15_0_1_1(op_O_15_0_1_1),
    .O_15_0_1_2(op_O_15_0_1_2),
    .O_15_0_2_0(op_O_15_0_2_0),
    .O_15_0_2_1(op_O_15_0_2_1),
    .O_15_0_2_2(op_O_15_0_2_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_0_2 = op_O_0_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_0_1_0 = op_O_0_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_0_1_1 = op_O_0_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_0_1_2 = op_O_0_0_1_2; // @[Map2T.scala 17:7]
  assign O_0_0_2_0 = op_O_0_0_2_0; // @[Map2T.scala 17:7]
  assign O_0_0_2_1 = op_O_0_0_2_1; // @[Map2T.scala 17:7]
  assign O_0_0_2_2 = op_O_0_0_2_2; // @[Map2T.scala 17:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_0_2 = op_O_1_0_0_2; // @[Map2T.scala 17:7]
  assign O_1_0_1_0 = op_O_1_0_1_0; // @[Map2T.scala 17:7]
  assign O_1_0_1_1 = op_O_1_0_1_1; // @[Map2T.scala 17:7]
  assign O_1_0_1_2 = op_O_1_0_1_2; // @[Map2T.scala 17:7]
  assign O_1_0_2_0 = op_O_1_0_2_0; // @[Map2T.scala 17:7]
  assign O_1_0_2_1 = op_O_1_0_2_1; // @[Map2T.scala 17:7]
  assign O_1_0_2_2 = op_O_1_0_2_2; // @[Map2T.scala 17:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_0_2 = op_O_2_0_0_2; // @[Map2T.scala 17:7]
  assign O_2_0_1_0 = op_O_2_0_1_0; // @[Map2T.scala 17:7]
  assign O_2_0_1_1 = op_O_2_0_1_1; // @[Map2T.scala 17:7]
  assign O_2_0_1_2 = op_O_2_0_1_2; // @[Map2T.scala 17:7]
  assign O_2_0_2_0 = op_O_2_0_2_0; // @[Map2T.scala 17:7]
  assign O_2_0_2_1 = op_O_2_0_2_1; // @[Map2T.scala 17:7]
  assign O_2_0_2_2 = op_O_2_0_2_2; // @[Map2T.scala 17:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_0_2 = op_O_3_0_0_2; // @[Map2T.scala 17:7]
  assign O_3_0_1_0 = op_O_3_0_1_0; // @[Map2T.scala 17:7]
  assign O_3_0_1_1 = op_O_3_0_1_1; // @[Map2T.scala 17:7]
  assign O_3_0_1_2 = op_O_3_0_1_2; // @[Map2T.scala 17:7]
  assign O_3_0_2_0 = op_O_3_0_2_0; // @[Map2T.scala 17:7]
  assign O_3_0_2_1 = op_O_3_0_2_1; // @[Map2T.scala 17:7]
  assign O_3_0_2_2 = op_O_3_0_2_2; // @[Map2T.scala 17:7]
  assign O_4_0_0_0 = op_O_4_0_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_0_1 = op_O_4_0_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_0_2 = op_O_4_0_0_2; // @[Map2T.scala 17:7]
  assign O_4_0_1_0 = op_O_4_0_1_0; // @[Map2T.scala 17:7]
  assign O_4_0_1_1 = op_O_4_0_1_1; // @[Map2T.scala 17:7]
  assign O_4_0_1_2 = op_O_4_0_1_2; // @[Map2T.scala 17:7]
  assign O_4_0_2_0 = op_O_4_0_2_0; // @[Map2T.scala 17:7]
  assign O_4_0_2_1 = op_O_4_0_2_1; // @[Map2T.scala 17:7]
  assign O_4_0_2_2 = op_O_4_0_2_2; // @[Map2T.scala 17:7]
  assign O_5_0_0_0 = op_O_5_0_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_0_1 = op_O_5_0_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_0_2 = op_O_5_0_0_2; // @[Map2T.scala 17:7]
  assign O_5_0_1_0 = op_O_5_0_1_0; // @[Map2T.scala 17:7]
  assign O_5_0_1_1 = op_O_5_0_1_1; // @[Map2T.scala 17:7]
  assign O_5_0_1_2 = op_O_5_0_1_2; // @[Map2T.scala 17:7]
  assign O_5_0_2_0 = op_O_5_0_2_0; // @[Map2T.scala 17:7]
  assign O_5_0_2_1 = op_O_5_0_2_1; // @[Map2T.scala 17:7]
  assign O_5_0_2_2 = op_O_5_0_2_2; // @[Map2T.scala 17:7]
  assign O_6_0_0_0 = op_O_6_0_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_0_1 = op_O_6_0_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_0_2 = op_O_6_0_0_2; // @[Map2T.scala 17:7]
  assign O_6_0_1_0 = op_O_6_0_1_0; // @[Map2T.scala 17:7]
  assign O_6_0_1_1 = op_O_6_0_1_1; // @[Map2T.scala 17:7]
  assign O_6_0_1_2 = op_O_6_0_1_2; // @[Map2T.scala 17:7]
  assign O_6_0_2_0 = op_O_6_0_2_0; // @[Map2T.scala 17:7]
  assign O_6_0_2_1 = op_O_6_0_2_1; // @[Map2T.scala 17:7]
  assign O_6_0_2_2 = op_O_6_0_2_2; // @[Map2T.scala 17:7]
  assign O_7_0_0_0 = op_O_7_0_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_0_1 = op_O_7_0_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_0_2 = op_O_7_0_0_2; // @[Map2T.scala 17:7]
  assign O_7_0_1_0 = op_O_7_0_1_0; // @[Map2T.scala 17:7]
  assign O_7_0_1_1 = op_O_7_0_1_1; // @[Map2T.scala 17:7]
  assign O_7_0_1_2 = op_O_7_0_1_2; // @[Map2T.scala 17:7]
  assign O_7_0_2_0 = op_O_7_0_2_0; // @[Map2T.scala 17:7]
  assign O_7_0_2_1 = op_O_7_0_2_1; // @[Map2T.scala 17:7]
  assign O_7_0_2_2 = op_O_7_0_2_2; // @[Map2T.scala 17:7]
  assign O_8_0_0_0 = op_O_8_0_0_0; // @[Map2T.scala 17:7]
  assign O_8_0_0_1 = op_O_8_0_0_1; // @[Map2T.scala 17:7]
  assign O_8_0_0_2 = op_O_8_0_0_2; // @[Map2T.scala 17:7]
  assign O_8_0_1_0 = op_O_8_0_1_0; // @[Map2T.scala 17:7]
  assign O_8_0_1_1 = op_O_8_0_1_1; // @[Map2T.scala 17:7]
  assign O_8_0_1_2 = op_O_8_0_1_2; // @[Map2T.scala 17:7]
  assign O_8_0_2_0 = op_O_8_0_2_0; // @[Map2T.scala 17:7]
  assign O_8_0_2_1 = op_O_8_0_2_1; // @[Map2T.scala 17:7]
  assign O_8_0_2_2 = op_O_8_0_2_2; // @[Map2T.scala 17:7]
  assign O_9_0_0_0 = op_O_9_0_0_0; // @[Map2T.scala 17:7]
  assign O_9_0_0_1 = op_O_9_0_0_1; // @[Map2T.scala 17:7]
  assign O_9_0_0_2 = op_O_9_0_0_2; // @[Map2T.scala 17:7]
  assign O_9_0_1_0 = op_O_9_0_1_0; // @[Map2T.scala 17:7]
  assign O_9_0_1_1 = op_O_9_0_1_1; // @[Map2T.scala 17:7]
  assign O_9_0_1_2 = op_O_9_0_1_2; // @[Map2T.scala 17:7]
  assign O_9_0_2_0 = op_O_9_0_2_0; // @[Map2T.scala 17:7]
  assign O_9_0_2_1 = op_O_9_0_2_1; // @[Map2T.scala 17:7]
  assign O_9_0_2_2 = op_O_9_0_2_2; // @[Map2T.scala 17:7]
  assign O_10_0_0_0 = op_O_10_0_0_0; // @[Map2T.scala 17:7]
  assign O_10_0_0_1 = op_O_10_0_0_1; // @[Map2T.scala 17:7]
  assign O_10_0_0_2 = op_O_10_0_0_2; // @[Map2T.scala 17:7]
  assign O_10_0_1_0 = op_O_10_0_1_0; // @[Map2T.scala 17:7]
  assign O_10_0_1_1 = op_O_10_0_1_1; // @[Map2T.scala 17:7]
  assign O_10_0_1_2 = op_O_10_0_1_2; // @[Map2T.scala 17:7]
  assign O_10_0_2_0 = op_O_10_0_2_0; // @[Map2T.scala 17:7]
  assign O_10_0_2_1 = op_O_10_0_2_1; // @[Map2T.scala 17:7]
  assign O_10_0_2_2 = op_O_10_0_2_2; // @[Map2T.scala 17:7]
  assign O_11_0_0_0 = op_O_11_0_0_0; // @[Map2T.scala 17:7]
  assign O_11_0_0_1 = op_O_11_0_0_1; // @[Map2T.scala 17:7]
  assign O_11_0_0_2 = op_O_11_0_0_2; // @[Map2T.scala 17:7]
  assign O_11_0_1_0 = op_O_11_0_1_0; // @[Map2T.scala 17:7]
  assign O_11_0_1_1 = op_O_11_0_1_1; // @[Map2T.scala 17:7]
  assign O_11_0_1_2 = op_O_11_0_1_2; // @[Map2T.scala 17:7]
  assign O_11_0_2_0 = op_O_11_0_2_0; // @[Map2T.scala 17:7]
  assign O_11_0_2_1 = op_O_11_0_2_1; // @[Map2T.scala 17:7]
  assign O_11_0_2_2 = op_O_11_0_2_2; // @[Map2T.scala 17:7]
  assign O_12_0_0_0 = op_O_12_0_0_0; // @[Map2T.scala 17:7]
  assign O_12_0_0_1 = op_O_12_0_0_1; // @[Map2T.scala 17:7]
  assign O_12_0_0_2 = op_O_12_0_0_2; // @[Map2T.scala 17:7]
  assign O_12_0_1_0 = op_O_12_0_1_0; // @[Map2T.scala 17:7]
  assign O_12_0_1_1 = op_O_12_0_1_1; // @[Map2T.scala 17:7]
  assign O_12_0_1_2 = op_O_12_0_1_2; // @[Map2T.scala 17:7]
  assign O_12_0_2_0 = op_O_12_0_2_0; // @[Map2T.scala 17:7]
  assign O_12_0_2_1 = op_O_12_0_2_1; // @[Map2T.scala 17:7]
  assign O_12_0_2_2 = op_O_12_0_2_2; // @[Map2T.scala 17:7]
  assign O_13_0_0_0 = op_O_13_0_0_0; // @[Map2T.scala 17:7]
  assign O_13_0_0_1 = op_O_13_0_0_1; // @[Map2T.scala 17:7]
  assign O_13_0_0_2 = op_O_13_0_0_2; // @[Map2T.scala 17:7]
  assign O_13_0_1_0 = op_O_13_0_1_0; // @[Map2T.scala 17:7]
  assign O_13_0_1_1 = op_O_13_0_1_1; // @[Map2T.scala 17:7]
  assign O_13_0_1_2 = op_O_13_0_1_2; // @[Map2T.scala 17:7]
  assign O_13_0_2_0 = op_O_13_0_2_0; // @[Map2T.scala 17:7]
  assign O_13_0_2_1 = op_O_13_0_2_1; // @[Map2T.scala 17:7]
  assign O_13_0_2_2 = op_O_13_0_2_2; // @[Map2T.scala 17:7]
  assign O_14_0_0_0 = op_O_14_0_0_0; // @[Map2T.scala 17:7]
  assign O_14_0_0_1 = op_O_14_0_0_1; // @[Map2T.scala 17:7]
  assign O_14_0_0_2 = op_O_14_0_0_2; // @[Map2T.scala 17:7]
  assign O_14_0_1_0 = op_O_14_0_1_0; // @[Map2T.scala 17:7]
  assign O_14_0_1_1 = op_O_14_0_1_1; // @[Map2T.scala 17:7]
  assign O_14_0_1_2 = op_O_14_0_1_2; // @[Map2T.scala 17:7]
  assign O_14_0_2_0 = op_O_14_0_2_0; // @[Map2T.scala 17:7]
  assign O_14_0_2_1 = op_O_14_0_2_1; // @[Map2T.scala 17:7]
  assign O_14_0_2_2 = op_O_14_0_2_2; // @[Map2T.scala 17:7]
  assign O_15_0_0_0 = op_O_15_0_0_0; // @[Map2T.scala 17:7]
  assign O_15_0_0_1 = op_O_15_0_0_1; // @[Map2T.scala 17:7]
  assign O_15_0_0_2 = op_O_15_0_0_2; // @[Map2T.scala 17:7]
  assign O_15_0_1_0 = op_O_15_0_1_0; // @[Map2T.scala 17:7]
  assign O_15_0_1_1 = op_O_15_0_1_1; // @[Map2T.scala 17:7]
  assign O_15_0_1_2 = op_O_15_0_1_2; // @[Map2T.scala 17:7]
  assign O_15_0_2_0 = op_O_15_0_2_0; // @[Map2T.scala 17:7]
  assign O_15_0_2_1 = op_O_15_0_2_1; // @[Map2T.scala 17:7]
  assign O_15_0_2_2 = op_O_15_0_2_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0_0 = I0_0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_0_1 = I0_0_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_0_0_2 = I0_0_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1_0 = I0_0_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1_1 = I0_0_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1_2 = I0_0_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0_0 = I0_1_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0_1 = I0_1_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0_2 = I0_1_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1_0 = I0_1_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1_1 = I0_1_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1_2 = I0_1_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0_0 = I0_2_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0_1 = I0_2_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0_2 = I0_2_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1_0 = I0_2_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1_1 = I0_2_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1_2 = I0_2_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0_0 = I0_3_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0_1 = I0_3_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0_2 = I0_3_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1_0 = I0_3_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1_1 = I0_3_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1_2 = I0_3_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0_0 = I0_4_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0_1 = I0_4_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0_2 = I0_4_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0_1_0 = I0_4_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_1_1 = I0_4_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0_1_2 = I0_4_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0_0 = I0_5_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0_1 = I0_5_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0_2 = I0_5_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0_1_0 = I0_5_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_1_1 = I0_5_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0_1_2 = I0_5_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0_0 = I0_6_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0_1 = I0_6_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0_2 = I0_6_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0_1_0 = I0_6_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_1_1 = I0_6_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0_1_2 = I0_6_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0_0 = I0_7_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0_1 = I0_7_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0_2 = I0_7_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0_1_0 = I0_7_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_1_1 = I0_7_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0_1_2 = I0_7_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_8_0_0_0 = I0_8_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_8_0_0_1 = I0_8_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_8_0_0_2 = I0_8_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_8_0_1_0 = I0_8_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_8_0_1_1 = I0_8_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_8_0_1_2 = I0_8_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_9_0_0_0 = I0_9_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_9_0_0_1 = I0_9_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_9_0_0_2 = I0_9_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_9_0_1_0 = I0_9_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_9_0_1_1 = I0_9_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_9_0_1_2 = I0_9_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_10_0_0_0 = I0_10_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_10_0_0_1 = I0_10_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_10_0_0_2 = I0_10_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_10_0_1_0 = I0_10_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_10_0_1_1 = I0_10_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_10_0_1_2 = I0_10_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_11_0_0_0 = I0_11_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_11_0_0_1 = I0_11_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_11_0_0_2 = I0_11_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_11_0_1_0 = I0_11_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_11_0_1_1 = I0_11_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_11_0_1_2 = I0_11_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_12_0_0_0 = I0_12_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_12_0_0_1 = I0_12_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_12_0_0_2 = I0_12_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_12_0_1_0 = I0_12_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_12_0_1_1 = I0_12_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_12_0_1_2 = I0_12_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_13_0_0_0 = I0_13_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_13_0_0_1 = I0_13_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_13_0_0_2 = I0_13_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_13_0_1_0 = I0_13_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_13_0_1_1 = I0_13_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_13_0_1_2 = I0_13_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_14_0_0_0 = I0_14_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_14_0_0_1 = I0_14_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_14_0_0_2 = I0_14_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_14_0_1_0 = I0_14_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_14_0_1_1 = I0_14_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_14_0_1_2 = I0_14_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_15_0_0_0 = I0_15_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_15_0_0_1 = I0_15_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_15_0_0_2 = I0_15_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_15_0_1_0 = I0_15_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_15_0_1_1 = I0_15_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_15_0_1_2 = I0_15_0_1_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0_0 = I1_0_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_0_1 = I1_0_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_0_2 = I1_0_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0_0 = I1_1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_1_0_1 = I1_1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_1_0_2 = I1_1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0_0 = I1_2_0_0; // @[Map2T.scala 16:11]
  assign op_I1_2_0_1 = I1_2_0_1; // @[Map2T.scala 16:11]
  assign op_I1_2_0_2 = I1_2_0_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0_0 = I1_3_0_0; // @[Map2T.scala 16:11]
  assign op_I1_3_0_1 = I1_3_0_1; // @[Map2T.scala 16:11]
  assign op_I1_3_0_2 = I1_3_0_2; // @[Map2T.scala 16:11]
  assign op_I1_4_0_0 = I1_4_0_0; // @[Map2T.scala 16:11]
  assign op_I1_4_0_1 = I1_4_0_1; // @[Map2T.scala 16:11]
  assign op_I1_4_0_2 = I1_4_0_2; // @[Map2T.scala 16:11]
  assign op_I1_5_0_0 = I1_5_0_0; // @[Map2T.scala 16:11]
  assign op_I1_5_0_1 = I1_5_0_1; // @[Map2T.scala 16:11]
  assign op_I1_5_0_2 = I1_5_0_2; // @[Map2T.scala 16:11]
  assign op_I1_6_0_0 = I1_6_0_0; // @[Map2T.scala 16:11]
  assign op_I1_6_0_1 = I1_6_0_1; // @[Map2T.scala 16:11]
  assign op_I1_6_0_2 = I1_6_0_2; // @[Map2T.scala 16:11]
  assign op_I1_7_0_0 = I1_7_0_0; // @[Map2T.scala 16:11]
  assign op_I1_7_0_1 = I1_7_0_1; // @[Map2T.scala 16:11]
  assign op_I1_7_0_2 = I1_7_0_2; // @[Map2T.scala 16:11]
  assign op_I1_8_0_0 = I1_8_0_0; // @[Map2T.scala 16:11]
  assign op_I1_8_0_1 = I1_8_0_1; // @[Map2T.scala 16:11]
  assign op_I1_8_0_2 = I1_8_0_2; // @[Map2T.scala 16:11]
  assign op_I1_9_0_0 = I1_9_0_0; // @[Map2T.scala 16:11]
  assign op_I1_9_0_1 = I1_9_0_1; // @[Map2T.scala 16:11]
  assign op_I1_9_0_2 = I1_9_0_2; // @[Map2T.scala 16:11]
  assign op_I1_10_0_0 = I1_10_0_0; // @[Map2T.scala 16:11]
  assign op_I1_10_0_1 = I1_10_0_1; // @[Map2T.scala 16:11]
  assign op_I1_10_0_2 = I1_10_0_2; // @[Map2T.scala 16:11]
  assign op_I1_11_0_0 = I1_11_0_0; // @[Map2T.scala 16:11]
  assign op_I1_11_0_1 = I1_11_0_1; // @[Map2T.scala 16:11]
  assign op_I1_11_0_2 = I1_11_0_2; // @[Map2T.scala 16:11]
  assign op_I1_12_0_0 = I1_12_0_0; // @[Map2T.scala 16:11]
  assign op_I1_12_0_1 = I1_12_0_1; // @[Map2T.scala 16:11]
  assign op_I1_12_0_2 = I1_12_0_2; // @[Map2T.scala 16:11]
  assign op_I1_13_0_0 = I1_13_0_0; // @[Map2T.scala 16:11]
  assign op_I1_13_0_1 = I1_13_0_1; // @[Map2T.scala 16:11]
  assign op_I1_13_0_2 = I1_13_0_2; // @[Map2T.scala 16:11]
  assign op_I1_14_0_0 = I1_14_0_0; // @[Map2T.scala 16:11]
  assign op_I1_14_0_1 = I1_14_0_1; // @[Map2T.scala 16:11]
  assign op_I1_14_0_2 = I1_14_0_2; // @[Map2T.scala 16:11]
  assign op_I1_15_0_0 = I1_15_0_0; // @[Map2T.scala 16:11]
  assign op_I1_15_0_1 = I1_15_0_1; // @[Map2T.scala 16:11]
  assign op_I1_15_0_2 = I1_15_0_2; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleToSSeq_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0_0 = I_0_0; // @[Tuple.scala 41:5]
  assign O_0_1 = I_0_1; // @[Tuple.scala 41:5]
  assign O_0_2 = I_0_2; // @[Tuple.scala 41:5]
  assign O_1_0 = I_1_0; // @[Tuple.scala 41:5]
  assign O_1_1 = I_1_1; // @[Tuple.scala 41:5]
  assign O_1_2 = I_1_2; // @[Tuple.scala 41:5]
  assign O_2_0 = I_2_0; // @[Tuple.scala 41:5]
  assign O_2_1 = I_2_1; // @[Tuple.scala 41:5]
  assign O_2_2 = I_2_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_3 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0_0(op_inst_I_0_0),
    .I_0_1(op_inst_I_0_1),
    .I_0_2(op_inst_I_0_2),
    .I_1_0(op_inst_I_1_0),
    .I_1_1(op_inst_I_1_1),
    .I_1_2(op_inst_I_1_2),
    .I_2_0(op_inst_I_2_0),
    .I_2_1(op_inst_I_2_1),
    .I_2_2(op_inst_I_2_2),
    .O_0_0(op_inst_O_0_0),
    .O_0_1(op_inst_O_0_1),
    .O_0_2(op_inst_O_0_2),
    .O_1_0(op_inst_O_1_0),
    .O_1_1(op_inst_O_1_1),
    .O_1_2(op_inst_O_1_2),
    .O_2_0(op_inst_O_2_0),
    .O_2_1(op_inst_O_2_1),
    .O_2_2(op_inst_O_2_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0_0 = op_inst_O_0_0; // @[Remove1S.scala 14:5]
  assign O_0_1 = op_inst_O_0_1; // @[Remove1S.scala 14:5]
  assign O_0_2 = op_inst_O_0_2; // @[Remove1S.scala 14:5]
  assign O_1_0 = op_inst_O_1_0; // @[Remove1S.scala 14:5]
  assign O_1_1 = op_inst_O_1_1; // @[Remove1S.scala 14:5]
  assign O_1_2 = op_inst_O_1_2; // @[Remove1S.scala 14:5]
  assign O_2_0 = op_inst_O_2_0; // @[Remove1S.scala 14:5]
  assign O_2_1 = op_inst_O_2_1; // @[Remove1S.scala 14:5]
  assign O_2_2 = op_inst_O_2_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0_0 = I_0_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_1 = I_0_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_2 = I_0_0_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_0 = I_0_1_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_1 = I_0_1_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_2 = I_0_1_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_0 = I_0_2_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_1 = I_0_2_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_2 = I_0_2_2; // @[Remove1S.scala 13:13]
endmodule
module MapS_6(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0_0,
  input  [7:0] I_0_0_0_1,
  input  [7:0] I_0_0_0_2,
  input  [7:0] I_0_0_1_0,
  input  [7:0] I_0_0_1_1,
  input  [7:0] I_0_0_1_2,
  input  [7:0] I_0_0_2_0,
  input  [7:0] I_0_0_2_1,
  input  [7:0] I_0_0_2_2,
  input  [7:0] I_1_0_0_0,
  input  [7:0] I_1_0_0_1,
  input  [7:0] I_1_0_0_2,
  input  [7:0] I_1_0_1_0,
  input  [7:0] I_1_0_1_1,
  input  [7:0] I_1_0_1_2,
  input  [7:0] I_1_0_2_0,
  input  [7:0] I_1_0_2_1,
  input  [7:0] I_1_0_2_2,
  input  [7:0] I_2_0_0_0,
  input  [7:0] I_2_0_0_1,
  input  [7:0] I_2_0_0_2,
  input  [7:0] I_2_0_1_0,
  input  [7:0] I_2_0_1_1,
  input  [7:0] I_2_0_1_2,
  input  [7:0] I_2_0_2_0,
  input  [7:0] I_2_0_2_1,
  input  [7:0] I_2_0_2_2,
  input  [7:0] I_3_0_0_0,
  input  [7:0] I_3_0_0_1,
  input  [7:0] I_3_0_0_2,
  input  [7:0] I_3_0_1_0,
  input  [7:0] I_3_0_1_1,
  input  [7:0] I_3_0_1_2,
  input  [7:0] I_3_0_2_0,
  input  [7:0] I_3_0_2_1,
  input  [7:0] I_3_0_2_2,
  input  [7:0] I_4_0_0_0,
  input  [7:0] I_4_0_0_1,
  input  [7:0] I_4_0_0_2,
  input  [7:0] I_4_0_1_0,
  input  [7:0] I_4_0_1_1,
  input  [7:0] I_4_0_1_2,
  input  [7:0] I_4_0_2_0,
  input  [7:0] I_4_0_2_1,
  input  [7:0] I_4_0_2_2,
  input  [7:0] I_5_0_0_0,
  input  [7:0] I_5_0_0_1,
  input  [7:0] I_5_0_0_2,
  input  [7:0] I_5_0_1_0,
  input  [7:0] I_5_0_1_1,
  input  [7:0] I_5_0_1_2,
  input  [7:0] I_5_0_2_0,
  input  [7:0] I_5_0_2_1,
  input  [7:0] I_5_0_2_2,
  input  [7:0] I_6_0_0_0,
  input  [7:0] I_6_0_0_1,
  input  [7:0] I_6_0_0_2,
  input  [7:0] I_6_0_1_0,
  input  [7:0] I_6_0_1_1,
  input  [7:0] I_6_0_1_2,
  input  [7:0] I_6_0_2_0,
  input  [7:0] I_6_0_2_1,
  input  [7:0] I_6_0_2_2,
  input  [7:0] I_7_0_0_0,
  input  [7:0] I_7_0_0_1,
  input  [7:0] I_7_0_0_2,
  input  [7:0] I_7_0_1_0,
  input  [7:0] I_7_0_1_1,
  input  [7:0] I_7_0_1_2,
  input  [7:0] I_7_0_2_0,
  input  [7:0] I_7_0_2_1,
  input  [7:0] I_7_0_2_2,
  input  [7:0] I_8_0_0_0,
  input  [7:0] I_8_0_0_1,
  input  [7:0] I_8_0_0_2,
  input  [7:0] I_8_0_1_0,
  input  [7:0] I_8_0_1_1,
  input  [7:0] I_8_0_1_2,
  input  [7:0] I_8_0_2_0,
  input  [7:0] I_8_0_2_1,
  input  [7:0] I_8_0_2_2,
  input  [7:0] I_9_0_0_0,
  input  [7:0] I_9_0_0_1,
  input  [7:0] I_9_0_0_2,
  input  [7:0] I_9_0_1_0,
  input  [7:0] I_9_0_1_1,
  input  [7:0] I_9_0_1_2,
  input  [7:0] I_9_0_2_0,
  input  [7:0] I_9_0_2_1,
  input  [7:0] I_9_0_2_2,
  input  [7:0] I_10_0_0_0,
  input  [7:0] I_10_0_0_1,
  input  [7:0] I_10_0_0_2,
  input  [7:0] I_10_0_1_0,
  input  [7:0] I_10_0_1_1,
  input  [7:0] I_10_0_1_2,
  input  [7:0] I_10_0_2_0,
  input  [7:0] I_10_0_2_1,
  input  [7:0] I_10_0_2_2,
  input  [7:0] I_11_0_0_0,
  input  [7:0] I_11_0_0_1,
  input  [7:0] I_11_0_0_2,
  input  [7:0] I_11_0_1_0,
  input  [7:0] I_11_0_1_1,
  input  [7:0] I_11_0_1_2,
  input  [7:0] I_11_0_2_0,
  input  [7:0] I_11_0_2_1,
  input  [7:0] I_11_0_2_2,
  input  [7:0] I_12_0_0_0,
  input  [7:0] I_12_0_0_1,
  input  [7:0] I_12_0_0_2,
  input  [7:0] I_12_0_1_0,
  input  [7:0] I_12_0_1_1,
  input  [7:0] I_12_0_1_2,
  input  [7:0] I_12_0_2_0,
  input  [7:0] I_12_0_2_1,
  input  [7:0] I_12_0_2_2,
  input  [7:0] I_13_0_0_0,
  input  [7:0] I_13_0_0_1,
  input  [7:0] I_13_0_0_2,
  input  [7:0] I_13_0_1_0,
  input  [7:0] I_13_0_1_1,
  input  [7:0] I_13_0_1_2,
  input  [7:0] I_13_0_2_0,
  input  [7:0] I_13_0_2_1,
  input  [7:0] I_13_0_2_2,
  input  [7:0] I_14_0_0_0,
  input  [7:0] I_14_0_0_1,
  input  [7:0] I_14_0_0_2,
  input  [7:0] I_14_0_1_0,
  input  [7:0] I_14_0_1_1,
  input  [7:0] I_14_0_1_2,
  input  [7:0] I_14_0_2_0,
  input  [7:0] I_14_0_2_1,
  input  [7:0] I_14_0_2_2,
  input  [7:0] I_15_0_0_0,
  input  [7:0] I_15_0_0_1,
  input  [7:0] I_15_0_0_2,
  input  [7:0] I_15_0_1_0,
  input  [7:0] I_15_0_1_1,
  input  [7:0] I_15_0_1_2,
  input  [7:0] I_15_0_2_0,
  input  [7:0] I_15_0_2_1,
  input  [7:0] I_15_0_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_1_2_0,
  output [7:0] O_1_2_1,
  output [7:0] O_1_2_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_2_1_2,
  output [7:0] O_2_2_0,
  output [7:0] O_2_2_1,
  output [7:0] O_2_2_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_3_1_2,
  output [7:0] O_3_2_0,
  output [7:0] O_3_2_1,
  output [7:0] O_3_2_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_4_1_2,
  output [7:0] O_4_2_0,
  output [7:0] O_4_2_1,
  output [7:0] O_4_2_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_5_1_2,
  output [7:0] O_5_2_0,
  output [7:0] O_5_2_1,
  output [7:0] O_5_2_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_6_1_2,
  output [7:0] O_6_2_0,
  output [7:0] O_6_2_1,
  output [7:0] O_6_2_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_7_1_2,
  output [7:0] O_7_2_0,
  output [7:0] O_7_2_1,
  output [7:0] O_7_2_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_8_1_0,
  output [7:0] O_8_1_1,
  output [7:0] O_8_1_2,
  output [7:0] O_8_2_0,
  output [7:0] O_8_2_1,
  output [7:0] O_8_2_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_9_1_0,
  output [7:0] O_9_1_1,
  output [7:0] O_9_1_2,
  output [7:0] O_9_2_0,
  output [7:0] O_9_2_1,
  output [7:0] O_9_2_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_10_1_0,
  output [7:0] O_10_1_1,
  output [7:0] O_10_1_2,
  output [7:0] O_10_2_0,
  output [7:0] O_10_2_1,
  output [7:0] O_10_2_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_11_1_0,
  output [7:0] O_11_1_1,
  output [7:0] O_11_1_2,
  output [7:0] O_11_2_0,
  output [7:0] O_11_2_1,
  output [7:0] O_11_2_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_12_1_0,
  output [7:0] O_12_1_1,
  output [7:0] O_12_1_2,
  output [7:0] O_12_2_0,
  output [7:0] O_12_2_1,
  output [7:0] O_12_2_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_13_1_0,
  output [7:0] O_13_1_1,
  output [7:0] O_13_1_2,
  output [7:0] O_13_2_0,
  output [7:0] O_13_2_1,
  output [7:0] O_13_2_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_14_1_0,
  output [7:0] O_14_1_1,
  output [7:0] O_14_1_2,
  output [7:0] O_14_2_0,
  output [7:0] O_14_2_1,
  output [7:0] O_14_2_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2,
  output [7:0] O_15_1_0,
  output [7:0] O_15_1_1,
  output [7:0] O_15_1_2,
  output [7:0] O_15_2_0,
  output [7:0] O_15_2_1,
  output [7:0] O_15_2_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_2_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Remove1S_3 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0_0(fst_op_I_0_0_0),
    .I_0_0_1(fst_op_I_0_0_1),
    .I_0_0_2(fst_op_I_0_0_2),
    .I_0_1_0(fst_op_I_0_1_0),
    .I_0_1_1(fst_op_I_0_1_1),
    .I_0_1_2(fst_op_I_0_1_2),
    .I_0_2_0(fst_op_I_0_2_0),
    .I_0_2_1(fst_op_I_0_2_1),
    .I_0_2_2(fst_op_I_0_2_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  Remove1S_3 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0_0(other_ops_0_I_0_0_0),
    .I_0_0_1(other_ops_0_I_0_0_1),
    .I_0_0_2(other_ops_0_I_0_0_2),
    .I_0_1_0(other_ops_0_I_0_1_0),
    .I_0_1_1(other_ops_0_I_0_1_1),
    .I_0_1_2(other_ops_0_I_0_1_2),
    .I_0_2_0(other_ops_0_I_0_2_0),
    .I_0_2_1(other_ops_0_I_0_2_1),
    .I_0_2_2(other_ops_0_I_0_2_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  Remove1S_3 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0_0(other_ops_1_I_0_0_0),
    .I_0_0_1(other_ops_1_I_0_0_1),
    .I_0_0_2(other_ops_1_I_0_0_2),
    .I_0_1_0(other_ops_1_I_0_1_0),
    .I_0_1_1(other_ops_1_I_0_1_1),
    .I_0_1_2(other_ops_1_I_0_1_2),
    .I_0_2_0(other_ops_1_I_0_2_0),
    .I_0_2_1(other_ops_1_I_0_2_1),
    .I_0_2_2(other_ops_1_I_0_2_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  Remove1S_3 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0_0(other_ops_2_I_0_0_0),
    .I_0_0_1(other_ops_2_I_0_0_1),
    .I_0_0_2(other_ops_2_I_0_0_2),
    .I_0_1_0(other_ops_2_I_0_1_0),
    .I_0_1_1(other_ops_2_I_0_1_1),
    .I_0_1_2(other_ops_2_I_0_1_2),
    .I_0_2_0(other_ops_2_I_0_2_0),
    .I_0_2_1(other_ops_2_I_0_2_1),
    .I_0_2_2(other_ops_2_I_0_2_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  Remove1S_3 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0_0(other_ops_3_I_0_0_0),
    .I_0_0_1(other_ops_3_I_0_0_1),
    .I_0_0_2(other_ops_3_I_0_0_2),
    .I_0_1_0(other_ops_3_I_0_1_0),
    .I_0_1_1(other_ops_3_I_0_1_1),
    .I_0_1_2(other_ops_3_I_0_1_2),
    .I_0_2_0(other_ops_3_I_0_2_0),
    .I_0_2_1(other_ops_3_I_0_2_1),
    .I_0_2_2(other_ops_3_I_0_2_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2),
    .O_2_0(other_ops_3_O_2_0),
    .O_2_1(other_ops_3_O_2_1),
    .O_2_2(other_ops_3_O_2_2)
  );
  Remove1S_3 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0_0(other_ops_4_I_0_0_0),
    .I_0_0_1(other_ops_4_I_0_0_1),
    .I_0_0_2(other_ops_4_I_0_0_2),
    .I_0_1_0(other_ops_4_I_0_1_0),
    .I_0_1_1(other_ops_4_I_0_1_1),
    .I_0_1_2(other_ops_4_I_0_1_2),
    .I_0_2_0(other_ops_4_I_0_2_0),
    .I_0_2_1(other_ops_4_I_0_2_1),
    .I_0_2_2(other_ops_4_I_0_2_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2),
    .O_2_0(other_ops_4_O_2_0),
    .O_2_1(other_ops_4_O_2_1),
    .O_2_2(other_ops_4_O_2_2)
  );
  Remove1S_3 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0_0(other_ops_5_I_0_0_0),
    .I_0_0_1(other_ops_5_I_0_0_1),
    .I_0_0_2(other_ops_5_I_0_0_2),
    .I_0_1_0(other_ops_5_I_0_1_0),
    .I_0_1_1(other_ops_5_I_0_1_1),
    .I_0_1_2(other_ops_5_I_0_1_2),
    .I_0_2_0(other_ops_5_I_0_2_0),
    .I_0_2_1(other_ops_5_I_0_2_1),
    .I_0_2_2(other_ops_5_I_0_2_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2),
    .O_2_0(other_ops_5_O_2_0),
    .O_2_1(other_ops_5_O_2_1),
    .O_2_2(other_ops_5_O_2_2)
  );
  Remove1S_3 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0_0(other_ops_6_I_0_0_0),
    .I_0_0_1(other_ops_6_I_0_0_1),
    .I_0_0_2(other_ops_6_I_0_0_2),
    .I_0_1_0(other_ops_6_I_0_1_0),
    .I_0_1_1(other_ops_6_I_0_1_1),
    .I_0_1_2(other_ops_6_I_0_1_2),
    .I_0_2_0(other_ops_6_I_0_2_0),
    .I_0_2_1(other_ops_6_I_0_2_1),
    .I_0_2_2(other_ops_6_I_0_2_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2),
    .O_2_0(other_ops_6_O_2_0),
    .O_2_1(other_ops_6_O_2_1),
    .O_2_2(other_ops_6_O_2_2)
  );
  Remove1S_3 other_ops_7 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0_0(other_ops_7_I_0_0_0),
    .I_0_0_1(other_ops_7_I_0_0_1),
    .I_0_0_2(other_ops_7_I_0_0_2),
    .I_0_1_0(other_ops_7_I_0_1_0),
    .I_0_1_1(other_ops_7_I_0_1_1),
    .I_0_1_2(other_ops_7_I_0_1_2),
    .I_0_2_0(other_ops_7_I_0_2_0),
    .I_0_2_1(other_ops_7_I_0_2_1),
    .I_0_2_2(other_ops_7_I_0_2_2),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_0_2(other_ops_7_O_0_2),
    .O_1_0(other_ops_7_O_1_0),
    .O_1_1(other_ops_7_O_1_1),
    .O_1_2(other_ops_7_O_1_2),
    .O_2_0(other_ops_7_O_2_0),
    .O_2_1(other_ops_7_O_2_1),
    .O_2_2(other_ops_7_O_2_2)
  );
  Remove1S_3 other_ops_8 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0_0(other_ops_8_I_0_0_0),
    .I_0_0_1(other_ops_8_I_0_0_1),
    .I_0_0_2(other_ops_8_I_0_0_2),
    .I_0_1_0(other_ops_8_I_0_1_0),
    .I_0_1_1(other_ops_8_I_0_1_1),
    .I_0_1_2(other_ops_8_I_0_1_2),
    .I_0_2_0(other_ops_8_I_0_2_0),
    .I_0_2_1(other_ops_8_I_0_2_1),
    .I_0_2_2(other_ops_8_I_0_2_2),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_0_2(other_ops_8_O_0_2),
    .O_1_0(other_ops_8_O_1_0),
    .O_1_1(other_ops_8_O_1_1),
    .O_1_2(other_ops_8_O_1_2),
    .O_2_0(other_ops_8_O_2_0),
    .O_2_1(other_ops_8_O_2_1),
    .O_2_2(other_ops_8_O_2_2)
  );
  Remove1S_3 other_ops_9 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0_0(other_ops_9_I_0_0_0),
    .I_0_0_1(other_ops_9_I_0_0_1),
    .I_0_0_2(other_ops_9_I_0_0_2),
    .I_0_1_0(other_ops_9_I_0_1_0),
    .I_0_1_1(other_ops_9_I_0_1_1),
    .I_0_1_2(other_ops_9_I_0_1_2),
    .I_0_2_0(other_ops_9_I_0_2_0),
    .I_0_2_1(other_ops_9_I_0_2_1),
    .I_0_2_2(other_ops_9_I_0_2_2),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_0_2(other_ops_9_O_0_2),
    .O_1_0(other_ops_9_O_1_0),
    .O_1_1(other_ops_9_O_1_1),
    .O_1_2(other_ops_9_O_1_2),
    .O_2_0(other_ops_9_O_2_0),
    .O_2_1(other_ops_9_O_2_1),
    .O_2_2(other_ops_9_O_2_2)
  );
  Remove1S_3 other_ops_10 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0_0(other_ops_10_I_0_0_0),
    .I_0_0_1(other_ops_10_I_0_0_1),
    .I_0_0_2(other_ops_10_I_0_0_2),
    .I_0_1_0(other_ops_10_I_0_1_0),
    .I_0_1_1(other_ops_10_I_0_1_1),
    .I_0_1_2(other_ops_10_I_0_1_2),
    .I_0_2_0(other_ops_10_I_0_2_0),
    .I_0_2_1(other_ops_10_I_0_2_1),
    .I_0_2_2(other_ops_10_I_0_2_2),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_0_2(other_ops_10_O_0_2),
    .O_1_0(other_ops_10_O_1_0),
    .O_1_1(other_ops_10_O_1_1),
    .O_1_2(other_ops_10_O_1_2),
    .O_2_0(other_ops_10_O_2_0),
    .O_2_1(other_ops_10_O_2_1),
    .O_2_2(other_ops_10_O_2_2)
  );
  Remove1S_3 other_ops_11 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0_0(other_ops_11_I_0_0_0),
    .I_0_0_1(other_ops_11_I_0_0_1),
    .I_0_0_2(other_ops_11_I_0_0_2),
    .I_0_1_0(other_ops_11_I_0_1_0),
    .I_0_1_1(other_ops_11_I_0_1_1),
    .I_0_1_2(other_ops_11_I_0_1_2),
    .I_0_2_0(other_ops_11_I_0_2_0),
    .I_0_2_1(other_ops_11_I_0_2_1),
    .I_0_2_2(other_ops_11_I_0_2_2),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_0_2(other_ops_11_O_0_2),
    .O_1_0(other_ops_11_O_1_0),
    .O_1_1(other_ops_11_O_1_1),
    .O_1_2(other_ops_11_O_1_2),
    .O_2_0(other_ops_11_O_2_0),
    .O_2_1(other_ops_11_O_2_1),
    .O_2_2(other_ops_11_O_2_2)
  );
  Remove1S_3 other_ops_12 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0_0(other_ops_12_I_0_0_0),
    .I_0_0_1(other_ops_12_I_0_0_1),
    .I_0_0_2(other_ops_12_I_0_0_2),
    .I_0_1_0(other_ops_12_I_0_1_0),
    .I_0_1_1(other_ops_12_I_0_1_1),
    .I_0_1_2(other_ops_12_I_0_1_2),
    .I_0_2_0(other_ops_12_I_0_2_0),
    .I_0_2_1(other_ops_12_I_0_2_1),
    .I_0_2_2(other_ops_12_I_0_2_2),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_0_2(other_ops_12_O_0_2),
    .O_1_0(other_ops_12_O_1_0),
    .O_1_1(other_ops_12_O_1_1),
    .O_1_2(other_ops_12_O_1_2),
    .O_2_0(other_ops_12_O_2_0),
    .O_2_1(other_ops_12_O_2_1),
    .O_2_2(other_ops_12_O_2_2)
  );
  Remove1S_3 other_ops_13 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0_0(other_ops_13_I_0_0_0),
    .I_0_0_1(other_ops_13_I_0_0_1),
    .I_0_0_2(other_ops_13_I_0_0_2),
    .I_0_1_0(other_ops_13_I_0_1_0),
    .I_0_1_1(other_ops_13_I_0_1_1),
    .I_0_1_2(other_ops_13_I_0_1_2),
    .I_0_2_0(other_ops_13_I_0_2_0),
    .I_0_2_1(other_ops_13_I_0_2_1),
    .I_0_2_2(other_ops_13_I_0_2_2),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_0_2(other_ops_13_O_0_2),
    .O_1_0(other_ops_13_O_1_0),
    .O_1_1(other_ops_13_O_1_1),
    .O_1_2(other_ops_13_O_1_2),
    .O_2_0(other_ops_13_O_2_0),
    .O_2_1(other_ops_13_O_2_1),
    .O_2_2(other_ops_13_O_2_2)
  );
  Remove1S_3 other_ops_14 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0_0(other_ops_14_I_0_0_0),
    .I_0_0_1(other_ops_14_I_0_0_1),
    .I_0_0_2(other_ops_14_I_0_0_2),
    .I_0_1_0(other_ops_14_I_0_1_0),
    .I_0_1_1(other_ops_14_I_0_1_1),
    .I_0_1_2(other_ops_14_I_0_1_2),
    .I_0_2_0(other_ops_14_I_0_2_0),
    .I_0_2_1(other_ops_14_I_0_2_1),
    .I_0_2_2(other_ops_14_I_0_2_2),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_0_2(other_ops_14_O_0_2),
    .O_1_0(other_ops_14_O_1_0),
    .O_1_1(other_ops_14_O_1_1),
    .O_1_2(other_ops_14_O_1_2),
    .O_2_0(other_ops_14_O_2_0),
    .O_2_1(other_ops_14_O_2_1),
    .O_2_2(other_ops_14_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[MapS.scala 17:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[MapS.scala 17:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[MapS.scala 17:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[MapS.scala 17:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[MapS.scala 17:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[MapS.scala 17:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[MapS.scala 17:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[MapS.scala 21:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[MapS.scala 21:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[MapS.scala 21:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[MapS.scala 21:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[MapS.scala 21:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[MapS.scala 21:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[MapS.scala 21:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[MapS.scala 21:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[MapS.scala 21:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[MapS.scala 21:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[MapS.scala 21:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[MapS.scala 21:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[MapS.scala 21:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[MapS.scala 21:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[MapS.scala 21:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[MapS.scala 21:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[MapS.scala 21:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[MapS.scala 21:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[MapS.scala 21:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[MapS.scala 21:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[MapS.scala 21:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[MapS.scala 21:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[MapS.scala 21:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[MapS.scala 21:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[MapS.scala 21:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[MapS.scala 21:12]
  assign O_4_2_0 = other_ops_3_O_2_0; // @[MapS.scala 21:12]
  assign O_4_2_1 = other_ops_3_O_2_1; // @[MapS.scala 21:12]
  assign O_4_2_2 = other_ops_3_O_2_2; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[MapS.scala 21:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[MapS.scala 21:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[MapS.scala 21:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[MapS.scala 21:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[MapS.scala 21:12]
  assign O_5_2_0 = other_ops_4_O_2_0; // @[MapS.scala 21:12]
  assign O_5_2_1 = other_ops_4_O_2_1; // @[MapS.scala 21:12]
  assign O_5_2_2 = other_ops_4_O_2_2; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[MapS.scala 21:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[MapS.scala 21:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[MapS.scala 21:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[MapS.scala 21:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[MapS.scala 21:12]
  assign O_6_2_0 = other_ops_5_O_2_0; // @[MapS.scala 21:12]
  assign O_6_2_1 = other_ops_5_O_2_1; // @[MapS.scala 21:12]
  assign O_6_2_2 = other_ops_5_O_2_2; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[MapS.scala 21:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[MapS.scala 21:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[MapS.scala 21:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[MapS.scala 21:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[MapS.scala 21:12]
  assign O_7_2_0 = other_ops_6_O_2_0; // @[MapS.scala 21:12]
  assign O_7_2_1 = other_ops_6_O_2_1; // @[MapS.scala 21:12]
  assign O_7_2_2 = other_ops_6_O_2_2; // @[MapS.scala 21:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[MapS.scala 21:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[MapS.scala 21:12]
  assign O_8_0_2 = other_ops_7_O_0_2; // @[MapS.scala 21:12]
  assign O_8_1_0 = other_ops_7_O_1_0; // @[MapS.scala 21:12]
  assign O_8_1_1 = other_ops_7_O_1_1; // @[MapS.scala 21:12]
  assign O_8_1_2 = other_ops_7_O_1_2; // @[MapS.scala 21:12]
  assign O_8_2_0 = other_ops_7_O_2_0; // @[MapS.scala 21:12]
  assign O_8_2_1 = other_ops_7_O_2_1; // @[MapS.scala 21:12]
  assign O_8_2_2 = other_ops_7_O_2_2; // @[MapS.scala 21:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[MapS.scala 21:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[MapS.scala 21:12]
  assign O_9_0_2 = other_ops_8_O_0_2; // @[MapS.scala 21:12]
  assign O_9_1_0 = other_ops_8_O_1_0; // @[MapS.scala 21:12]
  assign O_9_1_1 = other_ops_8_O_1_1; // @[MapS.scala 21:12]
  assign O_9_1_2 = other_ops_8_O_1_2; // @[MapS.scala 21:12]
  assign O_9_2_0 = other_ops_8_O_2_0; // @[MapS.scala 21:12]
  assign O_9_2_1 = other_ops_8_O_2_1; // @[MapS.scala 21:12]
  assign O_9_2_2 = other_ops_8_O_2_2; // @[MapS.scala 21:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[MapS.scala 21:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[MapS.scala 21:12]
  assign O_10_0_2 = other_ops_9_O_0_2; // @[MapS.scala 21:12]
  assign O_10_1_0 = other_ops_9_O_1_0; // @[MapS.scala 21:12]
  assign O_10_1_1 = other_ops_9_O_1_1; // @[MapS.scala 21:12]
  assign O_10_1_2 = other_ops_9_O_1_2; // @[MapS.scala 21:12]
  assign O_10_2_0 = other_ops_9_O_2_0; // @[MapS.scala 21:12]
  assign O_10_2_1 = other_ops_9_O_2_1; // @[MapS.scala 21:12]
  assign O_10_2_2 = other_ops_9_O_2_2; // @[MapS.scala 21:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[MapS.scala 21:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[MapS.scala 21:12]
  assign O_11_0_2 = other_ops_10_O_0_2; // @[MapS.scala 21:12]
  assign O_11_1_0 = other_ops_10_O_1_0; // @[MapS.scala 21:12]
  assign O_11_1_1 = other_ops_10_O_1_1; // @[MapS.scala 21:12]
  assign O_11_1_2 = other_ops_10_O_1_2; // @[MapS.scala 21:12]
  assign O_11_2_0 = other_ops_10_O_2_0; // @[MapS.scala 21:12]
  assign O_11_2_1 = other_ops_10_O_2_1; // @[MapS.scala 21:12]
  assign O_11_2_2 = other_ops_10_O_2_2; // @[MapS.scala 21:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[MapS.scala 21:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[MapS.scala 21:12]
  assign O_12_0_2 = other_ops_11_O_0_2; // @[MapS.scala 21:12]
  assign O_12_1_0 = other_ops_11_O_1_0; // @[MapS.scala 21:12]
  assign O_12_1_1 = other_ops_11_O_1_1; // @[MapS.scala 21:12]
  assign O_12_1_2 = other_ops_11_O_1_2; // @[MapS.scala 21:12]
  assign O_12_2_0 = other_ops_11_O_2_0; // @[MapS.scala 21:12]
  assign O_12_2_1 = other_ops_11_O_2_1; // @[MapS.scala 21:12]
  assign O_12_2_2 = other_ops_11_O_2_2; // @[MapS.scala 21:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[MapS.scala 21:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[MapS.scala 21:12]
  assign O_13_0_2 = other_ops_12_O_0_2; // @[MapS.scala 21:12]
  assign O_13_1_0 = other_ops_12_O_1_0; // @[MapS.scala 21:12]
  assign O_13_1_1 = other_ops_12_O_1_1; // @[MapS.scala 21:12]
  assign O_13_1_2 = other_ops_12_O_1_2; // @[MapS.scala 21:12]
  assign O_13_2_0 = other_ops_12_O_2_0; // @[MapS.scala 21:12]
  assign O_13_2_1 = other_ops_12_O_2_1; // @[MapS.scala 21:12]
  assign O_13_2_2 = other_ops_12_O_2_2; // @[MapS.scala 21:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[MapS.scala 21:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[MapS.scala 21:12]
  assign O_14_0_2 = other_ops_13_O_0_2; // @[MapS.scala 21:12]
  assign O_14_1_0 = other_ops_13_O_1_0; // @[MapS.scala 21:12]
  assign O_14_1_1 = other_ops_13_O_1_1; // @[MapS.scala 21:12]
  assign O_14_1_2 = other_ops_13_O_1_2; // @[MapS.scala 21:12]
  assign O_14_2_0 = other_ops_13_O_2_0; // @[MapS.scala 21:12]
  assign O_14_2_1 = other_ops_13_O_2_1; // @[MapS.scala 21:12]
  assign O_14_2_2 = other_ops_13_O_2_2; // @[MapS.scala 21:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[MapS.scala 21:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[MapS.scala 21:12]
  assign O_15_0_2 = other_ops_14_O_0_2; // @[MapS.scala 21:12]
  assign O_15_1_0 = other_ops_14_O_1_0; // @[MapS.scala 21:12]
  assign O_15_1_1 = other_ops_14_O_1_1; // @[MapS.scala 21:12]
  assign O_15_1_2 = other_ops_14_O_1_2; // @[MapS.scala 21:12]
  assign O_15_2_0 = other_ops_14_O_2_0; // @[MapS.scala 21:12]
  assign O_15_2_1 = other_ops_14_O_2_1; // @[MapS.scala 21:12]
  assign O_15_2_2 = other_ops_14_O_2_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0_0 = I_0_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_1 = I_0_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_2 = I_0_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_0 = I_0_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_1 = I_0_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_2 = I_0_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_0 = I_0_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_1 = I_0_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_2 = I_0_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0_0 = I_1_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_1 = I_1_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_2 = I_1_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_0 = I_1_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_1 = I_1_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_2 = I_1_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_0 = I_1_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_1 = I_1_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_2 = I_1_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0_0 = I_2_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_1 = I_2_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_2 = I_2_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_0 = I_2_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_1 = I_2_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_2 = I_2_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_0 = I_2_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_1 = I_2_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_2 = I_2_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0_0 = I_3_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_1 = I_3_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_2 = I_3_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_0 = I_3_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_1 = I_3_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_2 = I_3_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_0 = I_3_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_1 = I_3_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_2 = I_3_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0_0 = I_4_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_1 = I_4_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_2 = I_4_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_0 = I_4_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_1 = I_4_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_2 = I_4_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_0 = I_4_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_1 = I_4_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_2 = I_4_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0_0 = I_5_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_1 = I_5_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_2 = I_5_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_0 = I_5_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_1 = I_5_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_2 = I_5_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_0 = I_5_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_1 = I_5_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_2 = I_5_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0_0 = I_6_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_1 = I_6_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_2 = I_6_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_0 = I_6_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_1 = I_6_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_2 = I_6_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_0 = I_6_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_1 = I_6_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_2 = I_6_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0_0 = I_7_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_1 = I_7_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_2 = I_7_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_0 = I_7_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_1 = I_7_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_2 = I_7_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_0 = I_7_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_1 = I_7_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_2 = I_7_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0_0 = I_8_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_0_1 = I_8_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_0_2 = I_8_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_0 = I_8_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_1 = I_8_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_2 = I_8_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2_0 = I_8_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2_1 = I_8_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2_2 = I_8_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0_0 = I_9_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_0_1 = I_9_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_0_2 = I_9_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_0 = I_9_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_1 = I_9_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_2 = I_9_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2_0 = I_9_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2_1 = I_9_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2_2 = I_9_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0_0 = I_10_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_0_1 = I_10_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_0_2 = I_10_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_0 = I_10_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_1 = I_10_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_2 = I_10_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2_0 = I_10_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2_1 = I_10_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2_2 = I_10_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0_0 = I_11_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_0_1 = I_11_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_0_2 = I_11_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_0 = I_11_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_1 = I_11_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_2 = I_11_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2_0 = I_11_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2_1 = I_11_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2_2 = I_11_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0_0 = I_12_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_0_1 = I_12_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_0_2 = I_12_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_0 = I_12_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_1 = I_12_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_2 = I_12_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2_0 = I_12_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2_1 = I_12_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2_2 = I_12_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0_0 = I_13_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_0_1 = I_13_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_0_2 = I_13_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_0 = I_13_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_1 = I_13_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_2 = I_13_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2_0 = I_13_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2_1 = I_13_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2_2 = I_13_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0_0 = I_14_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_0_1 = I_14_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_0_2 = I_14_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_0 = I_14_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_1 = I_14_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_2 = I_14_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2_0 = I_14_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2_1 = I_14_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2_2 = I_14_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0_0 = I_15_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_0_1 = I_15_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_0_2 = I_15_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_0 = I_15_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_1 = I_15_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_2 = I_15_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2_0 = I_15_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2_1 = I_15_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2_2 = I_15_0_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0_0,
  input  [7:0] I_0_0_0_1,
  input  [7:0] I_0_0_0_2,
  input  [7:0] I_0_0_1_0,
  input  [7:0] I_0_0_1_1,
  input  [7:0] I_0_0_1_2,
  input  [7:0] I_0_0_2_0,
  input  [7:0] I_0_0_2_1,
  input  [7:0] I_0_0_2_2,
  input  [7:0] I_1_0_0_0,
  input  [7:0] I_1_0_0_1,
  input  [7:0] I_1_0_0_2,
  input  [7:0] I_1_0_1_0,
  input  [7:0] I_1_0_1_1,
  input  [7:0] I_1_0_1_2,
  input  [7:0] I_1_0_2_0,
  input  [7:0] I_1_0_2_1,
  input  [7:0] I_1_0_2_2,
  input  [7:0] I_2_0_0_0,
  input  [7:0] I_2_0_0_1,
  input  [7:0] I_2_0_0_2,
  input  [7:0] I_2_0_1_0,
  input  [7:0] I_2_0_1_1,
  input  [7:0] I_2_0_1_2,
  input  [7:0] I_2_0_2_0,
  input  [7:0] I_2_0_2_1,
  input  [7:0] I_2_0_2_2,
  input  [7:0] I_3_0_0_0,
  input  [7:0] I_3_0_0_1,
  input  [7:0] I_3_0_0_2,
  input  [7:0] I_3_0_1_0,
  input  [7:0] I_3_0_1_1,
  input  [7:0] I_3_0_1_2,
  input  [7:0] I_3_0_2_0,
  input  [7:0] I_3_0_2_1,
  input  [7:0] I_3_0_2_2,
  input  [7:0] I_4_0_0_0,
  input  [7:0] I_4_0_0_1,
  input  [7:0] I_4_0_0_2,
  input  [7:0] I_4_0_1_0,
  input  [7:0] I_4_0_1_1,
  input  [7:0] I_4_0_1_2,
  input  [7:0] I_4_0_2_0,
  input  [7:0] I_4_0_2_1,
  input  [7:0] I_4_0_2_2,
  input  [7:0] I_5_0_0_0,
  input  [7:0] I_5_0_0_1,
  input  [7:0] I_5_0_0_2,
  input  [7:0] I_5_0_1_0,
  input  [7:0] I_5_0_1_1,
  input  [7:0] I_5_0_1_2,
  input  [7:0] I_5_0_2_0,
  input  [7:0] I_5_0_2_1,
  input  [7:0] I_5_0_2_2,
  input  [7:0] I_6_0_0_0,
  input  [7:0] I_6_0_0_1,
  input  [7:0] I_6_0_0_2,
  input  [7:0] I_6_0_1_0,
  input  [7:0] I_6_0_1_1,
  input  [7:0] I_6_0_1_2,
  input  [7:0] I_6_0_2_0,
  input  [7:0] I_6_0_2_1,
  input  [7:0] I_6_0_2_2,
  input  [7:0] I_7_0_0_0,
  input  [7:0] I_7_0_0_1,
  input  [7:0] I_7_0_0_2,
  input  [7:0] I_7_0_1_0,
  input  [7:0] I_7_0_1_1,
  input  [7:0] I_7_0_1_2,
  input  [7:0] I_7_0_2_0,
  input  [7:0] I_7_0_2_1,
  input  [7:0] I_7_0_2_2,
  input  [7:0] I_8_0_0_0,
  input  [7:0] I_8_0_0_1,
  input  [7:0] I_8_0_0_2,
  input  [7:0] I_8_0_1_0,
  input  [7:0] I_8_0_1_1,
  input  [7:0] I_8_0_1_2,
  input  [7:0] I_8_0_2_0,
  input  [7:0] I_8_0_2_1,
  input  [7:0] I_8_0_2_2,
  input  [7:0] I_9_0_0_0,
  input  [7:0] I_9_0_0_1,
  input  [7:0] I_9_0_0_2,
  input  [7:0] I_9_0_1_0,
  input  [7:0] I_9_0_1_1,
  input  [7:0] I_9_0_1_2,
  input  [7:0] I_9_0_2_0,
  input  [7:0] I_9_0_2_1,
  input  [7:0] I_9_0_2_2,
  input  [7:0] I_10_0_0_0,
  input  [7:0] I_10_0_0_1,
  input  [7:0] I_10_0_0_2,
  input  [7:0] I_10_0_1_0,
  input  [7:0] I_10_0_1_1,
  input  [7:0] I_10_0_1_2,
  input  [7:0] I_10_0_2_0,
  input  [7:0] I_10_0_2_1,
  input  [7:0] I_10_0_2_2,
  input  [7:0] I_11_0_0_0,
  input  [7:0] I_11_0_0_1,
  input  [7:0] I_11_0_0_2,
  input  [7:0] I_11_0_1_0,
  input  [7:0] I_11_0_1_1,
  input  [7:0] I_11_0_1_2,
  input  [7:0] I_11_0_2_0,
  input  [7:0] I_11_0_2_1,
  input  [7:0] I_11_0_2_2,
  input  [7:0] I_12_0_0_0,
  input  [7:0] I_12_0_0_1,
  input  [7:0] I_12_0_0_2,
  input  [7:0] I_12_0_1_0,
  input  [7:0] I_12_0_1_1,
  input  [7:0] I_12_0_1_2,
  input  [7:0] I_12_0_2_0,
  input  [7:0] I_12_0_2_1,
  input  [7:0] I_12_0_2_2,
  input  [7:0] I_13_0_0_0,
  input  [7:0] I_13_0_0_1,
  input  [7:0] I_13_0_0_2,
  input  [7:0] I_13_0_1_0,
  input  [7:0] I_13_0_1_1,
  input  [7:0] I_13_0_1_2,
  input  [7:0] I_13_0_2_0,
  input  [7:0] I_13_0_2_1,
  input  [7:0] I_13_0_2_2,
  input  [7:0] I_14_0_0_0,
  input  [7:0] I_14_0_0_1,
  input  [7:0] I_14_0_0_2,
  input  [7:0] I_14_0_1_0,
  input  [7:0] I_14_0_1_1,
  input  [7:0] I_14_0_1_2,
  input  [7:0] I_14_0_2_0,
  input  [7:0] I_14_0_2_1,
  input  [7:0] I_14_0_2_2,
  input  [7:0] I_15_0_0_0,
  input  [7:0] I_15_0_0_1,
  input  [7:0] I_15_0_0_2,
  input  [7:0] I_15_0_1_0,
  input  [7:0] I_15_0_1_1,
  input  [7:0] I_15_0_1_2,
  input  [7:0] I_15_0_2_0,
  input  [7:0] I_15_0_2_1,
  input  [7:0] I_15_0_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_1_2_0,
  output [7:0] O_1_2_1,
  output [7:0] O_1_2_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_2_1_2,
  output [7:0] O_2_2_0,
  output [7:0] O_2_2_1,
  output [7:0] O_2_2_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_3_1_2,
  output [7:0] O_3_2_0,
  output [7:0] O_3_2_1,
  output [7:0] O_3_2_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_4_1_2,
  output [7:0] O_4_2_0,
  output [7:0] O_4_2_1,
  output [7:0] O_4_2_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_5_1_2,
  output [7:0] O_5_2_0,
  output [7:0] O_5_2_1,
  output [7:0] O_5_2_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_6_1_2,
  output [7:0] O_6_2_0,
  output [7:0] O_6_2_1,
  output [7:0] O_6_2_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_7_1_2,
  output [7:0] O_7_2_0,
  output [7:0] O_7_2_1,
  output [7:0] O_7_2_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_8_1_0,
  output [7:0] O_8_1_1,
  output [7:0] O_8_1_2,
  output [7:0] O_8_2_0,
  output [7:0] O_8_2_1,
  output [7:0] O_8_2_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_9_1_0,
  output [7:0] O_9_1_1,
  output [7:0] O_9_1_2,
  output [7:0] O_9_2_0,
  output [7:0] O_9_2_1,
  output [7:0] O_9_2_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_10_1_0,
  output [7:0] O_10_1_1,
  output [7:0] O_10_1_2,
  output [7:0] O_10_2_0,
  output [7:0] O_10_2_1,
  output [7:0] O_10_2_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_11_1_0,
  output [7:0] O_11_1_1,
  output [7:0] O_11_1_2,
  output [7:0] O_11_2_0,
  output [7:0] O_11_2_1,
  output [7:0] O_11_2_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_12_1_0,
  output [7:0] O_12_1_1,
  output [7:0] O_12_1_2,
  output [7:0] O_12_2_0,
  output [7:0] O_12_2_1,
  output [7:0] O_12_2_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_13_1_0,
  output [7:0] O_13_1_1,
  output [7:0] O_13_1_2,
  output [7:0] O_13_2_0,
  output [7:0] O_13_2_1,
  output [7:0] O_13_2_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_14_1_0,
  output [7:0] O_14_1_1,
  output [7:0] O_14_1_2,
  output [7:0] O_14_2_0,
  output [7:0] O_14_2_1,
  output [7:0] O_14_2_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2,
  output [7:0] O_15_1_0,
  output [7:0] O_15_1_1,
  output [7:0] O_15_1_2,
  output [7:0] O_15_2_0,
  output [7:0] O_15_2_1,
  output [7:0] O_15_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_2_2; // @[MapT.scala 8:20]
  MapS_6 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0_0(op_I_0_0_0_0),
    .I_0_0_0_1(op_I_0_0_0_1),
    .I_0_0_0_2(op_I_0_0_0_2),
    .I_0_0_1_0(op_I_0_0_1_0),
    .I_0_0_1_1(op_I_0_0_1_1),
    .I_0_0_1_2(op_I_0_0_1_2),
    .I_0_0_2_0(op_I_0_0_2_0),
    .I_0_0_2_1(op_I_0_0_2_1),
    .I_0_0_2_2(op_I_0_0_2_2),
    .I_1_0_0_0(op_I_1_0_0_0),
    .I_1_0_0_1(op_I_1_0_0_1),
    .I_1_0_0_2(op_I_1_0_0_2),
    .I_1_0_1_0(op_I_1_0_1_0),
    .I_1_0_1_1(op_I_1_0_1_1),
    .I_1_0_1_2(op_I_1_0_1_2),
    .I_1_0_2_0(op_I_1_0_2_0),
    .I_1_0_2_1(op_I_1_0_2_1),
    .I_1_0_2_2(op_I_1_0_2_2),
    .I_2_0_0_0(op_I_2_0_0_0),
    .I_2_0_0_1(op_I_2_0_0_1),
    .I_2_0_0_2(op_I_2_0_0_2),
    .I_2_0_1_0(op_I_2_0_1_0),
    .I_2_0_1_1(op_I_2_0_1_1),
    .I_2_0_1_2(op_I_2_0_1_2),
    .I_2_0_2_0(op_I_2_0_2_0),
    .I_2_0_2_1(op_I_2_0_2_1),
    .I_2_0_2_2(op_I_2_0_2_2),
    .I_3_0_0_0(op_I_3_0_0_0),
    .I_3_0_0_1(op_I_3_0_0_1),
    .I_3_0_0_2(op_I_3_0_0_2),
    .I_3_0_1_0(op_I_3_0_1_0),
    .I_3_0_1_1(op_I_3_0_1_1),
    .I_3_0_1_2(op_I_3_0_1_2),
    .I_3_0_2_0(op_I_3_0_2_0),
    .I_3_0_2_1(op_I_3_0_2_1),
    .I_3_0_2_2(op_I_3_0_2_2),
    .I_4_0_0_0(op_I_4_0_0_0),
    .I_4_0_0_1(op_I_4_0_0_1),
    .I_4_0_0_2(op_I_4_0_0_2),
    .I_4_0_1_0(op_I_4_0_1_0),
    .I_4_0_1_1(op_I_4_0_1_1),
    .I_4_0_1_2(op_I_4_0_1_2),
    .I_4_0_2_0(op_I_4_0_2_0),
    .I_4_0_2_1(op_I_4_0_2_1),
    .I_4_0_2_2(op_I_4_0_2_2),
    .I_5_0_0_0(op_I_5_0_0_0),
    .I_5_0_0_1(op_I_5_0_0_1),
    .I_5_0_0_2(op_I_5_0_0_2),
    .I_5_0_1_0(op_I_5_0_1_0),
    .I_5_0_1_1(op_I_5_0_1_1),
    .I_5_0_1_2(op_I_5_0_1_2),
    .I_5_0_2_0(op_I_5_0_2_0),
    .I_5_0_2_1(op_I_5_0_2_1),
    .I_5_0_2_2(op_I_5_0_2_2),
    .I_6_0_0_0(op_I_6_0_0_0),
    .I_6_0_0_1(op_I_6_0_0_1),
    .I_6_0_0_2(op_I_6_0_0_2),
    .I_6_0_1_0(op_I_6_0_1_0),
    .I_6_0_1_1(op_I_6_0_1_1),
    .I_6_0_1_2(op_I_6_0_1_2),
    .I_6_0_2_0(op_I_6_0_2_0),
    .I_6_0_2_1(op_I_6_0_2_1),
    .I_6_0_2_2(op_I_6_0_2_2),
    .I_7_0_0_0(op_I_7_0_0_0),
    .I_7_0_0_1(op_I_7_0_0_1),
    .I_7_0_0_2(op_I_7_0_0_2),
    .I_7_0_1_0(op_I_7_0_1_0),
    .I_7_0_1_1(op_I_7_0_1_1),
    .I_7_0_1_2(op_I_7_0_1_2),
    .I_7_0_2_0(op_I_7_0_2_0),
    .I_7_0_2_1(op_I_7_0_2_1),
    .I_7_0_2_2(op_I_7_0_2_2),
    .I_8_0_0_0(op_I_8_0_0_0),
    .I_8_0_0_1(op_I_8_0_0_1),
    .I_8_0_0_2(op_I_8_0_0_2),
    .I_8_0_1_0(op_I_8_0_1_0),
    .I_8_0_1_1(op_I_8_0_1_1),
    .I_8_0_1_2(op_I_8_0_1_2),
    .I_8_0_2_0(op_I_8_0_2_0),
    .I_8_0_2_1(op_I_8_0_2_1),
    .I_8_0_2_2(op_I_8_0_2_2),
    .I_9_0_0_0(op_I_9_0_0_0),
    .I_9_0_0_1(op_I_9_0_0_1),
    .I_9_0_0_2(op_I_9_0_0_2),
    .I_9_0_1_0(op_I_9_0_1_0),
    .I_9_0_1_1(op_I_9_0_1_1),
    .I_9_0_1_2(op_I_9_0_1_2),
    .I_9_0_2_0(op_I_9_0_2_0),
    .I_9_0_2_1(op_I_9_0_2_1),
    .I_9_0_2_2(op_I_9_0_2_2),
    .I_10_0_0_0(op_I_10_0_0_0),
    .I_10_0_0_1(op_I_10_0_0_1),
    .I_10_0_0_2(op_I_10_0_0_2),
    .I_10_0_1_0(op_I_10_0_1_0),
    .I_10_0_1_1(op_I_10_0_1_1),
    .I_10_0_1_2(op_I_10_0_1_2),
    .I_10_0_2_0(op_I_10_0_2_0),
    .I_10_0_2_1(op_I_10_0_2_1),
    .I_10_0_2_2(op_I_10_0_2_2),
    .I_11_0_0_0(op_I_11_0_0_0),
    .I_11_0_0_1(op_I_11_0_0_1),
    .I_11_0_0_2(op_I_11_0_0_2),
    .I_11_0_1_0(op_I_11_0_1_0),
    .I_11_0_1_1(op_I_11_0_1_1),
    .I_11_0_1_2(op_I_11_0_1_2),
    .I_11_0_2_0(op_I_11_0_2_0),
    .I_11_0_2_1(op_I_11_0_2_1),
    .I_11_0_2_2(op_I_11_0_2_2),
    .I_12_0_0_0(op_I_12_0_0_0),
    .I_12_0_0_1(op_I_12_0_0_1),
    .I_12_0_0_2(op_I_12_0_0_2),
    .I_12_0_1_0(op_I_12_0_1_0),
    .I_12_0_1_1(op_I_12_0_1_1),
    .I_12_0_1_2(op_I_12_0_1_2),
    .I_12_0_2_0(op_I_12_0_2_0),
    .I_12_0_2_1(op_I_12_0_2_1),
    .I_12_0_2_2(op_I_12_0_2_2),
    .I_13_0_0_0(op_I_13_0_0_0),
    .I_13_0_0_1(op_I_13_0_0_1),
    .I_13_0_0_2(op_I_13_0_0_2),
    .I_13_0_1_0(op_I_13_0_1_0),
    .I_13_0_1_1(op_I_13_0_1_1),
    .I_13_0_1_2(op_I_13_0_1_2),
    .I_13_0_2_0(op_I_13_0_2_0),
    .I_13_0_2_1(op_I_13_0_2_1),
    .I_13_0_2_2(op_I_13_0_2_2),
    .I_14_0_0_0(op_I_14_0_0_0),
    .I_14_0_0_1(op_I_14_0_0_1),
    .I_14_0_0_2(op_I_14_0_0_2),
    .I_14_0_1_0(op_I_14_0_1_0),
    .I_14_0_1_1(op_I_14_0_1_1),
    .I_14_0_1_2(op_I_14_0_1_2),
    .I_14_0_2_0(op_I_14_0_2_0),
    .I_14_0_2_1(op_I_14_0_2_1),
    .I_14_0_2_2(op_I_14_0_2_2),
    .I_15_0_0_0(op_I_15_0_0_0),
    .I_15_0_0_1(op_I_15_0_0_1),
    .I_15_0_0_2(op_I_15_0_0_2),
    .I_15_0_1_0(op_I_15_0_1_0),
    .I_15_0_1_1(op_I_15_0_1_1),
    .I_15_0_1_2(op_I_15_0_1_2),
    .I_15_0_2_0(op_I_15_0_2_0),
    .I_15_0_2_1(op_I_15_0_2_1),
    .I_15_0_2_2(op_I_15_0_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_2_2_0(op_O_2_2_0),
    .O_2_2_1(op_O_2_2_1),
    .O_2_2_2(op_O_2_2_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_3_2_0(op_O_3_2_0),
    .O_3_2_1(op_O_3_2_1),
    .O_3_2_2(op_O_3_2_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_4_2_0(op_O_4_2_0),
    .O_4_2_1(op_O_4_2_1),
    .O_4_2_2(op_O_4_2_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_5_2_0(op_O_5_2_0),
    .O_5_2_1(op_O_5_2_1),
    .O_5_2_2(op_O_5_2_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_6_2_0(op_O_6_2_0),
    .O_6_2_1(op_O_6_2_1),
    .O_6_2_2(op_O_6_2_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2),
    .O_7_2_0(op_O_7_2_0),
    .O_7_2_1(op_O_7_2_1),
    .O_7_2_2(op_O_7_2_2),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_0_2(op_O_8_0_2),
    .O_8_1_0(op_O_8_1_0),
    .O_8_1_1(op_O_8_1_1),
    .O_8_1_2(op_O_8_1_2),
    .O_8_2_0(op_O_8_2_0),
    .O_8_2_1(op_O_8_2_1),
    .O_8_2_2(op_O_8_2_2),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_0_2(op_O_9_0_2),
    .O_9_1_0(op_O_9_1_0),
    .O_9_1_1(op_O_9_1_1),
    .O_9_1_2(op_O_9_1_2),
    .O_9_2_0(op_O_9_2_0),
    .O_9_2_1(op_O_9_2_1),
    .O_9_2_2(op_O_9_2_2),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_0_2(op_O_10_0_2),
    .O_10_1_0(op_O_10_1_0),
    .O_10_1_1(op_O_10_1_1),
    .O_10_1_2(op_O_10_1_2),
    .O_10_2_0(op_O_10_2_0),
    .O_10_2_1(op_O_10_2_1),
    .O_10_2_2(op_O_10_2_2),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_0_2(op_O_11_0_2),
    .O_11_1_0(op_O_11_1_0),
    .O_11_1_1(op_O_11_1_1),
    .O_11_1_2(op_O_11_1_2),
    .O_11_2_0(op_O_11_2_0),
    .O_11_2_1(op_O_11_2_1),
    .O_11_2_2(op_O_11_2_2),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_0_2(op_O_12_0_2),
    .O_12_1_0(op_O_12_1_0),
    .O_12_1_1(op_O_12_1_1),
    .O_12_1_2(op_O_12_1_2),
    .O_12_2_0(op_O_12_2_0),
    .O_12_2_1(op_O_12_2_1),
    .O_12_2_2(op_O_12_2_2),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_0_2(op_O_13_0_2),
    .O_13_1_0(op_O_13_1_0),
    .O_13_1_1(op_O_13_1_1),
    .O_13_1_2(op_O_13_1_2),
    .O_13_2_0(op_O_13_2_0),
    .O_13_2_1(op_O_13_2_1),
    .O_13_2_2(op_O_13_2_2),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_0_2(op_O_14_0_2),
    .O_14_1_0(op_O_14_1_0),
    .O_14_1_1(op_O_14_1_1),
    .O_14_1_2(op_O_14_1_2),
    .O_14_2_0(op_O_14_2_0),
    .O_14_2_1(op_O_14_2_1),
    .O_14_2_2(op_O_14_2_2),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_0_2(op_O_15_0_2),
    .O_15_1_0(op_O_15_1_0),
    .O_15_1_1(op_O_15_1_1),
    .O_15_1_2(op_O_15_1_2),
    .O_15_2_0(op_O_15_2_0),
    .O_15_2_1(op_O_15_2_1),
    .O_15_2_2(op_O_15_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_0_1_0 = op_O_0_1_0; // @[MapT.scala 15:7]
  assign O_0_1_1 = op_O_0_1_1; // @[MapT.scala 15:7]
  assign O_0_1_2 = op_O_0_1_2; // @[MapT.scala 15:7]
  assign O_0_2_0 = op_O_0_2_0; // @[MapT.scala 15:7]
  assign O_0_2_1 = op_O_0_2_1; // @[MapT.scala 15:7]
  assign O_0_2_2 = op_O_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_1_1_0 = op_O_1_1_0; // @[MapT.scala 15:7]
  assign O_1_1_1 = op_O_1_1_1; // @[MapT.scala 15:7]
  assign O_1_1_2 = op_O_1_1_2; // @[MapT.scala 15:7]
  assign O_1_2_0 = op_O_1_2_0; // @[MapT.scala 15:7]
  assign O_1_2_1 = op_O_1_2_1; // @[MapT.scala 15:7]
  assign O_1_2_2 = op_O_1_2_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_2_1_0 = op_O_2_1_0; // @[MapT.scala 15:7]
  assign O_2_1_1 = op_O_2_1_1; // @[MapT.scala 15:7]
  assign O_2_1_2 = op_O_2_1_2; // @[MapT.scala 15:7]
  assign O_2_2_0 = op_O_2_2_0; // @[MapT.scala 15:7]
  assign O_2_2_1 = op_O_2_2_1; // @[MapT.scala 15:7]
  assign O_2_2_2 = op_O_2_2_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign O_3_1_0 = op_O_3_1_0; // @[MapT.scala 15:7]
  assign O_3_1_1 = op_O_3_1_1; // @[MapT.scala 15:7]
  assign O_3_1_2 = op_O_3_1_2; // @[MapT.scala 15:7]
  assign O_3_2_0 = op_O_3_2_0; // @[MapT.scala 15:7]
  assign O_3_2_1 = op_O_3_2_1; // @[MapT.scala 15:7]
  assign O_3_2_2 = op_O_3_2_2; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_4_0_2 = op_O_4_0_2; // @[MapT.scala 15:7]
  assign O_4_1_0 = op_O_4_1_0; // @[MapT.scala 15:7]
  assign O_4_1_1 = op_O_4_1_1; // @[MapT.scala 15:7]
  assign O_4_1_2 = op_O_4_1_2; // @[MapT.scala 15:7]
  assign O_4_2_0 = op_O_4_2_0; // @[MapT.scala 15:7]
  assign O_4_2_1 = op_O_4_2_1; // @[MapT.scala 15:7]
  assign O_4_2_2 = op_O_4_2_2; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_5_0_2 = op_O_5_0_2; // @[MapT.scala 15:7]
  assign O_5_1_0 = op_O_5_1_0; // @[MapT.scala 15:7]
  assign O_5_1_1 = op_O_5_1_1; // @[MapT.scala 15:7]
  assign O_5_1_2 = op_O_5_1_2; // @[MapT.scala 15:7]
  assign O_5_2_0 = op_O_5_2_0; // @[MapT.scala 15:7]
  assign O_5_2_1 = op_O_5_2_1; // @[MapT.scala 15:7]
  assign O_5_2_2 = op_O_5_2_2; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_6_0_2 = op_O_6_0_2; // @[MapT.scala 15:7]
  assign O_6_1_0 = op_O_6_1_0; // @[MapT.scala 15:7]
  assign O_6_1_1 = op_O_6_1_1; // @[MapT.scala 15:7]
  assign O_6_1_2 = op_O_6_1_2; // @[MapT.scala 15:7]
  assign O_6_2_0 = op_O_6_2_0; // @[MapT.scala 15:7]
  assign O_6_2_1 = op_O_6_2_1; // @[MapT.scala 15:7]
  assign O_6_2_2 = op_O_6_2_2; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_7_0_2 = op_O_7_0_2; // @[MapT.scala 15:7]
  assign O_7_1_0 = op_O_7_1_0; // @[MapT.scala 15:7]
  assign O_7_1_1 = op_O_7_1_1; // @[MapT.scala 15:7]
  assign O_7_1_2 = op_O_7_1_2; // @[MapT.scala 15:7]
  assign O_7_2_0 = op_O_7_2_0; // @[MapT.scala 15:7]
  assign O_7_2_1 = op_O_7_2_1; // @[MapT.scala 15:7]
  assign O_7_2_2 = op_O_7_2_2; // @[MapT.scala 15:7]
  assign O_8_0_0 = op_O_8_0_0; // @[MapT.scala 15:7]
  assign O_8_0_1 = op_O_8_0_1; // @[MapT.scala 15:7]
  assign O_8_0_2 = op_O_8_0_2; // @[MapT.scala 15:7]
  assign O_8_1_0 = op_O_8_1_0; // @[MapT.scala 15:7]
  assign O_8_1_1 = op_O_8_1_1; // @[MapT.scala 15:7]
  assign O_8_1_2 = op_O_8_1_2; // @[MapT.scala 15:7]
  assign O_8_2_0 = op_O_8_2_0; // @[MapT.scala 15:7]
  assign O_8_2_1 = op_O_8_2_1; // @[MapT.scala 15:7]
  assign O_8_2_2 = op_O_8_2_2; // @[MapT.scala 15:7]
  assign O_9_0_0 = op_O_9_0_0; // @[MapT.scala 15:7]
  assign O_9_0_1 = op_O_9_0_1; // @[MapT.scala 15:7]
  assign O_9_0_2 = op_O_9_0_2; // @[MapT.scala 15:7]
  assign O_9_1_0 = op_O_9_1_0; // @[MapT.scala 15:7]
  assign O_9_1_1 = op_O_9_1_1; // @[MapT.scala 15:7]
  assign O_9_1_2 = op_O_9_1_2; // @[MapT.scala 15:7]
  assign O_9_2_0 = op_O_9_2_0; // @[MapT.scala 15:7]
  assign O_9_2_1 = op_O_9_2_1; // @[MapT.scala 15:7]
  assign O_9_2_2 = op_O_9_2_2; // @[MapT.scala 15:7]
  assign O_10_0_0 = op_O_10_0_0; // @[MapT.scala 15:7]
  assign O_10_0_1 = op_O_10_0_1; // @[MapT.scala 15:7]
  assign O_10_0_2 = op_O_10_0_2; // @[MapT.scala 15:7]
  assign O_10_1_0 = op_O_10_1_0; // @[MapT.scala 15:7]
  assign O_10_1_1 = op_O_10_1_1; // @[MapT.scala 15:7]
  assign O_10_1_2 = op_O_10_1_2; // @[MapT.scala 15:7]
  assign O_10_2_0 = op_O_10_2_0; // @[MapT.scala 15:7]
  assign O_10_2_1 = op_O_10_2_1; // @[MapT.scala 15:7]
  assign O_10_2_2 = op_O_10_2_2; // @[MapT.scala 15:7]
  assign O_11_0_0 = op_O_11_0_0; // @[MapT.scala 15:7]
  assign O_11_0_1 = op_O_11_0_1; // @[MapT.scala 15:7]
  assign O_11_0_2 = op_O_11_0_2; // @[MapT.scala 15:7]
  assign O_11_1_0 = op_O_11_1_0; // @[MapT.scala 15:7]
  assign O_11_1_1 = op_O_11_1_1; // @[MapT.scala 15:7]
  assign O_11_1_2 = op_O_11_1_2; // @[MapT.scala 15:7]
  assign O_11_2_0 = op_O_11_2_0; // @[MapT.scala 15:7]
  assign O_11_2_1 = op_O_11_2_1; // @[MapT.scala 15:7]
  assign O_11_2_2 = op_O_11_2_2; // @[MapT.scala 15:7]
  assign O_12_0_0 = op_O_12_0_0; // @[MapT.scala 15:7]
  assign O_12_0_1 = op_O_12_0_1; // @[MapT.scala 15:7]
  assign O_12_0_2 = op_O_12_0_2; // @[MapT.scala 15:7]
  assign O_12_1_0 = op_O_12_1_0; // @[MapT.scala 15:7]
  assign O_12_1_1 = op_O_12_1_1; // @[MapT.scala 15:7]
  assign O_12_1_2 = op_O_12_1_2; // @[MapT.scala 15:7]
  assign O_12_2_0 = op_O_12_2_0; // @[MapT.scala 15:7]
  assign O_12_2_1 = op_O_12_2_1; // @[MapT.scala 15:7]
  assign O_12_2_2 = op_O_12_2_2; // @[MapT.scala 15:7]
  assign O_13_0_0 = op_O_13_0_0; // @[MapT.scala 15:7]
  assign O_13_0_1 = op_O_13_0_1; // @[MapT.scala 15:7]
  assign O_13_0_2 = op_O_13_0_2; // @[MapT.scala 15:7]
  assign O_13_1_0 = op_O_13_1_0; // @[MapT.scala 15:7]
  assign O_13_1_1 = op_O_13_1_1; // @[MapT.scala 15:7]
  assign O_13_1_2 = op_O_13_1_2; // @[MapT.scala 15:7]
  assign O_13_2_0 = op_O_13_2_0; // @[MapT.scala 15:7]
  assign O_13_2_1 = op_O_13_2_1; // @[MapT.scala 15:7]
  assign O_13_2_2 = op_O_13_2_2; // @[MapT.scala 15:7]
  assign O_14_0_0 = op_O_14_0_0; // @[MapT.scala 15:7]
  assign O_14_0_1 = op_O_14_0_1; // @[MapT.scala 15:7]
  assign O_14_0_2 = op_O_14_0_2; // @[MapT.scala 15:7]
  assign O_14_1_0 = op_O_14_1_0; // @[MapT.scala 15:7]
  assign O_14_1_1 = op_O_14_1_1; // @[MapT.scala 15:7]
  assign O_14_1_2 = op_O_14_1_2; // @[MapT.scala 15:7]
  assign O_14_2_0 = op_O_14_2_0; // @[MapT.scala 15:7]
  assign O_14_2_1 = op_O_14_2_1; // @[MapT.scala 15:7]
  assign O_14_2_2 = op_O_14_2_2; // @[MapT.scala 15:7]
  assign O_15_0_0 = op_O_15_0_0; // @[MapT.scala 15:7]
  assign O_15_0_1 = op_O_15_0_1; // @[MapT.scala 15:7]
  assign O_15_0_2 = op_O_15_0_2; // @[MapT.scala 15:7]
  assign O_15_1_0 = op_O_15_1_0; // @[MapT.scala 15:7]
  assign O_15_1_1 = op_O_15_1_1; // @[MapT.scala 15:7]
  assign O_15_1_2 = op_O_15_1_2; // @[MapT.scala 15:7]
  assign O_15_2_0 = op_O_15_2_0; // @[MapT.scala 15:7]
  assign O_15_2_1 = op_O_15_2_1; // @[MapT.scala 15:7]
  assign O_15_2_2 = op_O_15_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0_0 = I_0_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_0_1 = I_0_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_0_2 = I_0_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_0_1_0 = I_0_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1_1 = I_0_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_0_1_2 = I_0_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_0_2_0 = I_0_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_0_2_1 = I_0_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2_2 = I_0_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0_0 = I_1_0_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_0_1 = I_1_0_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0_2 = I_1_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_1_0 = I_1_0_1_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1_1 = I_1_0_1_1; // @[MapT.scala 14:10]
  assign op_I_1_0_1_2 = I_1_0_1_2; // @[MapT.scala 14:10]
  assign op_I_1_0_2_0 = I_1_0_2_0; // @[MapT.scala 14:10]
  assign op_I_1_0_2_1 = I_1_0_2_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2_2 = I_1_0_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0_0 = I_2_0_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_0_1 = I_2_0_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0_2 = I_2_0_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_1_0 = I_2_0_1_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1_1 = I_2_0_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0_1_2 = I_2_0_1_2; // @[MapT.scala 14:10]
  assign op_I_2_0_2_0 = I_2_0_2_0; // @[MapT.scala 14:10]
  assign op_I_2_0_2_1 = I_2_0_2_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2_2 = I_2_0_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0_0 = I_3_0_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_0_1 = I_3_0_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0_2 = I_3_0_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_1_0 = I_3_0_1_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1_1 = I_3_0_1_1; // @[MapT.scala 14:10]
  assign op_I_3_0_1_2 = I_3_0_1_2; // @[MapT.scala 14:10]
  assign op_I_3_0_2_0 = I_3_0_2_0; // @[MapT.scala 14:10]
  assign op_I_3_0_2_1 = I_3_0_2_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2_2 = I_3_0_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0_0 = I_4_0_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_0_1 = I_4_0_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_0_2 = I_4_0_0_2; // @[MapT.scala 14:10]
  assign op_I_4_0_1_0 = I_4_0_1_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1_1 = I_4_0_1_1; // @[MapT.scala 14:10]
  assign op_I_4_0_1_2 = I_4_0_1_2; // @[MapT.scala 14:10]
  assign op_I_4_0_2_0 = I_4_0_2_0; // @[MapT.scala 14:10]
  assign op_I_4_0_2_1 = I_4_0_2_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2_2 = I_4_0_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0_0 = I_5_0_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_0_1 = I_5_0_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_0_2 = I_5_0_0_2; // @[MapT.scala 14:10]
  assign op_I_5_0_1_0 = I_5_0_1_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1_1 = I_5_0_1_1; // @[MapT.scala 14:10]
  assign op_I_5_0_1_2 = I_5_0_1_2; // @[MapT.scala 14:10]
  assign op_I_5_0_2_0 = I_5_0_2_0; // @[MapT.scala 14:10]
  assign op_I_5_0_2_1 = I_5_0_2_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2_2 = I_5_0_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0_0 = I_6_0_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_0_1 = I_6_0_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_0_2 = I_6_0_0_2; // @[MapT.scala 14:10]
  assign op_I_6_0_1_0 = I_6_0_1_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1_1 = I_6_0_1_1; // @[MapT.scala 14:10]
  assign op_I_6_0_1_2 = I_6_0_1_2; // @[MapT.scala 14:10]
  assign op_I_6_0_2_0 = I_6_0_2_0; // @[MapT.scala 14:10]
  assign op_I_6_0_2_1 = I_6_0_2_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2_2 = I_6_0_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0_0 = I_7_0_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_0_1 = I_7_0_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_0_2 = I_7_0_0_2; // @[MapT.scala 14:10]
  assign op_I_7_0_1_0 = I_7_0_1_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1_1 = I_7_0_1_1; // @[MapT.scala 14:10]
  assign op_I_7_0_1_2 = I_7_0_1_2; // @[MapT.scala 14:10]
  assign op_I_7_0_2_0 = I_7_0_2_0; // @[MapT.scala 14:10]
  assign op_I_7_0_2_1 = I_7_0_2_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2_2 = I_7_0_2_2; // @[MapT.scala 14:10]
  assign op_I_8_0_0_0 = I_8_0_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_0_1 = I_8_0_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_0_2 = I_8_0_0_2; // @[MapT.scala 14:10]
  assign op_I_8_0_1_0 = I_8_0_1_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1_1 = I_8_0_1_1; // @[MapT.scala 14:10]
  assign op_I_8_0_1_2 = I_8_0_1_2; // @[MapT.scala 14:10]
  assign op_I_8_0_2_0 = I_8_0_2_0; // @[MapT.scala 14:10]
  assign op_I_8_0_2_1 = I_8_0_2_1; // @[MapT.scala 14:10]
  assign op_I_8_0_2_2 = I_8_0_2_2; // @[MapT.scala 14:10]
  assign op_I_9_0_0_0 = I_9_0_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_0_1 = I_9_0_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_0_2 = I_9_0_0_2; // @[MapT.scala 14:10]
  assign op_I_9_0_1_0 = I_9_0_1_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1_1 = I_9_0_1_1; // @[MapT.scala 14:10]
  assign op_I_9_0_1_2 = I_9_0_1_2; // @[MapT.scala 14:10]
  assign op_I_9_0_2_0 = I_9_0_2_0; // @[MapT.scala 14:10]
  assign op_I_9_0_2_1 = I_9_0_2_1; // @[MapT.scala 14:10]
  assign op_I_9_0_2_2 = I_9_0_2_2; // @[MapT.scala 14:10]
  assign op_I_10_0_0_0 = I_10_0_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_0_1 = I_10_0_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_0_2 = I_10_0_0_2; // @[MapT.scala 14:10]
  assign op_I_10_0_1_0 = I_10_0_1_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1_1 = I_10_0_1_1; // @[MapT.scala 14:10]
  assign op_I_10_0_1_2 = I_10_0_1_2; // @[MapT.scala 14:10]
  assign op_I_10_0_2_0 = I_10_0_2_0; // @[MapT.scala 14:10]
  assign op_I_10_0_2_1 = I_10_0_2_1; // @[MapT.scala 14:10]
  assign op_I_10_0_2_2 = I_10_0_2_2; // @[MapT.scala 14:10]
  assign op_I_11_0_0_0 = I_11_0_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_0_1 = I_11_0_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_0_2 = I_11_0_0_2; // @[MapT.scala 14:10]
  assign op_I_11_0_1_0 = I_11_0_1_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1_1 = I_11_0_1_1; // @[MapT.scala 14:10]
  assign op_I_11_0_1_2 = I_11_0_1_2; // @[MapT.scala 14:10]
  assign op_I_11_0_2_0 = I_11_0_2_0; // @[MapT.scala 14:10]
  assign op_I_11_0_2_1 = I_11_0_2_1; // @[MapT.scala 14:10]
  assign op_I_11_0_2_2 = I_11_0_2_2; // @[MapT.scala 14:10]
  assign op_I_12_0_0_0 = I_12_0_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_0_1 = I_12_0_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_0_2 = I_12_0_0_2; // @[MapT.scala 14:10]
  assign op_I_12_0_1_0 = I_12_0_1_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1_1 = I_12_0_1_1; // @[MapT.scala 14:10]
  assign op_I_12_0_1_2 = I_12_0_1_2; // @[MapT.scala 14:10]
  assign op_I_12_0_2_0 = I_12_0_2_0; // @[MapT.scala 14:10]
  assign op_I_12_0_2_1 = I_12_0_2_1; // @[MapT.scala 14:10]
  assign op_I_12_0_2_2 = I_12_0_2_2; // @[MapT.scala 14:10]
  assign op_I_13_0_0_0 = I_13_0_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_0_1 = I_13_0_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_0_2 = I_13_0_0_2; // @[MapT.scala 14:10]
  assign op_I_13_0_1_0 = I_13_0_1_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1_1 = I_13_0_1_1; // @[MapT.scala 14:10]
  assign op_I_13_0_1_2 = I_13_0_1_2; // @[MapT.scala 14:10]
  assign op_I_13_0_2_0 = I_13_0_2_0; // @[MapT.scala 14:10]
  assign op_I_13_0_2_1 = I_13_0_2_1; // @[MapT.scala 14:10]
  assign op_I_13_0_2_2 = I_13_0_2_2; // @[MapT.scala 14:10]
  assign op_I_14_0_0_0 = I_14_0_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_0_1 = I_14_0_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_0_2 = I_14_0_0_2; // @[MapT.scala 14:10]
  assign op_I_14_0_1_0 = I_14_0_1_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1_1 = I_14_0_1_1; // @[MapT.scala 14:10]
  assign op_I_14_0_1_2 = I_14_0_1_2; // @[MapT.scala 14:10]
  assign op_I_14_0_2_0 = I_14_0_2_0; // @[MapT.scala 14:10]
  assign op_I_14_0_2_1 = I_14_0_2_1; // @[MapT.scala 14:10]
  assign op_I_14_0_2_2 = I_14_0_2_2; // @[MapT.scala 14:10]
  assign op_I_15_0_0_0 = I_15_0_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_0_1 = I_15_0_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_0_2 = I_15_0_0_2; // @[MapT.scala 14:10]
  assign op_I_15_0_1_0 = I_15_0_1_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1_1 = I_15_0_1_1; // @[MapT.scala 14:10]
  assign op_I_15_0_1_2 = I_15_0_1_2; // @[MapT.scala 14:10]
  assign op_I_15_0_2_0 = I_15_0_2_0; // @[MapT.scala 14:10]
  assign op_I_15_0_2_1 = I_15_0_2_1; // @[MapT.scala 14:10]
  assign op_I_15_0_2_2 = I_15_0_2_2; // @[MapT.scala 14:10]
endmodule
module InitialDelayCounter(
  input   clock,
  input   reset,
  output  valid_down
);
  reg  value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire  _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 1'h1; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 1'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 1'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module AtomTuple(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_t0b,
  output [7:0] O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Map2S_22(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_t0b,
  output [7:0] O_0_t1b,
  output [7:0] O_1_t0b,
  output [7:0] O_1_t1b,
  output [7:0] O_2_t0b,
  output [7:0] O_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  AtomTuple other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  AtomTuple other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_t0b(other_ops_1_O_t0b),
    .O_t1b(other_ops_1_O_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign O_2_t0b = other_ops_1_O_t0b; // @[Map2S.scala 24:12]
  assign O_2_t1b = other_ops_1_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
endmodule
module Map2S_23(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_1_2,
  input  [7:0] I0_2_0,
  input  [7:0] I0_2_1,
  input  [7:0] I0_2_2,
  output [7:0] O_0_0_t0b,
  output [7:0] O_0_0_t1b,
  output [7:0] O_0_1_t0b,
  output [7:0] O_0_1_t1b,
  output [7:0] O_0_2_t0b,
  output [7:0] O_0_2_t1b,
  output [7:0] O_1_0_t0b,
  output [7:0] O_1_0_t1b,
  output [7:0] O_1_1_t0b,
  output [7:0] O_1_1_t1b,
  output [7:0] O_1_2_t0b,
  output [7:0] O_1_2_t1b,
  output [7:0] O_2_0_t0b,
  output [7:0] O_2_0_t1b,
  output [7:0] O_2_1_t0b,
  output [7:0] O_2_1_t1b,
  output [7:0] O_2_2_t0b,
  output [7:0] O_2_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_t1b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  Map2S_22 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b),
    .O_1_t0b(fst_op_O_1_t0b),
    .O_1_t1b(fst_op_O_1_t1b),
    .O_2_t0b(fst_op_O_2_t0b),
    .O_2_t1b(fst_op_O_2_t1b)
  );
  Map2S_22 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_t0b(other_ops_0_O_0_t0b),
    .O_0_t1b(other_ops_0_O_0_t1b),
    .O_1_t0b(other_ops_0_O_1_t0b),
    .O_1_t1b(other_ops_0_O_1_t1b),
    .O_2_t0b(other_ops_0_O_2_t0b),
    .O_2_t1b(other_ops_0_O_2_t1b)
  );
  Map2S_22 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_t0b(other_ops_1_O_0_t0b),
    .O_0_t1b(other_ops_1_O_0_t1b),
    .O_1_t0b(other_ops_1_O_1_t0b),
    .O_1_t1b(other_ops_1_O_1_t1b),
    .O_2_t0b(other_ops_1_O_2_t0b),
    .O_2_t1b(other_ops_1_O_2_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign O_0_1_t0b = fst_op_O_1_t0b; // @[Map2S.scala 19:8]
  assign O_0_1_t1b = fst_op_O_1_t1b; // @[Map2S.scala 19:8]
  assign O_0_2_t0b = fst_op_O_2_t0b; // @[Map2S.scala 19:8]
  assign O_0_2_t1b = fst_op_O_2_t1b; // @[Map2S.scala 19:8]
  assign O_1_0_t0b = other_ops_0_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_1_0_t1b = other_ops_0_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_1_1_t0b = other_ops_0_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_1_1_t1b = other_ops_0_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_1_2_t0b = other_ops_0_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_1_2_t1b = other_ops_0_O_2_t1b; // @[Map2S.scala 24:12]
  assign O_2_0_t0b = other_ops_1_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_2_0_t1b = other_ops_1_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_2_1_t0b = other_ops_1_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_2_1_t1b = other_ops_1_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_2_2_t0b = other_ops_1_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_2_2_t1b = other_ops_1_O_2_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = 8'h0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = 8'h1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = 8'h0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = 8'h2; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = 8'h0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = 8'h0; // @[Map2S.scala 23:43]
endmodule
module LShift(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  wire [262:0] _GEN_0; // @[Arithmetic.scala 163:23]
  wire [262:0] _T; // @[Arithmetic.scala 163:23]
  assign _GEN_0 = {{255'd0}, I_t0b}; // @[Arithmetic.scala 163:23]
  assign _T = _GEN_0 << I_t1b; // @[Arithmetic.scala 163:23]
  assign valid_down = valid_up; // @[Arithmetic.scala 164:14]
  assign O = _T[7:0]; // @[Arithmetic.scala 163:5]
endmodule
module MapS_7(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  input  [7:0] I_1_t0b,
  input  [7:0] I_1_t1b,
  input  [7:0] I_2_t0b,
  input  [7:0] I_2_t1b,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  LShift fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  LShift other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t0b(other_ops_0_I_t0b),
    .I_t1b(other_ops_0_I_t1b),
    .O(other_ops_0_O)
  );
  LShift other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_t0b(other_ops_1_I_t0b),
    .I_t1b(other_ops_1_I_t1b),
    .O(other_ops_1_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t0b = I_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_t1b = I_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_t0b = I_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_t1b = I_2_t1b; // @[MapS.scala 20:41]
endmodule
module MapS_8(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_t0b,
  input  [7:0] I_0_0_t1b,
  input  [7:0] I_0_1_t0b,
  input  [7:0] I_0_1_t1b,
  input  [7:0] I_0_2_t0b,
  input  [7:0] I_0_2_t1b,
  input  [7:0] I_1_0_t0b,
  input  [7:0] I_1_0_t1b,
  input  [7:0] I_1_1_t0b,
  input  [7:0] I_1_1_t1b,
  input  [7:0] I_1_2_t0b,
  input  [7:0] I_1_2_t1b,
  input  [7:0] I_2_0_t0b,
  input  [7:0] I_2_0_t1b,
  input  [7:0] I_2_1_t0b,
  input  [7:0] I_2_1_t1b,
  input  [7:0] I_2_2_t0b,
  input  [7:0] I_2_2_t1b,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  MapS_7 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .I_1_t0b(fst_op_I_1_t0b),
    .I_1_t1b(fst_op_I_1_t1b),
    .I_2_t0b(fst_op_I_2_t0b),
    .I_2_t1b(fst_op_I_2_t1b),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  MapS_7 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_t0b(other_ops_0_I_0_t0b),
    .I_0_t1b(other_ops_0_I_0_t1b),
    .I_1_t0b(other_ops_0_I_1_t0b),
    .I_1_t1b(other_ops_0_I_1_t1b),
    .I_2_t0b(other_ops_0_I_2_t0b),
    .I_2_t1b(other_ops_0_I_2_t1b),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  MapS_7 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_t0b(other_ops_1_I_0_t0b),
    .I_0_t1b(other_ops_1_I_0_t1b),
    .I_1_t0b(other_ops_1_I_1_t0b),
    .I_1_t1b(other_ops_1_I_1_t1b),
    .I_2_t0b(other_ops_1_I_2_t0b),
    .I_2_t1b(other_ops_1_I_2_t1b),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t0b = I_0_1_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t1b = I_0_1_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t0b = I_0_2_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t1b = I_0_2_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_t0b = I_1_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_t1b = I_1_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t0b = I_1_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t1b = I_1_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t0b = I_1_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t1b = I_1_2_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_t0b = I_2_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_t1b = I_2_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t0b = I_2_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t1b = I_2_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t0b = I_2_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t1b = I_2_2_t1b; // @[MapS.scala 20:41]
endmodule
module AddNoValid(
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  assign O = I_t0b + I_t1b; // @[Arithmetic.scala 69:5]
endmodule
module ReduceS(
  input        clock,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O_0
);
  wire [7:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_1_O; // @[ReduceS.scala 20:43]
  reg [7:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_1;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  AddNoValid AddNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_1_I_t0b),
    .I_t1b(AddNoValid_1_I_t1b),
    .O(AddNoValid_1_O)
  );
  assign valid_down = _T_1; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = I_0; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = AddNoValid_1_O; // @[ReduceS.scala 36:18]
  assign AddNoValid_1_I_t0b = I_1; // @[ReduceS.scala 43:18]
  assign AddNoValid_1_I_t1b = I_2; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    _T_1 <= valid_up;
  end
endmodule
module MapS_9(
  input        clock,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  output [7:0] O_0_0,
  output [7:0] O_1_0,
  output [7:0] O_2_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  ReduceS fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .O_0(fst_op_O_0)
  );
  ReduceS other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0(other_ops_0_I_0),
    .I_1(other_ops_0_I_1),
    .I_2(other_ops_0_I_2),
    .O_0(other_ops_0_O_0)
  );
  ReduceS other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0(other_ops_1_I_0),
    .I_1(other_ops_1_I_1),
    .I_2(other_ops_1_I_2),
    .O_0(other_ops_1_O_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0 = I_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1 = I_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2 = I_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0 = I_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1 = I_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2 = I_2_2; // @[MapS.scala 20:41]
endmodule
module MapSNoValid(
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  output [7:0] O_0
);
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 28:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 28:22]
  wire [7:0] fst_op_O; // @[MapS.scala 28:22]
  AddNoValid fst_op ( // @[MapS.scala 28:22]
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign O_0 = fst_op_O; // @[MapS.scala 35:8]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 34:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 34:12]
endmodule
module ReduceS_1(
  input        clock,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_1_0,
  input  [7:0] I_2_0,
  output [7:0] O_0_0
);
  wire [7:0] MapSNoValid_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_O_0; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_1_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_1_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_1_O_0; // @[ReduceS.scala 20:43]
  reg [7:0] _T_0; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_1;
  MapSNoValid MapSNoValid ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_I_0_t0b),
    .I_0_t1b(MapSNoValid_I_0_t1b),
    .O_0(MapSNoValid_O_0)
  );
  MapSNoValid MapSNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_1_I_0_t0b),
    .I_0_t1b(MapSNoValid_1_I_0_t1b),
    .O_0(MapSNoValid_1_O_0)
  );
  assign valid_down = _T_1; // @[ReduceS.scala 47:14]
  assign O_0_0 = _T_0; // @[ReduceS.scala 27:14]
  assign MapSNoValid_I_0_t0b = I_2_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_I_0_t1b = MapSNoValid_1_O_0; // @[ReduceS.scala 36:18]
  assign MapSNoValid_1_I_0_t0b = I_0_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_1_I_0_t1b = I_1_0; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= MapSNoValid_O_0;
    _T_1 <= valid_up;
  end
endmodule
module InitialDelayCounter_1(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [1:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [1:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 2'h3; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 2'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 2'h3; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 2'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Map2S_24(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  output [7:0] O_0_t0b,
  output [7:0] O_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = 8'h4; // @[Map2S.scala 18:13]
endmodule
module Map2S_25(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  output [7:0] O_0_0_t0b,
  output [7:0] O_0_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  Map2S_24 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
endmodule
module RShift(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 143:14]
  assign O = I_t0b >> I_t1b; // @[Arithmetic.scala 142:5]
endmodule
module MapS_10(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  output [7:0] O_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  RShift fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
endmodule
module MapS_11(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_t0b,
  input  [7:0] I_0_0_t1b,
  output [7:0] O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  MapS_10 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
endmodule
module Module_0(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  output [7:0] O_0_0
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n146_valid_up; // @[Top.scala 16:22]
  wire  n146_valid_down; // @[Top.scala 16:22]
  wire [7:0] n146_I0_0_0; // @[Top.scala 16:22]
  wire [7:0] n146_I0_0_1; // @[Top.scala 16:22]
  wire [7:0] n146_I0_0_2; // @[Top.scala 16:22]
  wire [7:0] n146_I0_1_0; // @[Top.scala 16:22]
  wire [7:0] n146_I0_1_1; // @[Top.scala 16:22]
  wire [7:0] n146_I0_1_2; // @[Top.scala 16:22]
  wire [7:0] n146_I0_2_0; // @[Top.scala 16:22]
  wire [7:0] n146_I0_2_1; // @[Top.scala 16:22]
  wire [7:0] n146_I0_2_2; // @[Top.scala 16:22]
  wire [7:0] n146_O_0_0_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_0_0_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_0_1_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_0_1_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_0_2_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_0_2_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_1_0_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_1_0_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_1_1_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_1_1_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_1_2_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_1_2_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_2_0_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_2_0_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_2_1_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_2_1_t1b; // @[Top.scala 16:22]
  wire [7:0] n146_O_2_2_t0b; // @[Top.scala 16:22]
  wire [7:0] n146_O_2_2_t1b; // @[Top.scala 16:22]
  wire  n157_valid_up; // @[Top.scala 20:22]
  wire  n157_valid_down; // @[Top.scala 20:22]
  wire [7:0] n157_I_0_0_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_0_0_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_0_1_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_0_1_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_0_2_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_0_2_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_1_0_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_1_0_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_1_1_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_1_1_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_1_2_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_1_2_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_2_0_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_2_0_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_2_1_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_2_1_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_I_2_2_t0b; // @[Top.scala 20:22]
  wire [7:0] n157_I_2_2_t1b; // @[Top.scala 20:22]
  wire [7:0] n157_O_0_0; // @[Top.scala 20:22]
  wire [7:0] n157_O_0_1; // @[Top.scala 20:22]
  wire [7:0] n157_O_0_2; // @[Top.scala 20:22]
  wire [7:0] n157_O_1_0; // @[Top.scala 20:22]
  wire [7:0] n157_O_1_1; // @[Top.scala 20:22]
  wire [7:0] n157_O_1_2; // @[Top.scala 20:22]
  wire [7:0] n157_O_2_0; // @[Top.scala 20:22]
  wire [7:0] n157_O_2_1; // @[Top.scala 20:22]
  wire [7:0] n157_O_2_2; // @[Top.scala 20:22]
  wire  n162_clock; // @[Top.scala 23:22]
  wire  n162_valid_up; // @[Top.scala 23:22]
  wire  n162_valid_down; // @[Top.scala 23:22]
  wire [7:0] n162_I_0_0; // @[Top.scala 23:22]
  wire [7:0] n162_I_0_1; // @[Top.scala 23:22]
  wire [7:0] n162_I_0_2; // @[Top.scala 23:22]
  wire [7:0] n162_I_1_0; // @[Top.scala 23:22]
  wire [7:0] n162_I_1_1; // @[Top.scala 23:22]
  wire [7:0] n162_I_1_2; // @[Top.scala 23:22]
  wire [7:0] n162_I_2_0; // @[Top.scala 23:22]
  wire [7:0] n162_I_2_1; // @[Top.scala 23:22]
  wire [7:0] n162_I_2_2; // @[Top.scala 23:22]
  wire [7:0] n162_O_0_0; // @[Top.scala 23:22]
  wire [7:0] n162_O_1_0; // @[Top.scala 23:22]
  wire [7:0] n162_O_2_0; // @[Top.scala 23:22]
  wire  n167_clock; // @[Top.scala 26:22]
  wire  n167_valid_up; // @[Top.scala 26:22]
  wire  n167_valid_down; // @[Top.scala 26:22]
  wire [7:0] n167_I_0_0; // @[Top.scala 26:22]
  wire [7:0] n167_I_1_0; // @[Top.scala 26:22]
  wire [7:0] n167_I_2_0; // @[Top.scala 26:22]
  wire [7:0] n167_O_0_0; // @[Top.scala 26:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n170_valid_up; // @[Top.scala 30:22]
  wire  n170_valid_down; // @[Top.scala 30:22]
  wire [7:0] n170_I0_0_0; // @[Top.scala 30:22]
  wire [7:0] n170_O_0_0_t0b; // @[Top.scala 30:22]
  wire [7:0] n170_O_0_0_t1b; // @[Top.scala 30:22]
  wire  n181_valid_up; // @[Top.scala 34:22]
  wire  n181_valid_down; // @[Top.scala 34:22]
  wire [7:0] n181_I_0_0_t0b; // @[Top.scala 34:22]
  wire [7:0] n181_I_0_0_t1b; // @[Top.scala 34:22]
  wire [7:0] n181_O_0_0; // @[Top.scala 34:22]
  InitialDelayCounter InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  Map2S_23 n146 ( // @[Top.scala 16:22]
    .valid_up(n146_valid_up),
    .valid_down(n146_valid_down),
    .I0_0_0(n146_I0_0_0),
    .I0_0_1(n146_I0_0_1),
    .I0_0_2(n146_I0_0_2),
    .I0_1_0(n146_I0_1_0),
    .I0_1_1(n146_I0_1_1),
    .I0_1_2(n146_I0_1_2),
    .I0_2_0(n146_I0_2_0),
    .I0_2_1(n146_I0_2_1),
    .I0_2_2(n146_I0_2_2),
    .O_0_0_t0b(n146_O_0_0_t0b),
    .O_0_0_t1b(n146_O_0_0_t1b),
    .O_0_1_t0b(n146_O_0_1_t0b),
    .O_0_1_t1b(n146_O_0_1_t1b),
    .O_0_2_t0b(n146_O_0_2_t0b),
    .O_0_2_t1b(n146_O_0_2_t1b),
    .O_1_0_t0b(n146_O_1_0_t0b),
    .O_1_0_t1b(n146_O_1_0_t1b),
    .O_1_1_t0b(n146_O_1_1_t0b),
    .O_1_1_t1b(n146_O_1_1_t1b),
    .O_1_2_t0b(n146_O_1_2_t0b),
    .O_1_2_t1b(n146_O_1_2_t1b),
    .O_2_0_t0b(n146_O_2_0_t0b),
    .O_2_0_t1b(n146_O_2_0_t1b),
    .O_2_1_t0b(n146_O_2_1_t0b),
    .O_2_1_t1b(n146_O_2_1_t1b),
    .O_2_2_t0b(n146_O_2_2_t0b),
    .O_2_2_t1b(n146_O_2_2_t1b)
  );
  MapS_8 n157 ( // @[Top.scala 20:22]
    .valid_up(n157_valid_up),
    .valid_down(n157_valid_down),
    .I_0_0_t0b(n157_I_0_0_t0b),
    .I_0_0_t1b(n157_I_0_0_t1b),
    .I_0_1_t0b(n157_I_0_1_t0b),
    .I_0_1_t1b(n157_I_0_1_t1b),
    .I_0_2_t0b(n157_I_0_2_t0b),
    .I_0_2_t1b(n157_I_0_2_t1b),
    .I_1_0_t0b(n157_I_1_0_t0b),
    .I_1_0_t1b(n157_I_1_0_t1b),
    .I_1_1_t0b(n157_I_1_1_t0b),
    .I_1_1_t1b(n157_I_1_1_t1b),
    .I_1_2_t0b(n157_I_1_2_t0b),
    .I_1_2_t1b(n157_I_1_2_t1b),
    .I_2_0_t0b(n157_I_2_0_t0b),
    .I_2_0_t1b(n157_I_2_0_t1b),
    .I_2_1_t0b(n157_I_2_1_t0b),
    .I_2_1_t1b(n157_I_2_1_t1b),
    .I_2_2_t0b(n157_I_2_2_t0b),
    .I_2_2_t1b(n157_I_2_2_t1b),
    .O_0_0(n157_O_0_0),
    .O_0_1(n157_O_0_1),
    .O_0_2(n157_O_0_2),
    .O_1_0(n157_O_1_0),
    .O_1_1(n157_O_1_1),
    .O_1_2(n157_O_1_2),
    .O_2_0(n157_O_2_0),
    .O_2_1(n157_O_2_1),
    .O_2_2(n157_O_2_2)
  );
  MapS_9 n162 ( // @[Top.scala 23:22]
    .clock(n162_clock),
    .valid_up(n162_valid_up),
    .valid_down(n162_valid_down),
    .I_0_0(n162_I_0_0),
    .I_0_1(n162_I_0_1),
    .I_0_2(n162_I_0_2),
    .I_1_0(n162_I_1_0),
    .I_1_1(n162_I_1_1),
    .I_1_2(n162_I_1_2),
    .I_2_0(n162_I_2_0),
    .I_2_1(n162_I_2_1),
    .I_2_2(n162_I_2_2),
    .O_0_0(n162_O_0_0),
    .O_1_0(n162_O_1_0),
    .O_2_0(n162_O_2_0)
  );
  ReduceS_1 n167 ( // @[Top.scala 26:22]
    .clock(n167_clock),
    .valid_up(n167_valid_up),
    .valid_down(n167_valid_down),
    .I_0_0(n167_I_0_0),
    .I_1_0(n167_I_1_0),
    .I_2_0(n167_I_2_0),
    .O_0_0(n167_O_0_0)
  );
  InitialDelayCounter_1 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  Map2S_25 n170 ( // @[Top.scala 30:22]
    .valid_up(n170_valid_up),
    .valid_down(n170_valid_down),
    .I0_0_0(n170_I0_0_0),
    .O_0_0_t0b(n170_O_0_0_t0b),
    .O_0_0_t1b(n170_O_0_0_t1b)
  );
  MapS_11 n181 ( // @[Top.scala 34:22]
    .valid_up(n181_valid_up),
    .valid_down(n181_valid_down),
    .I_0_0_t0b(n181_I_0_0_t0b),
    .I_0_0_t1b(n181_I_0_0_t1b),
    .O_0_0(n181_O_0_0)
  );
  assign valid_down = n181_valid_down; // @[Top.scala 38:16]
  assign O_0_0 = n181_O_0_0; // @[Top.scala 37:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n146_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 19:19]
  assign n146_I0_0_0 = I_0_0; // @[Top.scala 17:13]
  assign n146_I0_0_1 = I_0_1; // @[Top.scala 17:13]
  assign n146_I0_0_2 = I_0_2; // @[Top.scala 17:13]
  assign n146_I0_1_0 = I_1_0; // @[Top.scala 17:13]
  assign n146_I0_1_1 = I_1_1; // @[Top.scala 17:13]
  assign n146_I0_1_2 = I_1_2; // @[Top.scala 17:13]
  assign n146_I0_2_0 = I_2_0; // @[Top.scala 17:13]
  assign n146_I0_2_1 = I_2_1; // @[Top.scala 17:13]
  assign n146_I0_2_2 = I_2_2; // @[Top.scala 17:13]
  assign n157_valid_up = n146_valid_down; // @[Top.scala 22:19]
  assign n157_I_0_0_t0b = n146_O_0_0_t0b; // @[Top.scala 21:12]
  assign n157_I_0_0_t1b = n146_O_0_0_t1b; // @[Top.scala 21:12]
  assign n157_I_0_1_t0b = n146_O_0_1_t0b; // @[Top.scala 21:12]
  assign n157_I_0_1_t1b = n146_O_0_1_t1b; // @[Top.scala 21:12]
  assign n157_I_0_2_t0b = n146_O_0_2_t0b; // @[Top.scala 21:12]
  assign n157_I_0_2_t1b = n146_O_0_2_t1b; // @[Top.scala 21:12]
  assign n157_I_1_0_t0b = n146_O_1_0_t0b; // @[Top.scala 21:12]
  assign n157_I_1_0_t1b = n146_O_1_0_t1b; // @[Top.scala 21:12]
  assign n157_I_1_1_t0b = n146_O_1_1_t0b; // @[Top.scala 21:12]
  assign n157_I_1_1_t1b = n146_O_1_1_t1b; // @[Top.scala 21:12]
  assign n157_I_1_2_t0b = n146_O_1_2_t0b; // @[Top.scala 21:12]
  assign n157_I_1_2_t1b = n146_O_1_2_t1b; // @[Top.scala 21:12]
  assign n157_I_2_0_t0b = n146_O_2_0_t0b; // @[Top.scala 21:12]
  assign n157_I_2_0_t1b = n146_O_2_0_t1b; // @[Top.scala 21:12]
  assign n157_I_2_1_t0b = n146_O_2_1_t0b; // @[Top.scala 21:12]
  assign n157_I_2_1_t1b = n146_O_2_1_t1b; // @[Top.scala 21:12]
  assign n157_I_2_2_t0b = n146_O_2_2_t0b; // @[Top.scala 21:12]
  assign n157_I_2_2_t1b = n146_O_2_2_t1b; // @[Top.scala 21:12]
  assign n162_clock = clock;
  assign n162_valid_up = n157_valid_down; // @[Top.scala 25:19]
  assign n162_I_0_0 = n157_O_0_0; // @[Top.scala 24:12]
  assign n162_I_0_1 = n157_O_0_1; // @[Top.scala 24:12]
  assign n162_I_0_2 = n157_O_0_2; // @[Top.scala 24:12]
  assign n162_I_1_0 = n157_O_1_0; // @[Top.scala 24:12]
  assign n162_I_1_1 = n157_O_1_1; // @[Top.scala 24:12]
  assign n162_I_1_2 = n157_O_1_2; // @[Top.scala 24:12]
  assign n162_I_2_0 = n157_O_2_0; // @[Top.scala 24:12]
  assign n162_I_2_1 = n157_O_2_1; // @[Top.scala 24:12]
  assign n162_I_2_2 = n157_O_2_2; // @[Top.scala 24:12]
  assign n167_clock = clock;
  assign n167_valid_up = n162_valid_down; // @[Top.scala 28:19]
  assign n167_I_0_0 = n162_O_0_0; // @[Top.scala 27:12]
  assign n167_I_1_0 = n162_O_1_0; // @[Top.scala 27:12]
  assign n167_I_2_0 = n162_O_2_0; // @[Top.scala 27:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n170_valid_up = n167_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 33:19]
  assign n170_I0_0_0 = n167_O_0_0; // @[Top.scala 31:13]
  assign n181_valid_up = n170_valid_down; // @[Top.scala 36:19]
  assign n181_I_0_0_t0b = n170_O_0_0_t0b; // @[Top.scala 35:12]
  assign n181_I_0_0_t1b = n170_O_0_0_t1b; // @[Top.scala 35:12]
endmodule
module MapS_12(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_1_1_2,
  input  [7:0] I_1_2_0,
  input  [7:0] I_1_2_1,
  input  [7:0] I_1_2_2,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_0_2,
  input  [7:0] I_2_1_0,
  input  [7:0] I_2_1_1,
  input  [7:0] I_2_1_2,
  input  [7:0] I_2_2_0,
  input  [7:0] I_2_2_1,
  input  [7:0] I_2_2_2,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_0_2,
  input  [7:0] I_3_1_0,
  input  [7:0] I_3_1_1,
  input  [7:0] I_3_1_2,
  input  [7:0] I_3_2_0,
  input  [7:0] I_3_2_1,
  input  [7:0] I_3_2_2,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_0_2,
  input  [7:0] I_4_1_0,
  input  [7:0] I_4_1_1,
  input  [7:0] I_4_1_2,
  input  [7:0] I_4_2_0,
  input  [7:0] I_4_2_1,
  input  [7:0] I_4_2_2,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_0_2,
  input  [7:0] I_5_1_0,
  input  [7:0] I_5_1_1,
  input  [7:0] I_5_1_2,
  input  [7:0] I_5_2_0,
  input  [7:0] I_5_2_1,
  input  [7:0] I_5_2_2,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_0_2,
  input  [7:0] I_6_1_0,
  input  [7:0] I_6_1_1,
  input  [7:0] I_6_1_2,
  input  [7:0] I_6_2_0,
  input  [7:0] I_6_2_1,
  input  [7:0] I_6_2_2,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_0_2,
  input  [7:0] I_7_1_0,
  input  [7:0] I_7_1_1,
  input  [7:0] I_7_1_2,
  input  [7:0] I_7_2_0,
  input  [7:0] I_7_2_1,
  input  [7:0] I_7_2_2,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_8_0_2,
  input  [7:0] I_8_1_0,
  input  [7:0] I_8_1_1,
  input  [7:0] I_8_1_2,
  input  [7:0] I_8_2_0,
  input  [7:0] I_8_2_1,
  input  [7:0] I_8_2_2,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_9_0_2,
  input  [7:0] I_9_1_0,
  input  [7:0] I_9_1_1,
  input  [7:0] I_9_1_2,
  input  [7:0] I_9_2_0,
  input  [7:0] I_9_2_1,
  input  [7:0] I_9_2_2,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_10_0_2,
  input  [7:0] I_10_1_0,
  input  [7:0] I_10_1_1,
  input  [7:0] I_10_1_2,
  input  [7:0] I_10_2_0,
  input  [7:0] I_10_2_1,
  input  [7:0] I_10_2_2,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_11_0_2,
  input  [7:0] I_11_1_0,
  input  [7:0] I_11_1_1,
  input  [7:0] I_11_1_2,
  input  [7:0] I_11_2_0,
  input  [7:0] I_11_2_1,
  input  [7:0] I_11_2_2,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_12_0_2,
  input  [7:0] I_12_1_0,
  input  [7:0] I_12_1_1,
  input  [7:0] I_12_1_2,
  input  [7:0] I_12_2_0,
  input  [7:0] I_12_2_1,
  input  [7:0] I_12_2_2,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_13_0_2,
  input  [7:0] I_13_1_0,
  input  [7:0] I_13_1_1,
  input  [7:0] I_13_1_2,
  input  [7:0] I_13_2_0,
  input  [7:0] I_13_2_1,
  input  [7:0] I_13_2_2,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_14_0_2,
  input  [7:0] I_14_1_0,
  input  [7:0] I_14_1_1,
  input  [7:0] I_14_1_2,
  input  [7:0] I_14_2_0,
  input  [7:0] I_14_2_1,
  input  [7:0] I_14_2_2,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  input  [7:0] I_15_0_2,
  input  [7:0] I_15_1_0,
  input  [7:0] I_15_1_1,
  input  [7:0] I_15_1_2,
  input  [7:0] I_15_2_0,
  input  [7:0] I_15_2_1,
  input  [7:0] I_15_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0,
  output [7:0] O_8_0_0,
  output [7:0] O_9_0_0,
  output [7:0] O_10_0_0,
  output [7:0] O_11_0_0,
  output [7:0] O_12_0_0,
  output [7:0] O_13_0_0,
  output [7:0] O_14_0_0,
  output [7:0] O_15_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_2_clock; // @[MapS.scala 10:86]
  wire  other_ops_2_reset; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_3_clock; // @[MapS.scala 10:86]
  wire  other_ops_3_reset; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_4_clock; // @[MapS.scala 10:86]
  wire  other_ops_4_reset; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_5_clock; // @[MapS.scala 10:86]
  wire  other_ops_5_reset; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_6_clock; // @[MapS.scala 10:86]
  wire  other_ops_6_reset; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_7_clock; // @[MapS.scala 10:86]
  wire  other_ops_7_reset; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_8_clock; // @[MapS.scala 10:86]
  wire  other_ops_8_reset; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_9_clock; // @[MapS.scala 10:86]
  wire  other_ops_9_reset; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_10_clock; // @[MapS.scala 10:86]
  wire  other_ops_10_reset; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_11_clock; // @[MapS.scala 10:86]
  wire  other_ops_11_reset; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_12_clock; // @[MapS.scala 10:86]
  wire  other_ops_12_reset; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_13_clock; // @[MapS.scala 10:86]
  wire  other_ops_13_reset; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_14_clock; // @[MapS.scala 10:86]
  wire  other_ops_14_reset; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Module_0 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .I_1_0(fst_op_I_1_0),
    .I_1_1(fst_op_I_1_1),
    .I_1_2(fst_op_I_1_2),
    .I_2_0(fst_op_I_2_0),
    .I_2_1(fst_op_I_2_1),
    .I_2_2(fst_op_I_2_2),
    .O_0_0(fst_op_O_0_0)
  );
  Module_0 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .I_1_0(other_ops_0_I_1_0),
    .I_1_1(other_ops_0_I_1_1),
    .I_1_2(other_ops_0_I_1_2),
    .I_2_0(other_ops_0_I_2_0),
    .I_2_1(other_ops_0_I_2_1),
    .I_2_2(other_ops_0_I_2_2),
    .O_0_0(other_ops_0_O_0_0)
  );
  Module_0 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .I_1_0(other_ops_1_I_1_0),
    .I_1_1(other_ops_1_I_1_1),
    .I_1_2(other_ops_1_I_1_2),
    .I_2_0(other_ops_1_I_2_0),
    .I_2_1(other_ops_1_I_2_1),
    .I_2_2(other_ops_1_I_2_2),
    .O_0_0(other_ops_1_O_0_0)
  );
  Module_0 other_ops_2 ( // @[MapS.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .I_1_0(other_ops_2_I_1_0),
    .I_1_1(other_ops_2_I_1_1),
    .I_1_2(other_ops_2_I_1_2),
    .I_2_0(other_ops_2_I_2_0),
    .I_2_1(other_ops_2_I_2_1),
    .I_2_2(other_ops_2_I_2_2),
    .O_0_0(other_ops_2_O_0_0)
  );
  Module_0 other_ops_3 ( // @[MapS.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_0_2(other_ops_3_I_0_2),
    .I_1_0(other_ops_3_I_1_0),
    .I_1_1(other_ops_3_I_1_1),
    .I_1_2(other_ops_3_I_1_2),
    .I_2_0(other_ops_3_I_2_0),
    .I_2_1(other_ops_3_I_2_1),
    .I_2_2(other_ops_3_I_2_2),
    .O_0_0(other_ops_3_O_0_0)
  );
  Module_0 other_ops_4 ( // @[MapS.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_0_2(other_ops_4_I_0_2),
    .I_1_0(other_ops_4_I_1_0),
    .I_1_1(other_ops_4_I_1_1),
    .I_1_2(other_ops_4_I_1_2),
    .I_2_0(other_ops_4_I_2_0),
    .I_2_1(other_ops_4_I_2_1),
    .I_2_2(other_ops_4_I_2_2),
    .O_0_0(other_ops_4_O_0_0)
  );
  Module_0 other_ops_5 ( // @[MapS.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_0_2(other_ops_5_I_0_2),
    .I_1_0(other_ops_5_I_1_0),
    .I_1_1(other_ops_5_I_1_1),
    .I_1_2(other_ops_5_I_1_2),
    .I_2_0(other_ops_5_I_2_0),
    .I_2_1(other_ops_5_I_2_1),
    .I_2_2(other_ops_5_I_2_2),
    .O_0_0(other_ops_5_O_0_0)
  );
  Module_0 other_ops_6 ( // @[MapS.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_0_2(other_ops_6_I_0_2),
    .I_1_0(other_ops_6_I_1_0),
    .I_1_1(other_ops_6_I_1_1),
    .I_1_2(other_ops_6_I_1_2),
    .I_2_0(other_ops_6_I_2_0),
    .I_2_1(other_ops_6_I_2_1),
    .I_2_2(other_ops_6_I_2_2),
    .O_0_0(other_ops_6_O_0_0)
  );
  Module_0 other_ops_7 ( // @[MapS.scala 10:86]
    .clock(other_ops_7_clock),
    .reset(other_ops_7_reset),
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0(other_ops_7_I_0_0),
    .I_0_1(other_ops_7_I_0_1),
    .I_0_2(other_ops_7_I_0_2),
    .I_1_0(other_ops_7_I_1_0),
    .I_1_1(other_ops_7_I_1_1),
    .I_1_2(other_ops_7_I_1_2),
    .I_2_0(other_ops_7_I_2_0),
    .I_2_1(other_ops_7_I_2_1),
    .I_2_2(other_ops_7_I_2_2),
    .O_0_0(other_ops_7_O_0_0)
  );
  Module_0 other_ops_8 ( // @[MapS.scala 10:86]
    .clock(other_ops_8_clock),
    .reset(other_ops_8_reset),
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0(other_ops_8_I_0_0),
    .I_0_1(other_ops_8_I_0_1),
    .I_0_2(other_ops_8_I_0_2),
    .I_1_0(other_ops_8_I_1_0),
    .I_1_1(other_ops_8_I_1_1),
    .I_1_2(other_ops_8_I_1_2),
    .I_2_0(other_ops_8_I_2_0),
    .I_2_1(other_ops_8_I_2_1),
    .I_2_2(other_ops_8_I_2_2),
    .O_0_0(other_ops_8_O_0_0)
  );
  Module_0 other_ops_9 ( // @[MapS.scala 10:86]
    .clock(other_ops_9_clock),
    .reset(other_ops_9_reset),
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0(other_ops_9_I_0_0),
    .I_0_1(other_ops_9_I_0_1),
    .I_0_2(other_ops_9_I_0_2),
    .I_1_0(other_ops_9_I_1_0),
    .I_1_1(other_ops_9_I_1_1),
    .I_1_2(other_ops_9_I_1_2),
    .I_2_0(other_ops_9_I_2_0),
    .I_2_1(other_ops_9_I_2_1),
    .I_2_2(other_ops_9_I_2_2),
    .O_0_0(other_ops_9_O_0_0)
  );
  Module_0 other_ops_10 ( // @[MapS.scala 10:86]
    .clock(other_ops_10_clock),
    .reset(other_ops_10_reset),
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0(other_ops_10_I_0_0),
    .I_0_1(other_ops_10_I_0_1),
    .I_0_2(other_ops_10_I_0_2),
    .I_1_0(other_ops_10_I_1_0),
    .I_1_1(other_ops_10_I_1_1),
    .I_1_2(other_ops_10_I_1_2),
    .I_2_0(other_ops_10_I_2_0),
    .I_2_1(other_ops_10_I_2_1),
    .I_2_2(other_ops_10_I_2_2),
    .O_0_0(other_ops_10_O_0_0)
  );
  Module_0 other_ops_11 ( // @[MapS.scala 10:86]
    .clock(other_ops_11_clock),
    .reset(other_ops_11_reset),
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0(other_ops_11_I_0_0),
    .I_0_1(other_ops_11_I_0_1),
    .I_0_2(other_ops_11_I_0_2),
    .I_1_0(other_ops_11_I_1_0),
    .I_1_1(other_ops_11_I_1_1),
    .I_1_2(other_ops_11_I_1_2),
    .I_2_0(other_ops_11_I_2_0),
    .I_2_1(other_ops_11_I_2_1),
    .I_2_2(other_ops_11_I_2_2),
    .O_0_0(other_ops_11_O_0_0)
  );
  Module_0 other_ops_12 ( // @[MapS.scala 10:86]
    .clock(other_ops_12_clock),
    .reset(other_ops_12_reset),
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0(other_ops_12_I_0_0),
    .I_0_1(other_ops_12_I_0_1),
    .I_0_2(other_ops_12_I_0_2),
    .I_1_0(other_ops_12_I_1_0),
    .I_1_1(other_ops_12_I_1_1),
    .I_1_2(other_ops_12_I_1_2),
    .I_2_0(other_ops_12_I_2_0),
    .I_2_1(other_ops_12_I_2_1),
    .I_2_2(other_ops_12_I_2_2),
    .O_0_0(other_ops_12_O_0_0)
  );
  Module_0 other_ops_13 ( // @[MapS.scala 10:86]
    .clock(other_ops_13_clock),
    .reset(other_ops_13_reset),
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0(other_ops_13_I_0_0),
    .I_0_1(other_ops_13_I_0_1),
    .I_0_2(other_ops_13_I_0_2),
    .I_1_0(other_ops_13_I_1_0),
    .I_1_1(other_ops_13_I_1_1),
    .I_1_2(other_ops_13_I_1_2),
    .I_2_0(other_ops_13_I_2_0),
    .I_2_1(other_ops_13_I_2_1),
    .I_2_2(other_ops_13_I_2_2),
    .O_0_0(other_ops_13_O_0_0)
  );
  Module_0 other_ops_14 ( // @[MapS.scala 10:86]
    .clock(other_ops_14_clock),
    .reset(other_ops_14_reset),
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0(other_ops_14_I_0_0),
    .I_0_1(other_ops_14_I_0_1),
    .I_0_2(other_ops_14_I_0_2),
    .I_1_0(other_ops_14_I_1_0),
    .I_1_1(other_ops_14_I_1_1),
    .I_1_2(other_ops_14_I_1_2),
    .I_2_0(other_ops_14_I_2_0),
    .I_2_1(other_ops_14_I_2_1),
    .I_2_2(other_ops_14_I_2_2),
    .O_0_0(other_ops_14_O_0_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[MapS.scala 21:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[MapS.scala 21:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[MapS.scala 21:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[MapS.scala 21:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[MapS.scala 21:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[MapS.scala 21:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[MapS.scala 21:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_1_0 = I_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_1_1 = I_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_1_2 = I_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_2_0 = I_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_2_1 = I_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_2_2 = I_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_0 = I_1_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_1 = I_1_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_2 = I_1_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_0 = I_1_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_1 = I_1_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_2 = I_1_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_0 = I_2_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_1 = I_2_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_2 = I_2_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_0 = I_2_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_1 = I_2_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_2 = I_2_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_2_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_0 = I_3_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_1 = I_3_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_2 = I_3_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_0 = I_3_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_1 = I_3_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_2 = I_3_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_3_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2 = I_4_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_0 = I_4_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_1 = I_4_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_2 = I_4_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_0 = I_4_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_1 = I_4_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_2 = I_4_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_4_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2 = I_5_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_0 = I_5_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_1 = I_5_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_2 = I_5_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_0 = I_5_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_1 = I_5_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_2 = I_5_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_5_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2 = I_6_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_0 = I_6_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_1 = I_6_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_2 = I_6_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_0 = I_6_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_1 = I_6_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_2 = I_6_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_6_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2 = I_7_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_0 = I_7_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_1 = I_7_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_2 = I_7_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_0 = I_7_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_1 = I_7_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_2 = I_7_2_2; // @[MapS.scala 20:41]
  assign other_ops_7_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_7_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0 = I_8_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1 = I_8_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2 = I_8_0_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_1_0 = I_8_1_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_1_1 = I_8_1_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_1_2 = I_8_1_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_2_0 = I_8_2_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_2_1 = I_8_2_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_2_2 = I_8_2_2; // @[MapS.scala 20:41]
  assign other_ops_8_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_8_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0 = I_9_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1 = I_9_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2 = I_9_0_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_1_0 = I_9_1_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_1_1 = I_9_1_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_1_2 = I_9_1_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_2_0 = I_9_2_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_2_1 = I_9_2_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_2_2 = I_9_2_2; // @[MapS.scala 20:41]
  assign other_ops_9_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_9_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0 = I_10_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1 = I_10_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2 = I_10_0_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_1_0 = I_10_1_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_1_1 = I_10_1_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_1_2 = I_10_1_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_2_0 = I_10_2_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_2_1 = I_10_2_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_2_2 = I_10_2_2; // @[MapS.scala 20:41]
  assign other_ops_10_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_10_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0 = I_11_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1 = I_11_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2 = I_11_0_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_1_0 = I_11_1_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_1_1 = I_11_1_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_1_2 = I_11_1_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_2_0 = I_11_2_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_2_1 = I_11_2_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_2_2 = I_11_2_2; // @[MapS.scala 20:41]
  assign other_ops_11_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_11_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0 = I_12_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1 = I_12_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2 = I_12_0_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_1_0 = I_12_1_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_1_1 = I_12_1_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_1_2 = I_12_1_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_2_0 = I_12_2_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_2_1 = I_12_2_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_2_2 = I_12_2_2; // @[MapS.scala 20:41]
  assign other_ops_12_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_12_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0 = I_13_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1 = I_13_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2 = I_13_0_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_1_0 = I_13_1_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_1_1 = I_13_1_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_1_2 = I_13_1_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_2_0 = I_13_2_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_2_1 = I_13_2_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_2_2 = I_13_2_2; // @[MapS.scala 20:41]
  assign other_ops_13_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_13_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0 = I_14_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1 = I_14_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2 = I_14_0_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_1_0 = I_14_1_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_1_1 = I_14_1_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_1_2 = I_14_1_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_2_0 = I_14_2_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_2_1 = I_14_2_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_2_2 = I_14_2_2; // @[MapS.scala 20:41]
  assign other_ops_14_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_14_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0 = I_15_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1 = I_15_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2 = I_15_0_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_1_0 = I_15_1_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_1_1 = I_15_1_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_1_2 = I_15_1_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_2_0 = I_15_2_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_2_1 = I_15_2_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_2_2 = I_15_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_4(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_1_1_2,
  input  [7:0] I_1_2_0,
  input  [7:0] I_1_2_1,
  input  [7:0] I_1_2_2,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_0_2,
  input  [7:0] I_2_1_0,
  input  [7:0] I_2_1_1,
  input  [7:0] I_2_1_2,
  input  [7:0] I_2_2_0,
  input  [7:0] I_2_2_1,
  input  [7:0] I_2_2_2,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_0_2,
  input  [7:0] I_3_1_0,
  input  [7:0] I_3_1_1,
  input  [7:0] I_3_1_2,
  input  [7:0] I_3_2_0,
  input  [7:0] I_3_2_1,
  input  [7:0] I_3_2_2,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_0_2,
  input  [7:0] I_4_1_0,
  input  [7:0] I_4_1_1,
  input  [7:0] I_4_1_2,
  input  [7:0] I_4_2_0,
  input  [7:0] I_4_2_1,
  input  [7:0] I_4_2_2,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_0_2,
  input  [7:0] I_5_1_0,
  input  [7:0] I_5_1_1,
  input  [7:0] I_5_1_2,
  input  [7:0] I_5_2_0,
  input  [7:0] I_5_2_1,
  input  [7:0] I_5_2_2,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_0_2,
  input  [7:0] I_6_1_0,
  input  [7:0] I_6_1_1,
  input  [7:0] I_6_1_2,
  input  [7:0] I_6_2_0,
  input  [7:0] I_6_2_1,
  input  [7:0] I_6_2_2,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_0_2,
  input  [7:0] I_7_1_0,
  input  [7:0] I_7_1_1,
  input  [7:0] I_7_1_2,
  input  [7:0] I_7_2_0,
  input  [7:0] I_7_2_1,
  input  [7:0] I_7_2_2,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_8_0_2,
  input  [7:0] I_8_1_0,
  input  [7:0] I_8_1_1,
  input  [7:0] I_8_1_2,
  input  [7:0] I_8_2_0,
  input  [7:0] I_8_2_1,
  input  [7:0] I_8_2_2,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_9_0_2,
  input  [7:0] I_9_1_0,
  input  [7:0] I_9_1_1,
  input  [7:0] I_9_1_2,
  input  [7:0] I_9_2_0,
  input  [7:0] I_9_2_1,
  input  [7:0] I_9_2_2,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_10_0_2,
  input  [7:0] I_10_1_0,
  input  [7:0] I_10_1_1,
  input  [7:0] I_10_1_2,
  input  [7:0] I_10_2_0,
  input  [7:0] I_10_2_1,
  input  [7:0] I_10_2_2,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_11_0_2,
  input  [7:0] I_11_1_0,
  input  [7:0] I_11_1_1,
  input  [7:0] I_11_1_2,
  input  [7:0] I_11_2_0,
  input  [7:0] I_11_2_1,
  input  [7:0] I_11_2_2,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_12_0_2,
  input  [7:0] I_12_1_0,
  input  [7:0] I_12_1_1,
  input  [7:0] I_12_1_2,
  input  [7:0] I_12_2_0,
  input  [7:0] I_12_2_1,
  input  [7:0] I_12_2_2,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_13_0_2,
  input  [7:0] I_13_1_0,
  input  [7:0] I_13_1_1,
  input  [7:0] I_13_1_2,
  input  [7:0] I_13_2_0,
  input  [7:0] I_13_2_1,
  input  [7:0] I_13_2_2,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_14_0_2,
  input  [7:0] I_14_1_0,
  input  [7:0] I_14_1_1,
  input  [7:0] I_14_1_2,
  input  [7:0] I_14_2_0,
  input  [7:0] I_14_2_1,
  input  [7:0] I_14_2_2,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  input  [7:0] I_15_0_2,
  input  [7:0] I_15_1_0,
  input  [7:0] I_15_1_1,
  input  [7:0] I_15_1_2,
  input  [7:0] I_15_2_0,
  input  [7:0] I_15_2_1,
  input  [7:0] I_15_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0,
  output [7:0] O_8_0_0,
  output [7:0] O_9_0_0,
  output [7:0] O_10_0_0,
  output [7:0] O_11_0_0,
  output [7:0] O_12_0_0,
  output [7:0] O_13_0_0,
  output [7:0] O_14_0_0,
  output [7:0] O_15_0_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_0; // @[MapT.scala 8:20]
  MapS_12 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_4_1_2(op_I_4_1_2),
    .I_4_2_0(op_I_4_2_0),
    .I_4_2_1(op_I_4_2_1),
    .I_4_2_2(op_I_4_2_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_5_1_2(op_I_5_1_2),
    .I_5_2_0(op_I_5_2_0),
    .I_5_2_1(op_I_5_2_1),
    .I_5_2_2(op_I_5_2_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_6_1_2(op_I_6_1_2),
    .I_6_2_0(op_I_6_2_0),
    .I_6_2_1(op_I_6_2_1),
    .I_6_2_2(op_I_6_2_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_7_1_2(op_I_7_1_2),
    .I_7_2_0(op_I_7_2_0),
    .I_7_2_1(op_I_7_2_1),
    .I_7_2_2(op_I_7_2_2),
    .I_8_0_0(op_I_8_0_0),
    .I_8_0_1(op_I_8_0_1),
    .I_8_0_2(op_I_8_0_2),
    .I_8_1_0(op_I_8_1_0),
    .I_8_1_1(op_I_8_1_1),
    .I_8_1_2(op_I_8_1_2),
    .I_8_2_0(op_I_8_2_0),
    .I_8_2_1(op_I_8_2_1),
    .I_8_2_2(op_I_8_2_2),
    .I_9_0_0(op_I_9_0_0),
    .I_9_0_1(op_I_9_0_1),
    .I_9_0_2(op_I_9_0_2),
    .I_9_1_0(op_I_9_1_0),
    .I_9_1_1(op_I_9_1_1),
    .I_9_1_2(op_I_9_1_2),
    .I_9_2_0(op_I_9_2_0),
    .I_9_2_1(op_I_9_2_1),
    .I_9_2_2(op_I_9_2_2),
    .I_10_0_0(op_I_10_0_0),
    .I_10_0_1(op_I_10_0_1),
    .I_10_0_2(op_I_10_0_2),
    .I_10_1_0(op_I_10_1_0),
    .I_10_1_1(op_I_10_1_1),
    .I_10_1_2(op_I_10_1_2),
    .I_10_2_0(op_I_10_2_0),
    .I_10_2_1(op_I_10_2_1),
    .I_10_2_2(op_I_10_2_2),
    .I_11_0_0(op_I_11_0_0),
    .I_11_0_1(op_I_11_0_1),
    .I_11_0_2(op_I_11_0_2),
    .I_11_1_0(op_I_11_1_0),
    .I_11_1_1(op_I_11_1_1),
    .I_11_1_2(op_I_11_1_2),
    .I_11_2_0(op_I_11_2_0),
    .I_11_2_1(op_I_11_2_1),
    .I_11_2_2(op_I_11_2_2),
    .I_12_0_0(op_I_12_0_0),
    .I_12_0_1(op_I_12_0_1),
    .I_12_0_2(op_I_12_0_2),
    .I_12_1_0(op_I_12_1_0),
    .I_12_1_1(op_I_12_1_1),
    .I_12_1_2(op_I_12_1_2),
    .I_12_2_0(op_I_12_2_0),
    .I_12_2_1(op_I_12_2_1),
    .I_12_2_2(op_I_12_2_2),
    .I_13_0_0(op_I_13_0_0),
    .I_13_0_1(op_I_13_0_1),
    .I_13_0_2(op_I_13_0_2),
    .I_13_1_0(op_I_13_1_0),
    .I_13_1_1(op_I_13_1_1),
    .I_13_1_2(op_I_13_1_2),
    .I_13_2_0(op_I_13_2_0),
    .I_13_2_1(op_I_13_2_1),
    .I_13_2_2(op_I_13_2_2),
    .I_14_0_0(op_I_14_0_0),
    .I_14_0_1(op_I_14_0_1),
    .I_14_0_2(op_I_14_0_2),
    .I_14_1_0(op_I_14_1_0),
    .I_14_1_1(op_I_14_1_1),
    .I_14_1_2(op_I_14_1_2),
    .I_14_2_0(op_I_14_2_0),
    .I_14_2_1(op_I_14_2_1),
    .I_14_2_2(op_I_14_2_2),
    .I_15_0_0(op_I_15_0_0),
    .I_15_0_1(op_I_15_0_1),
    .I_15_0_2(op_I_15_0_2),
    .I_15_1_0(op_I_15_1_0),
    .I_15_1_1(op_I_15_1_1),
    .I_15_1_2(op_I_15_1_2),
    .I_15_2_0(op_I_15_2_0),
    .I_15_2_1(op_I_15_2_1),
    .I_15_2_2(op_I_15_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_1_0_0(op_O_1_0_0),
    .O_2_0_0(op_O_2_0_0),
    .O_3_0_0(op_O_3_0_0),
    .O_4_0_0(op_O_4_0_0),
    .O_5_0_0(op_O_5_0_0),
    .O_6_0_0(op_O_6_0_0),
    .O_7_0_0(op_O_7_0_0),
    .O_8_0_0(op_O_8_0_0),
    .O_9_0_0(op_O_9_0_0),
    .O_10_0_0(op_O_10_0_0),
    .O_11_0_0(op_O_11_0_0),
    .O_12_0_0(op_O_12_0_0),
    .O_13_0_0(op_O_13_0_0),
    .O_14_0_0(op_O_14_0_0),
    .O_15_0_0(op_O_15_0_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_8_0_0 = op_O_8_0_0; // @[MapT.scala 15:7]
  assign O_9_0_0 = op_O_9_0_0; // @[MapT.scala 15:7]
  assign O_10_0_0 = op_O_10_0_0; // @[MapT.scala 15:7]
  assign O_11_0_0 = op_O_11_0_0; // @[MapT.scala 15:7]
  assign O_12_0_0 = op_O_12_0_0; // @[MapT.scala 15:7]
  assign O_13_0_0 = op_O_13_0_0; // @[MapT.scala 15:7]
  assign O_14_0_0 = op_O_14_0_0; // @[MapT.scala 15:7]
  assign O_15_0_0 = op_O_15_0_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_4_1_2 = I_4_1_2; // @[MapT.scala 14:10]
  assign op_I_4_2_0 = I_4_2_0; // @[MapT.scala 14:10]
  assign op_I_4_2_1 = I_4_2_1; // @[MapT.scala 14:10]
  assign op_I_4_2_2 = I_4_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_5_1_2 = I_5_1_2; // @[MapT.scala 14:10]
  assign op_I_5_2_0 = I_5_2_0; // @[MapT.scala 14:10]
  assign op_I_5_2_1 = I_5_2_1; // @[MapT.scala 14:10]
  assign op_I_5_2_2 = I_5_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_6_1_2 = I_6_1_2; // @[MapT.scala 14:10]
  assign op_I_6_2_0 = I_6_2_0; // @[MapT.scala 14:10]
  assign op_I_6_2_1 = I_6_2_1; // @[MapT.scala 14:10]
  assign op_I_6_2_2 = I_6_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_7_1_2 = I_7_1_2; // @[MapT.scala 14:10]
  assign op_I_7_2_0 = I_7_2_0; // @[MapT.scala 14:10]
  assign op_I_7_2_1 = I_7_2_1; // @[MapT.scala 14:10]
  assign op_I_7_2_2 = I_7_2_2; // @[MapT.scala 14:10]
  assign op_I_8_0_0 = I_8_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1 = I_8_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_2 = I_8_0_2; // @[MapT.scala 14:10]
  assign op_I_8_1_0 = I_8_1_0; // @[MapT.scala 14:10]
  assign op_I_8_1_1 = I_8_1_1; // @[MapT.scala 14:10]
  assign op_I_8_1_2 = I_8_1_2; // @[MapT.scala 14:10]
  assign op_I_8_2_0 = I_8_2_0; // @[MapT.scala 14:10]
  assign op_I_8_2_1 = I_8_2_1; // @[MapT.scala 14:10]
  assign op_I_8_2_2 = I_8_2_2; // @[MapT.scala 14:10]
  assign op_I_9_0_0 = I_9_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1 = I_9_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_2 = I_9_0_2; // @[MapT.scala 14:10]
  assign op_I_9_1_0 = I_9_1_0; // @[MapT.scala 14:10]
  assign op_I_9_1_1 = I_9_1_1; // @[MapT.scala 14:10]
  assign op_I_9_1_2 = I_9_1_2; // @[MapT.scala 14:10]
  assign op_I_9_2_0 = I_9_2_0; // @[MapT.scala 14:10]
  assign op_I_9_2_1 = I_9_2_1; // @[MapT.scala 14:10]
  assign op_I_9_2_2 = I_9_2_2; // @[MapT.scala 14:10]
  assign op_I_10_0_0 = I_10_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1 = I_10_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_2 = I_10_0_2; // @[MapT.scala 14:10]
  assign op_I_10_1_0 = I_10_1_0; // @[MapT.scala 14:10]
  assign op_I_10_1_1 = I_10_1_1; // @[MapT.scala 14:10]
  assign op_I_10_1_2 = I_10_1_2; // @[MapT.scala 14:10]
  assign op_I_10_2_0 = I_10_2_0; // @[MapT.scala 14:10]
  assign op_I_10_2_1 = I_10_2_1; // @[MapT.scala 14:10]
  assign op_I_10_2_2 = I_10_2_2; // @[MapT.scala 14:10]
  assign op_I_11_0_0 = I_11_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1 = I_11_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_2 = I_11_0_2; // @[MapT.scala 14:10]
  assign op_I_11_1_0 = I_11_1_0; // @[MapT.scala 14:10]
  assign op_I_11_1_1 = I_11_1_1; // @[MapT.scala 14:10]
  assign op_I_11_1_2 = I_11_1_2; // @[MapT.scala 14:10]
  assign op_I_11_2_0 = I_11_2_0; // @[MapT.scala 14:10]
  assign op_I_11_2_1 = I_11_2_1; // @[MapT.scala 14:10]
  assign op_I_11_2_2 = I_11_2_2; // @[MapT.scala 14:10]
  assign op_I_12_0_0 = I_12_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1 = I_12_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_2 = I_12_0_2; // @[MapT.scala 14:10]
  assign op_I_12_1_0 = I_12_1_0; // @[MapT.scala 14:10]
  assign op_I_12_1_1 = I_12_1_1; // @[MapT.scala 14:10]
  assign op_I_12_1_2 = I_12_1_2; // @[MapT.scala 14:10]
  assign op_I_12_2_0 = I_12_2_0; // @[MapT.scala 14:10]
  assign op_I_12_2_1 = I_12_2_1; // @[MapT.scala 14:10]
  assign op_I_12_2_2 = I_12_2_2; // @[MapT.scala 14:10]
  assign op_I_13_0_0 = I_13_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1 = I_13_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_2 = I_13_0_2; // @[MapT.scala 14:10]
  assign op_I_13_1_0 = I_13_1_0; // @[MapT.scala 14:10]
  assign op_I_13_1_1 = I_13_1_1; // @[MapT.scala 14:10]
  assign op_I_13_1_2 = I_13_1_2; // @[MapT.scala 14:10]
  assign op_I_13_2_0 = I_13_2_0; // @[MapT.scala 14:10]
  assign op_I_13_2_1 = I_13_2_1; // @[MapT.scala 14:10]
  assign op_I_13_2_2 = I_13_2_2; // @[MapT.scala 14:10]
  assign op_I_14_0_0 = I_14_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1 = I_14_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_2 = I_14_0_2; // @[MapT.scala 14:10]
  assign op_I_14_1_0 = I_14_1_0; // @[MapT.scala 14:10]
  assign op_I_14_1_1 = I_14_1_1; // @[MapT.scala 14:10]
  assign op_I_14_1_2 = I_14_1_2; // @[MapT.scala 14:10]
  assign op_I_14_2_0 = I_14_2_0; // @[MapT.scala 14:10]
  assign op_I_14_2_1 = I_14_2_1; // @[MapT.scala 14:10]
  assign op_I_14_2_2 = I_14_2_2; // @[MapT.scala 14:10]
  assign op_I_15_0_0 = I_15_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1 = I_15_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_2 = I_15_0_2; // @[MapT.scala 14:10]
  assign op_I_15_1_0 = I_15_1_0; // @[MapT.scala 14:10]
  assign op_I_15_1_1 = I_15_1_1; // @[MapT.scala 14:10]
  assign op_I_15_1_2 = I_15_1_2; // @[MapT.scala 14:10]
  assign op_I_15_2_0 = I_15_2_0; // @[MapT.scala 14:10]
  assign op_I_15_2_1 = I_15_2_1; // @[MapT.scala 14:10]
  assign op_I_15_2_2 = I_15_2_2; // @[MapT.scala 14:10]
endmodule
module FIFO_1(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_1_0_0,
  input  [7:0] I_2_0_0,
  input  [7:0] I_3_0_0,
  input  [7:0] I_4_0_0,
  input  [7:0] I_5_0_0,
  input  [7:0] I_6_0_0,
  input  [7:0] I_7_0_0,
  input  [7:0] I_8_0_0,
  input  [7:0] I_9_0_0,
  input  [7:0] I_10_0_0,
  input  [7:0] I_11_0_0,
  input  [7:0] I_12_0_0,
  input  [7:0] I_13_0_0,
  input  [7:0] I_14_0_0,
  input  [7:0] I_15_0_0,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0,
  output [7:0] O_8_0_0,
  output [7:0] O_9_0_0,
  output [7:0] O_10_0_0,
  output [7:0] O_11_0_0,
  output [7:0] O_12_0_0,
  output [7:0] O_13_0_0,
  output [7:0] O_14_0_0,
  output [7:0] O_15_0_0
);
  reg [7:0] _T__0_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_0;
  wire [7:0] _T__0_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__0_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_1;
  wire [7:0] _T__0_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__0_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__0_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__0_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__0_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [1:0] _T__0_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [7:0] _T__1_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_4;
  wire [7:0] _T__1_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__1_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_5;
  wire [7:0] _T__1_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__1_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__1_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__1_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__1_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_6;
  reg [1:0] _T__1_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_7;
  reg [7:0] _T__2_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_8;
  wire [7:0] _T__2_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__2_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_9;
  wire [7:0] _T__2_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__2_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__2_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__2_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__2_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [1:0] _T__2_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [7:0] _T__3_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_12;
  wire [7:0] _T__3_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__3_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_13;
  wire [7:0] _T__3_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__3_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__3_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__3_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__3_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_14;
  reg [1:0] _T__3_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_15;
  reg [7:0] _T__4_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_16;
  wire [7:0] _T__4_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__4_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_17;
  wire [7:0] _T__4_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__4_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__4_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__4_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__4_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_18;
  reg [1:0] _T__4_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_19;
  reg [7:0] _T__5_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_20;
  wire [7:0] _T__5_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__5_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_21;
  wire [7:0] _T__5_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__5_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__5_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__5_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__5_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_22;
  reg [1:0] _T__5_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_23;
  reg [7:0] _T__6_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_24;
  wire [7:0] _T__6_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__6_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_25;
  wire [7:0] _T__6_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__6_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__6_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__6_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__6_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_26;
  reg [1:0] _T__6_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_27;
  reg [7:0] _T__7_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_28;
  wire [7:0] _T__7_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__7_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_29;
  wire [7:0] _T__7_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__7_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__7_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__7_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__7_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_30;
  reg [1:0] _T__7_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_31;
  reg [7:0] _T__8_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_32;
  wire [7:0] _T__8_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__8_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_33;
  wire [7:0] _T__8_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__8_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__8_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__8_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__8_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_34;
  reg [1:0] _T__8_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_35;
  reg [7:0] _T__9_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_36;
  wire [7:0] _T__9_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__9_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_37;
  wire [7:0] _T__9_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__9_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__9_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__9_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__9_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_38;
  reg [1:0] _T__9_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_39;
  reg [7:0] _T__10_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_40;
  wire [7:0] _T__10_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__10_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_41;
  wire [7:0] _T__10_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__10_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__10_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__10_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__10_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_42;
  reg [1:0] _T__10_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_43;
  reg [7:0] _T__11_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_44;
  wire [7:0] _T__11_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__11_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_45;
  wire [7:0] _T__11_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__11_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__11_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__11_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__11_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_46;
  reg [1:0] _T__11_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_47;
  reg [7:0] _T__12_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_48;
  wire [7:0] _T__12_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__12_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_49;
  wire [7:0] _T__12_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__12_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__12_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__12_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__12_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_50;
  reg [1:0] _T__12_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_51;
  reg [7:0] _T__13_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_52;
  wire [7:0] _T__13_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__13_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_53;
  wire [7:0] _T__13_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__13_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__13_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__13_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__13_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_54;
  reg [1:0] _T__13_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_55;
  reg [7:0] _T__14_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_56;
  wire [7:0] _T__14_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__14_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_57;
  wire [7:0] _T__14_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__14_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__14_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__14_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__14_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_58;
  reg [1:0] _T__14_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_59;
  reg [7:0] _T__15_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_60;
  wire [7:0] _T__15_0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__15_0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_61;
  wire [7:0] _T__15_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__15_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__15_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__15_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__15_0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_62;
  reg [1:0] _T__15_0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_63;
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_64;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_65;
  reg [1:0] value_2; // @[Counter.scala 29:33]
  reg [31:0] _RAND_66;
  wire  _T_1; // @[FIFO.scala 33:46]
  wire  _T_2; // @[Counter.scala 37:24]
  wire [1:0] _T_4; // @[Counter.scala 38:22]
  wire  _T_6; // @[FIFO.scala 38:39]
  wire  _T_7; // @[FIFO.scala 39:15]
  wire  _T_8; // @[FIFO.scala 39:15]
  wire [1:0] _T_11; // @[Counter.scala 38:22]
  wire  _T_12; // @[FIFO.scala 42:39]
  wire  _T_18; // @[Counter.scala 37:24]
  wire [1:0] _T_20; // @[Counter.scala 38:22]
  wire  _GEN_8; // @[FIFO.scala 42:57]
  wire  _GEN_70; // @[FIFO.scala 39:15]
  assign _T__0_0_0__T_17_addr = _T__0_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__0_0_0__T_17_data = _T__0_0_0[_T__0_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__0_0_0__T_17_data = _T__0_0_0__T_17_addr >= 2'h3 ? _RAND_1[7:0] : _T__0_0_0[_T__0_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__0_0_0__T_5_data = I_0_0_0;
  assign _T__0_0_0__T_5_addr = value_2;
  assign _T__0_0_0__T_5_mask = 1'h1;
  assign _T__0_0_0__T_5_en = valid_up;
  assign _T__1_0_0__T_17_addr = _T__1_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__1_0_0__T_17_data = _T__1_0_0[_T__1_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__1_0_0__T_17_data = _T__1_0_0__T_17_addr >= 2'h3 ? _RAND_5[7:0] : _T__1_0_0[_T__1_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__1_0_0__T_5_data = I_1_0_0;
  assign _T__1_0_0__T_5_addr = value_2;
  assign _T__1_0_0__T_5_mask = 1'h1;
  assign _T__1_0_0__T_5_en = valid_up;
  assign _T__2_0_0__T_17_addr = _T__2_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__2_0_0__T_17_data = _T__2_0_0[_T__2_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__2_0_0__T_17_data = _T__2_0_0__T_17_addr >= 2'h3 ? _RAND_9[7:0] : _T__2_0_0[_T__2_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__2_0_0__T_5_data = I_2_0_0;
  assign _T__2_0_0__T_5_addr = value_2;
  assign _T__2_0_0__T_5_mask = 1'h1;
  assign _T__2_0_0__T_5_en = valid_up;
  assign _T__3_0_0__T_17_addr = _T__3_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__3_0_0__T_17_data = _T__3_0_0[_T__3_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__3_0_0__T_17_data = _T__3_0_0__T_17_addr >= 2'h3 ? _RAND_13[7:0] : _T__3_0_0[_T__3_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__3_0_0__T_5_data = I_3_0_0;
  assign _T__3_0_0__T_5_addr = value_2;
  assign _T__3_0_0__T_5_mask = 1'h1;
  assign _T__3_0_0__T_5_en = valid_up;
  assign _T__4_0_0__T_17_addr = _T__4_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__4_0_0__T_17_data = _T__4_0_0[_T__4_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__4_0_0__T_17_data = _T__4_0_0__T_17_addr >= 2'h3 ? _RAND_17[7:0] : _T__4_0_0[_T__4_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__4_0_0__T_5_data = I_4_0_0;
  assign _T__4_0_0__T_5_addr = value_2;
  assign _T__4_0_0__T_5_mask = 1'h1;
  assign _T__4_0_0__T_5_en = valid_up;
  assign _T__5_0_0__T_17_addr = _T__5_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__5_0_0__T_17_data = _T__5_0_0[_T__5_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__5_0_0__T_17_data = _T__5_0_0__T_17_addr >= 2'h3 ? _RAND_21[7:0] : _T__5_0_0[_T__5_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__5_0_0__T_5_data = I_5_0_0;
  assign _T__5_0_0__T_5_addr = value_2;
  assign _T__5_0_0__T_5_mask = 1'h1;
  assign _T__5_0_0__T_5_en = valid_up;
  assign _T__6_0_0__T_17_addr = _T__6_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__6_0_0__T_17_data = _T__6_0_0[_T__6_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__6_0_0__T_17_data = _T__6_0_0__T_17_addr >= 2'h3 ? _RAND_25[7:0] : _T__6_0_0[_T__6_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__6_0_0__T_5_data = I_6_0_0;
  assign _T__6_0_0__T_5_addr = value_2;
  assign _T__6_0_0__T_5_mask = 1'h1;
  assign _T__6_0_0__T_5_en = valid_up;
  assign _T__7_0_0__T_17_addr = _T__7_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__7_0_0__T_17_data = _T__7_0_0[_T__7_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__7_0_0__T_17_data = _T__7_0_0__T_17_addr >= 2'h3 ? _RAND_29[7:0] : _T__7_0_0[_T__7_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__7_0_0__T_5_data = I_7_0_0;
  assign _T__7_0_0__T_5_addr = value_2;
  assign _T__7_0_0__T_5_mask = 1'h1;
  assign _T__7_0_0__T_5_en = valid_up;
  assign _T__8_0_0__T_17_addr = _T__8_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__8_0_0__T_17_data = _T__8_0_0[_T__8_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__8_0_0__T_17_data = _T__8_0_0__T_17_addr >= 2'h3 ? _RAND_33[7:0] : _T__8_0_0[_T__8_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__8_0_0__T_5_data = I_8_0_0;
  assign _T__8_0_0__T_5_addr = value_2;
  assign _T__8_0_0__T_5_mask = 1'h1;
  assign _T__8_0_0__T_5_en = valid_up;
  assign _T__9_0_0__T_17_addr = _T__9_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__9_0_0__T_17_data = _T__9_0_0[_T__9_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__9_0_0__T_17_data = _T__9_0_0__T_17_addr >= 2'h3 ? _RAND_37[7:0] : _T__9_0_0[_T__9_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__9_0_0__T_5_data = I_9_0_0;
  assign _T__9_0_0__T_5_addr = value_2;
  assign _T__9_0_0__T_5_mask = 1'h1;
  assign _T__9_0_0__T_5_en = valid_up;
  assign _T__10_0_0__T_17_addr = _T__10_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__10_0_0__T_17_data = _T__10_0_0[_T__10_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__10_0_0__T_17_data = _T__10_0_0__T_17_addr >= 2'h3 ? _RAND_41[7:0] : _T__10_0_0[_T__10_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__10_0_0__T_5_data = I_10_0_0;
  assign _T__10_0_0__T_5_addr = value_2;
  assign _T__10_0_0__T_5_mask = 1'h1;
  assign _T__10_0_0__T_5_en = valid_up;
  assign _T__11_0_0__T_17_addr = _T__11_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__11_0_0__T_17_data = _T__11_0_0[_T__11_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__11_0_0__T_17_data = _T__11_0_0__T_17_addr >= 2'h3 ? _RAND_45[7:0] : _T__11_0_0[_T__11_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__11_0_0__T_5_data = I_11_0_0;
  assign _T__11_0_0__T_5_addr = value_2;
  assign _T__11_0_0__T_5_mask = 1'h1;
  assign _T__11_0_0__T_5_en = valid_up;
  assign _T__12_0_0__T_17_addr = _T__12_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__12_0_0__T_17_data = _T__12_0_0[_T__12_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__12_0_0__T_17_data = _T__12_0_0__T_17_addr >= 2'h3 ? _RAND_49[7:0] : _T__12_0_0[_T__12_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__12_0_0__T_5_data = I_12_0_0;
  assign _T__12_0_0__T_5_addr = value_2;
  assign _T__12_0_0__T_5_mask = 1'h1;
  assign _T__12_0_0__T_5_en = valid_up;
  assign _T__13_0_0__T_17_addr = _T__13_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__13_0_0__T_17_data = _T__13_0_0[_T__13_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__13_0_0__T_17_data = _T__13_0_0__T_17_addr >= 2'h3 ? _RAND_53[7:0] : _T__13_0_0[_T__13_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__13_0_0__T_5_data = I_13_0_0;
  assign _T__13_0_0__T_5_addr = value_2;
  assign _T__13_0_0__T_5_mask = 1'h1;
  assign _T__13_0_0__T_5_en = valid_up;
  assign _T__14_0_0__T_17_addr = _T__14_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__14_0_0__T_17_data = _T__14_0_0[_T__14_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__14_0_0__T_17_data = _T__14_0_0__T_17_addr >= 2'h3 ? _RAND_57[7:0] : _T__14_0_0[_T__14_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__14_0_0__T_5_data = I_14_0_0;
  assign _T__14_0_0__T_5_addr = value_2;
  assign _T__14_0_0__T_5_mask = 1'h1;
  assign _T__14_0_0__T_5_en = valid_up;
  assign _T__15_0_0__T_17_addr = _T__15_0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__15_0_0__T_17_data = _T__15_0_0[_T__15_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__15_0_0__T_17_data = _T__15_0_0__T_17_addr >= 2'h3 ? _RAND_61[7:0] : _T__15_0_0[_T__15_0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__15_0_0__T_5_data = I_15_0_0;
  assign _T__15_0_0__T_5_addr = value_2;
  assign _T__15_0_0__T_5_mask = 1'h1;
  assign _T__15_0_0__T_5_en = valid_up;
  assign _T_1 = value == 2'h2; // @[FIFO.scala 33:46]
  assign _T_2 = value_2 == 2'h2; // @[Counter.scala 37:24]
  assign _T_4 = value_2 + 2'h1; // @[Counter.scala 38:22]
  assign _T_6 = value < 2'h2; // @[FIFO.scala 38:39]
  assign _T_7 = $unsigned(reset); // @[FIFO.scala 39:15]
  assign _T_8 = _T_7 == 1'h0; // @[FIFO.scala 39:15]
  assign _T_11 = value + 2'h1; // @[Counter.scala 38:22]
  assign _T_12 = value >= 2'h1; // @[FIFO.scala 42:39]
  assign _T_18 = value_1 == 2'h2; // @[Counter.scala 37:24]
  assign _T_20 = value_1 + 2'h1; // @[Counter.scala 38:22]
  assign _GEN_8 = _T_12 & _T_12; // @[FIFO.scala 42:57]
  assign valid_down = value == 2'h2; // @[FIFO.scala 33:16]
  assign O_0_0_0 = _T__0_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_1_0_0 = _T__1_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_2_0_0 = _T__2_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_3_0_0 = _T__3_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_4_0_0 = _T__4_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_5_0_0 = _T__5_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_6_0_0 = _T__6_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_7_0_0 = _T__7_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_8_0_0 = _T__8_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_9_0_0 = _T__9_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_10_0_0 = _T__10_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_11_0_0 = _T__11_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_12_0_0 = _T__12_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_13_0_0 = _T__13_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_14_0_0 = _T__14_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_15_0_0 = _T__15_0_0__T_17_data; // @[FIFO.scala 43:11]
  assign _GEN_70 = valid_up & _T_6; // @[FIFO.scala 39:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__0_0_0[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__0_0_0__T_17_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__0_0_0__T_17_addr_pipe_0 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__1_0_0[initvar] = _RAND_4[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__1_0_0__T_17_en_pipe_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__1_0_0__T_17_addr_pipe_0 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__2_0_0[initvar] = _RAND_8[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__2_0_0__T_17_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__2_0_0__T_17_addr_pipe_0 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__3_0_0[initvar] = _RAND_12[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__3_0_0__T_17_en_pipe_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__3_0_0__T_17_addr_pipe_0 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__4_0_0[initvar] = _RAND_16[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_17 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T__4_0_0__T_17_en_pipe_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T__4_0_0__T_17_addr_pipe_0 = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__5_0_0[initvar] = _RAND_20[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_21 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T__5_0_0__T_17_en_pipe_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T__5_0_0__T_17_addr_pipe_0 = _RAND_23[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__6_0_0[initvar] = _RAND_24[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_25 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T__6_0_0__T_17_en_pipe_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T__6_0_0__T_17_addr_pipe_0 = _RAND_27[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__7_0_0[initvar] = _RAND_28[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_29 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T__7_0_0__T_17_en_pipe_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T__7_0_0__T_17_addr_pipe_0 = _RAND_31[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__8_0_0[initvar] = _RAND_32[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_33 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T__8_0_0__T_17_en_pipe_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T__8_0_0__T_17_addr_pipe_0 = _RAND_35[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__9_0_0[initvar] = _RAND_36[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_37 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T__9_0_0__T_17_en_pipe_0 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T__9_0_0__T_17_addr_pipe_0 = _RAND_39[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__10_0_0[initvar] = _RAND_40[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_41 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T__10_0_0__T_17_en_pipe_0 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T__10_0_0__T_17_addr_pipe_0 = _RAND_43[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__11_0_0[initvar] = _RAND_44[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_45 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T__11_0_0__T_17_en_pipe_0 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T__11_0_0__T_17_addr_pipe_0 = _RAND_47[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__12_0_0[initvar] = _RAND_48[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_49 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T__12_0_0__T_17_en_pipe_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T__12_0_0__T_17_addr_pipe_0 = _RAND_51[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__13_0_0[initvar] = _RAND_52[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_53 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T__13_0_0__T_17_en_pipe_0 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T__13_0_0__T_17_addr_pipe_0 = _RAND_55[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__14_0_0[initvar] = _RAND_56[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_57 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T__14_0_0__T_17_en_pipe_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T__14_0_0__T_17_addr_pipe_0 = _RAND_59[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__15_0_0[initvar] = _RAND_60[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_61 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T__15_0_0__T_17_en_pipe_0 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T__15_0_0__T_17_addr_pipe_0 = _RAND_63[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  value = _RAND_64[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  value_1 = _RAND_65[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  value_2 = _RAND_66[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__0_0_0__T_5_en & _T__0_0_0__T_5_mask) begin
      _T__0_0_0[_T__0_0_0__T_5_addr] <= _T__0_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__0_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__0_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__1_0_0__T_5_en & _T__1_0_0__T_5_mask) begin
      _T__1_0_0[_T__1_0_0__T_5_addr] <= _T__1_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__1_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__1_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__2_0_0__T_5_en & _T__2_0_0__T_5_mask) begin
      _T__2_0_0[_T__2_0_0__T_5_addr] <= _T__2_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__2_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__2_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__3_0_0__T_5_en & _T__3_0_0__T_5_mask) begin
      _T__3_0_0[_T__3_0_0__T_5_addr] <= _T__3_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__3_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__3_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__4_0_0__T_5_en & _T__4_0_0__T_5_mask) begin
      _T__4_0_0[_T__4_0_0__T_5_addr] <= _T__4_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__4_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__4_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__5_0_0__T_5_en & _T__5_0_0__T_5_mask) begin
      _T__5_0_0[_T__5_0_0__T_5_addr] <= _T__5_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__5_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__5_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__6_0_0__T_5_en & _T__6_0_0__T_5_mask) begin
      _T__6_0_0[_T__6_0_0__T_5_addr] <= _T__6_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__6_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__6_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__7_0_0__T_5_en & _T__7_0_0__T_5_mask) begin
      _T__7_0_0[_T__7_0_0__T_5_addr] <= _T__7_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__7_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__7_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__8_0_0__T_5_en & _T__8_0_0__T_5_mask) begin
      _T__8_0_0[_T__8_0_0__T_5_addr] <= _T__8_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__8_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__8_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__9_0_0__T_5_en & _T__9_0_0__T_5_mask) begin
      _T__9_0_0[_T__9_0_0__T_5_addr] <= _T__9_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__9_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__9_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__10_0_0__T_5_en & _T__10_0_0__T_5_mask) begin
      _T__10_0_0[_T__10_0_0__T_5_addr] <= _T__10_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__10_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__10_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__11_0_0__T_5_en & _T__11_0_0__T_5_mask) begin
      _T__11_0_0[_T__11_0_0__T_5_addr] <= _T__11_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__11_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__11_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__12_0_0__T_5_en & _T__12_0_0__T_5_mask) begin
      _T__12_0_0[_T__12_0_0__T_5_addr] <= _T__12_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__12_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__12_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__13_0_0__T_5_en & _T__13_0_0__T_5_mask) begin
      _T__13_0_0[_T__13_0_0__T_5_addr] <= _T__13_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__13_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__13_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__14_0_0__T_5_en & _T__14_0_0__T_5_mask) begin
      _T__14_0_0[_T__14_0_0__T_5_addr] <= _T__14_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__14_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__14_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__15_0_0__T_5_en & _T__15_0_0__T_5_mask) begin
      _T__15_0_0[_T__15_0_0__T_5_addr] <= _T__15_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__15_0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__15_0_0__T_17_addr_pipe_0 <= value_1;
    end
    if (reset) begin
      value <= 2'h0;
    end else if (valid_up) begin
      if (_T_6) begin
        if (_T_1) begin
          value <= 2'h0;
        end else begin
          value <= _T_11;
        end
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (valid_up) begin
      if (_T_12) begin
        if (_T_18) begin
          value_1 <= 2'h0;
        end else begin
          value_1 <= _T_20;
        end
      end
    end
    if (reset) begin
      value_2 <= 2'h0;
    end else if (valid_up) begin
      if (_T_2) begin
        value_2 <= 2'h0;
      end else begin
        value_2 <= _T_4;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_70 & _T_8) begin
          $fwrite(32'h80000002,"idc inc\n"); // @[FIFO.scala 39:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module FIFO_2(
  input        clock,
  input        valid_up,
  output       valid_down,
  input  [7:0] I,
  output [7:0] O
);
  reg [7:0] _T; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_1;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O = _T; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= I;
    _T_1 <= valid_up;
  end
endmodule
module InitialDelayCounter_2(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [2:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [2:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 3'h4; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 3'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 3'h4; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 3'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Sub(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 80:14]
  assign O = I_t0b - I_t1b; // @[Arithmetic.scala 79:5]
endmodule
module Abs(
  input        clock,
  input        valid_up,
  output       valid_down,
  input  [7:0] I,
  output [7:0] O
);
  reg [7:0] out_reg; // @[Arithmetic.scala 14:20]
  reg [31:0] _RAND_0;
  wire [7:0] _T; // @[Arithmetic.scala 15:16]
  wire  _T_1; // @[Arithmetic.scala 15:19]
  wire [7:0] _T_3; // @[Arithmetic.scala 15:43]
  reg  _T_4; // @[Arithmetic.scala 17:24]
  reg [31:0] _RAND_1;
  assign _T = $signed(I); // @[Arithmetic.scala 15:16]
  assign _T_1 = $signed(_T) < $signed(8'sh0); // @[Arithmetic.scala 15:19]
  assign _T_3 = 8'h0 - I; // @[Arithmetic.scala 15:43]
  assign valid_down = _T_4; // @[Arithmetic.scala 17:14]
  assign O = out_reg; // @[Arithmetic.scala 16:5]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_reg = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_4 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_1) begin
      out_reg <= _T_3;
    end else begin
      out_reg <= I;
    end
    _T_4 <= valid_up;
  end
endmodule
module Lt(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  wire  _T; // @[Arithmetic.scala 184:23]
  assign _T = I_t0b < I_t1b; // @[Arithmetic.scala 184:23]
  assign valid_down = valid_up; // @[Arithmetic.scala 185:14]
  assign O = {{7'd0}, _T}; // @[Arithmetic.scala 184:5]
endmodule
module FIFO_3(
  input        clock,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O_t0b,
  output [7:0] O_t1b
);
  reg [7:0] _T_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [7:0] _T_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_2;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_t0b = _T_t0b; // @[FIFO.scala 14:7]
  assign O_t1b = _T_t1b; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_t0b = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_t1b = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_t0b <= I_t0b;
    _T_t1b <= I_t1b;
    _T_1 <= valid_up;
  end
endmodule
module AtomTuple_5(
  input        valid_up,
  output       valid_down,
  input        I0,
  input  [7:0] I1_t0b,
  input  [7:0] I1_t1b,
  output       O_t0b,
  output [7:0] O_t1b_t0b,
  output [7:0] O_t1b_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b_t0b = I1_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t1b = I1_t1b; // @[Tuple.scala 50:9]
endmodule
module If(
  input        valid_up,
  output       valid_down,
  input        I_t0b,
  input  [7:0] I_t1b_t0b,
  input  [7:0] I_t1b_t1b,
  output [7:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 231:14]
  assign O = I_t0b ? I_t1b_t0b : I_t1b_t1b; // @[Arithmetic.scala 229:9 Arithmetic.scala 230:20]
endmodule
module Add(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 59:14]
  assign O = I_t0b + I_t1b; // @[Arithmetic.scala 58:5]
endmodule
module Module_1(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O
);
  wire  n214_clock; // @[Top.scala 45:22]
  wire  n214_valid_up; // @[Top.scala 45:22]
  wire  n214_valid_down; // @[Top.scala 45:22]
  wire [7:0] n214_I; // @[Top.scala 45:22]
  wire [7:0] n214_O; // @[Top.scala 45:22]
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n198_valid_up; // @[Top.scala 49:22]
  wire  n198_valid_down; // @[Top.scala 49:22]
  wire [7:0] n198_I0; // @[Top.scala 49:22]
  wire [7:0] n198_I1; // @[Top.scala 49:22]
  wire [7:0] n198_O_t0b; // @[Top.scala 49:22]
  wire [7:0] n198_O_t1b; // @[Top.scala 49:22]
  wire  n199_valid_up; // @[Top.scala 53:22]
  wire  n199_valid_down; // @[Top.scala 53:22]
  wire [7:0] n199_I_t0b; // @[Top.scala 53:22]
  wire [7:0] n199_I_t1b; // @[Top.scala 53:22]
  wire [7:0] n199_O; // @[Top.scala 53:22]
  wire  n200_clock; // @[Top.scala 56:22]
  wire  n200_valid_up; // @[Top.scala 56:22]
  wire  n200_valid_down; // @[Top.scala 56:22]
  wire [7:0] n200_I; // @[Top.scala 56:22]
  wire [7:0] n200_O; // @[Top.scala 56:22]
  wire  n202_valid_up; // @[Top.scala 59:22]
  wire  n202_valid_down; // @[Top.scala 59:22]
  wire [7:0] n202_I0; // @[Top.scala 59:22]
  wire [7:0] n202_I1; // @[Top.scala 59:22]
  wire [7:0] n202_O_t0b; // @[Top.scala 59:22]
  wire [7:0] n202_O_t1b; // @[Top.scala 59:22]
  wire  n203_valid_up; // @[Top.scala 63:22]
  wire  n203_valid_down; // @[Top.scala 63:22]
  wire [7:0] n203_I_t0b; // @[Top.scala 63:22]
  wire [7:0] n203_I_t1b; // @[Top.scala 63:22]
  wire [7:0] n203_O; // @[Top.scala 63:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n206_valid_up; // @[Top.scala 67:22]
  wire  n206_valid_down; // @[Top.scala 67:22]
  wire [7:0] n206_I0; // @[Top.scala 67:22]
  wire [7:0] n206_I1; // @[Top.scala 67:22]
  wire [7:0] n206_O_t0b; // @[Top.scala 67:22]
  wire [7:0] n206_O_t1b; // @[Top.scala 67:22]
  wire  n207_clock; // @[Top.scala 71:22]
  wire  n207_valid_up; // @[Top.scala 71:22]
  wire  n207_valid_down; // @[Top.scala 71:22]
  wire [7:0] n207_I_t0b; // @[Top.scala 71:22]
  wire [7:0] n207_I_t1b; // @[Top.scala 71:22]
  wire [7:0] n207_O_t0b; // @[Top.scala 71:22]
  wire [7:0] n207_O_t1b; // @[Top.scala 71:22]
  wire  n208_valid_up; // @[Top.scala 74:22]
  wire  n208_valid_down; // @[Top.scala 74:22]
  wire  n208_I0; // @[Top.scala 74:22]
  wire [7:0] n208_I1_t0b; // @[Top.scala 74:22]
  wire [7:0] n208_I1_t1b; // @[Top.scala 74:22]
  wire  n208_O_t0b; // @[Top.scala 74:22]
  wire [7:0] n208_O_t1b_t0b; // @[Top.scala 74:22]
  wire [7:0] n208_O_t1b_t1b; // @[Top.scala 74:22]
  wire  n209_valid_up; // @[Top.scala 78:22]
  wire  n209_valid_down; // @[Top.scala 78:22]
  wire  n209_I_t0b; // @[Top.scala 78:22]
  wire [7:0] n209_I_t1b_t0b; // @[Top.scala 78:22]
  wire [7:0] n209_I_t1b_t1b; // @[Top.scala 78:22]
  wire [7:0] n209_O; // @[Top.scala 78:22]
  wire  InitialDelayCounter_2_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_2_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_2_valid_down; // @[Const.scala 11:33]
  wire  n212_valid_up; // @[Top.scala 82:22]
  wire  n212_valid_down; // @[Top.scala 82:22]
  wire [7:0] n212_I0; // @[Top.scala 82:22]
  wire [7:0] n212_I1; // @[Top.scala 82:22]
  wire [7:0] n212_O_t0b; // @[Top.scala 82:22]
  wire [7:0] n212_O_t1b; // @[Top.scala 82:22]
  wire  n213_valid_up; // @[Top.scala 86:22]
  wire  n213_valid_down; // @[Top.scala 86:22]
  wire [7:0] n213_I_t0b; // @[Top.scala 86:22]
  wire [7:0] n213_I_t1b; // @[Top.scala 86:22]
  wire [7:0] n213_O; // @[Top.scala 86:22]
  wire  n215_valid_up; // @[Top.scala 89:22]
  wire  n215_valid_down; // @[Top.scala 89:22]
  wire [7:0] n215_I0; // @[Top.scala 89:22]
  wire [7:0] n215_I1; // @[Top.scala 89:22]
  wire [7:0] n215_O_t0b; // @[Top.scala 89:22]
  wire [7:0] n215_O_t1b; // @[Top.scala 89:22]
  wire  n216_valid_up; // @[Top.scala 93:22]
  wire  n216_valid_down; // @[Top.scala 93:22]
  wire [7:0] n216_I_t0b; // @[Top.scala 93:22]
  wire [7:0] n216_I_t1b; // @[Top.scala 93:22]
  wire [7:0] n216_O; // @[Top.scala 93:22]
  FIFO_2 n214 ( // @[Top.scala 45:22]
    .clock(n214_clock),
    .valid_up(n214_valid_up),
    .valid_down(n214_valid_down),
    .I(n214_I),
    .O(n214_O)
  );
  InitialDelayCounter_2 InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  AtomTuple n198 ( // @[Top.scala 49:22]
    .valid_up(n198_valid_up),
    .valid_down(n198_valid_down),
    .I0(n198_I0),
    .I1(n198_I1),
    .O_t0b(n198_O_t0b),
    .O_t1b(n198_O_t1b)
  );
  Sub n199 ( // @[Top.scala 53:22]
    .valid_up(n199_valid_up),
    .valid_down(n199_valid_down),
    .I_t0b(n199_I_t0b),
    .I_t1b(n199_I_t1b),
    .O(n199_O)
  );
  Abs n200 ( // @[Top.scala 56:22]
    .clock(n200_clock),
    .valid_up(n200_valid_up),
    .valid_down(n200_valid_down),
    .I(n200_I),
    .O(n200_O)
  );
  AtomTuple n202 ( // @[Top.scala 59:22]
    .valid_up(n202_valid_up),
    .valid_down(n202_valid_down),
    .I0(n202_I0),
    .I1(n202_I1),
    .O_t0b(n202_O_t0b),
    .O_t1b(n202_O_t1b)
  );
  Lt n203 ( // @[Top.scala 63:22]
    .valid_up(n203_valid_up),
    .valid_down(n203_valid_down),
    .I_t0b(n203_I_t0b),
    .I_t1b(n203_I_t1b),
    .O(n203_O)
  );
  InitialDelayCounter_1 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  AtomTuple n206 ( // @[Top.scala 67:22]
    .valid_up(n206_valid_up),
    .valid_down(n206_valid_down),
    .I0(n206_I0),
    .I1(n206_I1),
    .O_t0b(n206_O_t0b),
    .O_t1b(n206_O_t1b)
  );
  FIFO_3 n207 ( // @[Top.scala 71:22]
    .clock(n207_clock),
    .valid_up(n207_valid_up),
    .valid_down(n207_valid_down),
    .I_t0b(n207_I_t0b),
    .I_t1b(n207_I_t1b),
    .O_t0b(n207_O_t0b),
    .O_t1b(n207_O_t1b)
  );
  AtomTuple_5 n208 ( // @[Top.scala 74:22]
    .valid_up(n208_valid_up),
    .valid_down(n208_valid_down),
    .I0(n208_I0),
    .I1_t0b(n208_I1_t0b),
    .I1_t1b(n208_I1_t1b),
    .O_t0b(n208_O_t0b),
    .O_t1b_t0b(n208_O_t1b_t0b),
    .O_t1b_t1b(n208_O_t1b_t1b)
  );
  If n209 ( // @[Top.scala 78:22]
    .valid_up(n209_valid_up),
    .valid_down(n209_valid_down),
    .I_t0b(n209_I_t0b),
    .I_t1b_t0b(n209_I_t1b_t0b),
    .I_t1b_t1b(n209_I_t1b_t1b),
    .O(n209_O)
  );
  InitialDelayCounter_2 InitialDelayCounter_2 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_2_clock),
    .reset(InitialDelayCounter_2_reset),
    .valid_down(InitialDelayCounter_2_valid_down)
  );
  AtomTuple n212 ( // @[Top.scala 82:22]
    .valid_up(n212_valid_up),
    .valid_down(n212_valid_down),
    .I0(n212_I0),
    .I1(n212_I1),
    .O_t0b(n212_O_t0b),
    .O_t1b(n212_O_t1b)
  );
  RShift n213 ( // @[Top.scala 86:22]
    .valid_up(n213_valid_up),
    .valid_down(n213_valid_down),
    .I_t0b(n213_I_t0b),
    .I_t1b(n213_I_t1b),
    .O(n213_O)
  );
  AtomTuple n215 ( // @[Top.scala 89:22]
    .valid_up(n215_valid_up),
    .valid_down(n215_valid_down),
    .I0(n215_I0),
    .I1(n215_I1),
    .O_t0b(n215_O_t0b),
    .O_t1b(n215_O_t1b)
  );
  Add n216 ( // @[Top.scala 93:22]
    .valid_up(n216_valid_up),
    .valid_down(n216_valid_down),
    .I_t0b(n216_I_t0b),
    .I_t1b(n216_I_t1b),
    .O(n216_O)
  );
  assign valid_down = n216_valid_down; // @[Top.scala 97:16]
  assign O = n216_O; // @[Top.scala 96:7]
  assign n214_clock = clock;
  assign n214_valid_up = valid_up; // @[Top.scala 47:19]
  assign n214_I = I1; // @[Top.scala 46:12]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n198_valid_up = valid_up & valid_up; // @[Top.scala 52:19]
  assign n198_I0 = I1; // @[Top.scala 50:13]
  assign n198_I1 = I0; // @[Top.scala 51:13]
  assign n199_valid_up = n198_valid_down; // @[Top.scala 55:19]
  assign n199_I_t0b = n198_O_t0b; // @[Top.scala 54:12]
  assign n199_I_t1b = n198_O_t1b; // @[Top.scala 54:12]
  assign n200_clock = clock;
  assign n200_valid_up = n199_valid_down; // @[Top.scala 58:19]
  assign n200_I = n199_O; // @[Top.scala 57:12]
  assign n202_valid_up = InitialDelayCounter_valid_down & n200_valid_down; // @[Top.scala 62:19]
  assign n202_I0 = 8'hf; // @[Top.scala 60:13]
  assign n202_I1 = n200_O; // @[Top.scala 61:13]
  assign n203_valid_up = n202_valid_down; // @[Top.scala 65:19]
  assign n203_I_t0b = n202_O_t0b; // @[Top.scala 64:12]
  assign n203_I_t1b = n202_O_t1b; // @[Top.scala 64:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n206_valid_up = n199_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 70:19]
  assign n206_I0 = n199_O; // @[Top.scala 68:13]
  assign n206_I1 = 8'h0; // @[Top.scala 69:13]
  assign n207_clock = clock;
  assign n207_valid_up = n206_valid_down; // @[Top.scala 73:19]
  assign n207_I_t0b = n206_O_t0b; // @[Top.scala 72:12]
  assign n207_I_t1b = n206_O_t1b; // @[Top.scala 72:12]
  assign n208_valid_up = n203_valid_down & n207_valid_down; // @[Top.scala 77:19]
  assign n208_I0 = n203_O[0]; // @[Top.scala 75:13]
  assign n208_I1_t0b = n207_O_t0b; // @[Top.scala 76:13]
  assign n208_I1_t1b = n207_O_t1b; // @[Top.scala 76:13]
  assign n209_valid_up = n208_valid_down; // @[Top.scala 80:19]
  assign n209_I_t0b = n208_O_t0b; // @[Top.scala 79:12]
  assign n209_I_t1b_t0b = n208_O_t1b_t0b; // @[Top.scala 79:12]
  assign n209_I_t1b_t1b = n208_O_t1b_t1b; // @[Top.scala 79:12]
  assign InitialDelayCounter_2_clock = clock;
  assign InitialDelayCounter_2_reset = reset;
  assign n212_valid_up = n209_valid_down & InitialDelayCounter_2_valid_down; // @[Top.scala 85:19]
  assign n212_I0 = n209_O; // @[Top.scala 83:13]
  assign n212_I1 = 8'h2; // @[Top.scala 84:13]
  assign n213_valid_up = n212_valid_down; // @[Top.scala 88:19]
  assign n213_I_t0b = n212_O_t0b; // @[Top.scala 87:12]
  assign n213_I_t1b = n212_O_t1b; // @[Top.scala 87:12]
  assign n215_valid_up = n214_valid_down & n213_valid_down; // @[Top.scala 92:19]
  assign n215_I0 = n214_O; // @[Top.scala 90:13]
  assign n215_I1 = n213_O; // @[Top.scala 91:13]
  assign n216_valid_up = n215_valid_down; // @[Top.scala 95:19]
  assign n216_I_t0b = n215_O_t0b; // @[Top.scala 94:12]
  assign n216_I_t1b = n215_O_t1b; // @[Top.scala 94:12]
endmodule
module Map2S_26(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I1_0,
  output [7:0] O_0
);
  wire  fst_op_clock; // @[Map2S.scala 9:22]
  wire  fst_op_reset; // @[Map2S.scala 9:22]
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O; // @[Map2S.scala 9:22]
  Module_1 fst_op ( // @[Map2S.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0 = fst_op_O; // @[Map2S.scala 19:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_27(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I1_0_0,
  output [7:0] O_0_0
);
  wire  fst_op_clock; // @[Map2S.scala 9:22]
  wire  fst_op_reset; // @[Map2S.scala 9:22]
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0; // @[Map2S.scala 9:22]
  Map2S_26 fst_op ( // @[Map2S.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I1_0(fst_op_I1_0),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_28(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_1_0_0,
  input  [7:0] I0_2_0_0,
  input  [7:0] I0_3_0_0,
  input  [7:0] I0_4_0_0,
  input  [7:0] I0_5_0_0,
  input  [7:0] I0_6_0_0,
  input  [7:0] I0_7_0_0,
  input  [7:0] I0_8_0_0,
  input  [7:0] I0_9_0_0,
  input  [7:0] I0_10_0_0,
  input  [7:0] I0_11_0_0,
  input  [7:0] I0_12_0_0,
  input  [7:0] I0_13_0_0,
  input  [7:0] I0_14_0_0,
  input  [7:0] I0_15_0_0,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_7_0_0,
  input  [7:0] I1_8_0_0,
  input  [7:0] I1_9_0_0,
  input  [7:0] I1_10_0_0,
  input  [7:0] I1_11_0_0,
  input  [7:0] I1_12_0_0,
  input  [7:0] I1_13_0_0,
  input  [7:0] I1_14_0_0,
  input  [7:0] I1_15_0_0,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0,
  output [7:0] O_8_0_0,
  output [7:0] O_9_0_0,
  output [7:0] O_10_0_0,
  output [7:0] O_11_0_0,
  output [7:0] O_12_0_0,
  output [7:0] O_13_0_0,
  output [7:0] O_14_0_0,
  output [7:0] O_15_0_0
);
  wire  fst_op_clock; // @[Map2S.scala 9:22]
  wire  fst_op_reset; // @[Map2S.scala 9:22]
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire  other_ops_0_clock; // @[Map2S.scala 10:86]
  wire  other_ops_0_reset; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire  other_ops_1_clock; // @[Map2S.scala 10:86]
  wire  other_ops_1_reset; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire  other_ops_2_clock; // @[Map2S.scala 10:86]
  wire  other_ops_2_reset; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire  other_ops_3_clock; // @[Map2S.scala 10:86]
  wire  other_ops_3_reset; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[Map2S.scala 10:86]
  wire  other_ops_4_clock; // @[Map2S.scala 10:86]
  wire  other_ops_4_reset; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[Map2S.scala 10:86]
  wire  other_ops_5_clock; // @[Map2S.scala 10:86]
  wire  other_ops_5_reset; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[Map2S.scala 10:86]
  wire  other_ops_6_clock; // @[Map2S.scala 10:86]
  wire  other_ops_6_reset; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[Map2S.scala 10:86]
  wire  other_ops_7_clock; // @[Map2S.scala 10:86]
  wire  other_ops_7_reset; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0; // @[Map2S.scala 10:86]
  wire  other_ops_8_clock; // @[Map2S.scala 10:86]
  wire  other_ops_8_reset; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0; // @[Map2S.scala 10:86]
  wire  other_ops_9_clock; // @[Map2S.scala 10:86]
  wire  other_ops_9_reset; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0; // @[Map2S.scala 10:86]
  wire  other_ops_10_clock; // @[Map2S.scala 10:86]
  wire  other_ops_10_reset; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0; // @[Map2S.scala 10:86]
  wire  other_ops_11_clock; // @[Map2S.scala 10:86]
  wire  other_ops_11_reset; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0; // @[Map2S.scala 10:86]
  wire  other_ops_12_clock; // @[Map2S.scala 10:86]
  wire  other_ops_12_reset; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0; // @[Map2S.scala 10:86]
  wire  other_ops_13_clock; // @[Map2S.scala 10:86]
  wire  other_ops_13_reset; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0; // @[Map2S.scala 10:86]
  wire  other_ops_14_clock; // @[Map2S.scala 10:86]
  wire  other_ops_14_reset; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  Map2S_27 fst_op ( // @[Map2S.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I1_0_0(fst_op_I1_0_0),
    .O_0_0(fst_op_O_0_0)
  );
  Map2S_27 other_ops_0 ( // @[Map2S.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0(other_ops_0_I0_0_0),
    .I1_0_0(other_ops_0_I1_0_0),
    .O_0_0(other_ops_0_O_0_0)
  );
  Map2S_27 other_ops_1 ( // @[Map2S.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0(other_ops_1_I0_0_0),
    .I1_0_0(other_ops_1_I1_0_0),
    .O_0_0(other_ops_1_O_0_0)
  );
  Map2S_27 other_ops_2 ( // @[Map2S.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0(other_ops_2_I0_0_0),
    .I1_0_0(other_ops_2_I1_0_0),
    .O_0_0(other_ops_2_O_0_0)
  );
  Map2S_27 other_ops_3 ( // @[Map2S.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0(other_ops_3_I0_0_0),
    .I1_0_0(other_ops_3_I1_0_0),
    .O_0_0(other_ops_3_O_0_0)
  );
  Map2S_27 other_ops_4 ( // @[Map2S.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0(other_ops_4_I0_0_0),
    .I1_0_0(other_ops_4_I1_0_0),
    .O_0_0(other_ops_4_O_0_0)
  );
  Map2S_27 other_ops_5 ( // @[Map2S.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0(other_ops_5_I0_0_0),
    .I1_0_0(other_ops_5_I1_0_0),
    .O_0_0(other_ops_5_O_0_0)
  );
  Map2S_27 other_ops_6 ( // @[Map2S.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0(other_ops_6_I0_0_0),
    .I1_0_0(other_ops_6_I1_0_0),
    .O_0_0(other_ops_6_O_0_0)
  );
  Map2S_27 other_ops_7 ( // @[Map2S.scala 10:86]
    .clock(other_ops_7_clock),
    .reset(other_ops_7_reset),
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0_0(other_ops_7_I0_0_0),
    .I1_0_0(other_ops_7_I1_0_0),
    .O_0_0(other_ops_7_O_0_0)
  );
  Map2S_27 other_ops_8 ( // @[Map2S.scala 10:86]
    .clock(other_ops_8_clock),
    .reset(other_ops_8_reset),
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0_0(other_ops_8_I0_0_0),
    .I1_0_0(other_ops_8_I1_0_0),
    .O_0_0(other_ops_8_O_0_0)
  );
  Map2S_27 other_ops_9 ( // @[Map2S.scala 10:86]
    .clock(other_ops_9_clock),
    .reset(other_ops_9_reset),
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0_0(other_ops_9_I0_0_0),
    .I1_0_0(other_ops_9_I1_0_0),
    .O_0_0(other_ops_9_O_0_0)
  );
  Map2S_27 other_ops_10 ( // @[Map2S.scala 10:86]
    .clock(other_ops_10_clock),
    .reset(other_ops_10_reset),
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0_0(other_ops_10_I0_0_0),
    .I1_0_0(other_ops_10_I1_0_0),
    .O_0_0(other_ops_10_O_0_0)
  );
  Map2S_27 other_ops_11 ( // @[Map2S.scala 10:86]
    .clock(other_ops_11_clock),
    .reset(other_ops_11_reset),
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0_0(other_ops_11_I0_0_0),
    .I1_0_0(other_ops_11_I1_0_0),
    .O_0_0(other_ops_11_O_0_0)
  );
  Map2S_27 other_ops_12 ( // @[Map2S.scala 10:86]
    .clock(other_ops_12_clock),
    .reset(other_ops_12_reset),
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0_0(other_ops_12_I0_0_0),
    .I1_0_0(other_ops_12_I1_0_0),
    .O_0_0(other_ops_12_O_0_0)
  );
  Map2S_27 other_ops_13 ( // @[Map2S.scala 10:86]
    .clock(other_ops_13_clock),
    .reset(other_ops_13_reset),
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0_0(other_ops_13_I0_0_0),
    .I1_0_0(other_ops_13_I1_0_0),
    .O_0_0(other_ops_13_O_0_0)
  );
  Map2S_27 other_ops_14 ( // @[Map2S.scala 10:86]
    .clock(other_ops_14_clock),
    .reset(other_ops_14_reset),
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0_0(other_ops_14_I0_0_0),
    .I1_0_0(other_ops_14_I1_0_0),
    .O_0_0(other_ops_14_O_0_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[Map2S.scala 24:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[Map2S.scala 24:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[Map2S.scala 24:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[Map2S.scala 24:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[Map2S.scala 24:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[Map2S.scala 24:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[Map2S.scala 24:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[Map2S.scala 24:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[Map2S.scala 24:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_0 = I1_0_0_0; // @[Map2S.scala 18:13]
  assign other_ops_0_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_0_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0 = I0_1_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0_0 = I1_1_0_0; // @[Map2S.scala 23:43]
  assign other_ops_1_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_1_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0 = I0_2_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0_0 = I1_2_0_0; // @[Map2S.scala 23:43]
  assign other_ops_2_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_2_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0 = I0_3_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0_0 = I1_3_0_0; // @[Map2S.scala 23:43]
  assign other_ops_3_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_3_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0 = I0_4_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0_0 = I1_4_0_0; // @[Map2S.scala 23:43]
  assign other_ops_4_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_4_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0 = I0_5_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0_0 = I1_5_0_0; // @[Map2S.scala 23:43]
  assign other_ops_5_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_5_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0 = I0_6_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0_0 = I1_6_0_0; // @[Map2S.scala 23:43]
  assign other_ops_6_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_6_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0 = I0_7_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0_0 = I1_7_0_0; // @[Map2S.scala 23:43]
  assign other_ops_7_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_7_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0_0 = I0_8_0_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I1_0_0 = I1_8_0_0; // @[Map2S.scala 23:43]
  assign other_ops_8_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_8_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0_0 = I0_9_0_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I1_0_0 = I1_9_0_0; // @[Map2S.scala 23:43]
  assign other_ops_9_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_9_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0_0 = I0_10_0_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I1_0_0 = I1_10_0_0; // @[Map2S.scala 23:43]
  assign other_ops_10_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_10_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0_0 = I0_11_0_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I1_0_0 = I1_11_0_0; // @[Map2S.scala 23:43]
  assign other_ops_11_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_11_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0_0 = I0_12_0_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I1_0_0 = I1_12_0_0; // @[Map2S.scala 23:43]
  assign other_ops_12_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_12_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0_0 = I0_13_0_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I1_0_0 = I1_13_0_0; // @[Map2S.scala 23:43]
  assign other_ops_13_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_13_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0_0 = I0_14_0_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I1_0_0 = I1_14_0_0; // @[Map2S.scala 23:43]
  assign other_ops_14_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_14_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0_0 = I0_15_0_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I1_0_0 = I1_15_0_0; // @[Map2S.scala 23:43]
endmodule
module Map2T_8(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_1_0_0,
  input  [7:0] I0_2_0_0,
  input  [7:0] I0_3_0_0,
  input  [7:0] I0_4_0_0,
  input  [7:0] I0_5_0_0,
  input  [7:0] I0_6_0_0,
  input  [7:0] I0_7_0_0,
  input  [7:0] I0_8_0_0,
  input  [7:0] I0_9_0_0,
  input  [7:0] I0_10_0_0,
  input  [7:0] I0_11_0_0,
  input  [7:0] I0_12_0_0,
  input  [7:0] I0_13_0_0,
  input  [7:0] I0_14_0_0,
  input  [7:0] I0_15_0_0,
  input  [7:0] I1_0_0_0,
  input  [7:0] I1_1_0_0,
  input  [7:0] I1_2_0_0,
  input  [7:0] I1_3_0_0,
  input  [7:0] I1_4_0_0,
  input  [7:0] I1_5_0_0,
  input  [7:0] I1_6_0_0,
  input  [7:0] I1_7_0_0,
  input  [7:0] I1_8_0_0,
  input  [7:0] I1_9_0_0,
  input  [7:0] I1_10_0_0,
  input  [7:0] I1_11_0_0,
  input  [7:0] I1_12_0_0,
  input  [7:0] I1_13_0_0,
  input  [7:0] I1_14_0_0,
  input  [7:0] I1_15_0_0,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0,
  output [7:0] O_8_0_0,
  output [7:0] O_9_0_0,
  output [7:0] O_10_0_0,
  output [7:0] O_11_0_0,
  output [7:0] O_12_0_0,
  output [7:0] O_13_0_0,
  output [7:0] O_14_0_0,
  output [7:0] O_15_0_0
);
  wire  op_clock; // @[Map2T.scala 8:20]
  wire  op_reset; // @[Map2T.scala 8:20]
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_0; // @[Map2T.scala 8:20]
  Map2S_28 op ( // @[Map2T.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0(op_I0_0_0_0),
    .I0_1_0_0(op_I0_1_0_0),
    .I0_2_0_0(op_I0_2_0_0),
    .I0_3_0_0(op_I0_3_0_0),
    .I0_4_0_0(op_I0_4_0_0),
    .I0_5_0_0(op_I0_5_0_0),
    .I0_6_0_0(op_I0_6_0_0),
    .I0_7_0_0(op_I0_7_0_0),
    .I0_8_0_0(op_I0_8_0_0),
    .I0_9_0_0(op_I0_9_0_0),
    .I0_10_0_0(op_I0_10_0_0),
    .I0_11_0_0(op_I0_11_0_0),
    .I0_12_0_0(op_I0_12_0_0),
    .I0_13_0_0(op_I0_13_0_0),
    .I0_14_0_0(op_I0_14_0_0),
    .I0_15_0_0(op_I0_15_0_0),
    .I1_0_0_0(op_I1_0_0_0),
    .I1_1_0_0(op_I1_1_0_0),
    .I1_2_0_0(op_I1_2_0_0),
    .I1_3_0_0(op_I1_3_0_0),
    .I1_4_0_0(op_I1_4_0_0),
    .I1_5_0_0(op_I1_5_0_0),
    .I1_6_0_0(op_I1_6_0_0),
    .I1_7_0_0(op_I1_7_0_0),
    .I1_8_0_0(op_I1_8_0_0),
    .I1_9_0_0(op_I1_9_0_0),
    .I1_10_0_0(op_I1_10_0_0),
    .I1_11_0_0(op_I1_11_0_0),
    .I1_12_0_0(op_I1_12_0_0),
    .I1_13_0_0(op_I1_13_0_0),
    .I1_14_0_0(op_I1_14_0_0),
    .I1_15_0_0(op_I1_15_0_0),
    .O_0_0_0(op_O_0_0_0),
    .O_1_0_0(op_O_1_0_0),
    .O_2_0_0(op_O_2_0_0),
    .O_3_0_0(op_O_3_0_0),
    .O_4_0_0(op_O_4_0_0),
    .O_5_0_0(op_O_5_0_0),
    .O_6_0_0(op_O_6_0_0),
    .O_7_0_0(op_O_7_0_0),
    .O_8_0_0(op_O_8_0_0),
    .O_9_0_0(op_O_9_0_0),
    .O_10_0_0(op_O_10_0_0),
    .O_11_0_0(op_O_11_0_0),
    .O_12_0_0(op_O_12_0_0),
    .O_13_0_0(op_O_13_0_0),
    .O_14_0_0(op_O_14_0_0),
    .O_15_0_0(op_O_15_0_0)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_0 = op_O_2_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_0 = op_O_3_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_0 = op_O_4_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_0 = op_O_5_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_0 = op_O_6_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_0 = op_O_7_0_0; // @[Map2T.scala 17:7]
  assign O_8_0_0 = op_O_8_0_0; // @[Map2T.scala 17:7]
  assign O_9_0_0 = op_O_9_0_0; // @[Map2T.scala 17:7]
  assign O_10_0_0 = op_O_10_0_0; // @[Map2T.scala 17:7]
  assign O_11_0_0 = op_O_11_0_0; // @[Map2T.scala 17:7]
  assign O_12_0_0 = op_O_12_0_0; // @[Map2T.scala 17:7]
  assign O_13_0_0 = op_O_13_0_0; // @[Map2T.scala 17:7]
  assign O_14_0_0 = op_O_14_0_0; // @[Map2T.scala 17:7]
  assign O_15_0_0 = op_O_15_0_0; // @[Map2T.scala 17:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0 = I0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0 = I0_1_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0 = I0_2_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0 = I0_3_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0 = I0_4_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0 = I0_5_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0 = I0_6_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0 = I0_7_0_0; // @[Map2T.scala 15:11]
  assign op_I0_8_0_0 = I0_8_0_0; // @[Map2T.scala 15:11]
  assign op_I0_9_0_0 = I0_9_0_0; // @[Map2T.scala 15:11]
  assign op_I0_10_0_0 = I0_10_0_0; // @[Map2T.scala 15:11]
  assign op_I0_11_0_0 = I0_11_0_0; // @[Map2T.scala 15:11]
  assign op_I0_12_0_0 = I0_12_0_0; // @[Map2T.scala 15:11]
  assign op_I0_13_0_0 = I0_13_0_0; // @[Map2T.scala 15:11]
  assign op_I0_14_0_0 = I0_14_0_0; // @[Map2T.scala 15:11]
  assign op_I0_15_0_0 = I0_15_0_0; // @[Map2T.scala 15:11]
  assign op_I1_0_0_0 = I1_0_0_0; // @[Map2T.scala 16:11]
  assign op_I1_1_0_0 = I1_1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_2_0_0 = I1_2_0_0; // @[Map2T.scala 16:11]
  assign op_I1_3_0_0 = I1_3_0_0; // @[Map2T.scala 16:11]
  assign op_I1_4_0_0 = I1_4_0_0; // @[Map2T.scala 16:11]
  assign op_I1_5_0_0 = I1_5_0_0; // @[Map2T.scala 16:11]
  assign op_I1_6_0_0 = I1_6_0_0; // @[Map2T.scala 16:11]
  assign op_I1_7_0_0 = I1_7_0_0; // @[Map2T.scala 16:11]
  assign op_I1_8_0_0 = I1_8_0_0; // @[Map2T.scala 16:11]
  assign op_I1_9_0_0 = I1_9_0_0; // @[Map2T.scala 16:11]
  assign op_I1_10_0_0 = I1_10_0_0; // @[Map2T.scala 16:11]
  assign op_I1_11_0_0 = I1_11_0_0; // @[Map2T.scala 16:11]
  assign op_I1_12_0_0 = I1_12_0_0; // @[Map2T.scala 16:11]
  assign op_I1_13_0_0 = I1_13_0_0; // @[Map2T.scala 16:11]
  assign op_I1_14_0_0 = I1_14_0_0; // @[Map2T.scala 16:11]
  assign op_I1_15_0_0 = I1_15_0_0; // @[Map2T.scala 16:11]
endmodule
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_1_0_0,
  input  [7:0] I_2_0_0,
  input  [7:0] I_3_0_0,
  input  [7:0] I_4_0_0,
  input  [7:0] I_5_0_0,
  input  [7:0] I_6_0_0,
  input  [7:0] I_7_0_0,
  input  [7:0] I_8_0_0,
  input  [7:0] I_9_0_0,
  input  [7:0] I_10_0_0,
  input  [7:0] I_11_0_0,
  input  [7:0] I_12_0_0,
  input  [7:0] I_13_0_0,
  input  [7:0] I_14_0_0,
  input  [7:0] I_15_0_0,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0,
  output [7:0] O_8_0_0,
  output [7:0] O_9_0_0,
  output [7:0] O_10_0_0,
  output [7:0] O_11_0_0,
  output [7:0] O_12_0_0,
  output [7:0] O_13_0_0,
  output [7:0] O_14_0_0,
  output [7:0] O_15_0_0
);
  wire  n1_clock; // @[Top.scala 103:20]
  wire  n1_valid_up; // @[Top.scala 103:20]
  wire  n1_valid_down; // @[Top.scala 103:20]
  wire [7:0] n1_I_0_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_I_1_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_I_2_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_I_3_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_I_4_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_I_5_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_I_6_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_I_7_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_I_8_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_I_9_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_I_10_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_I_11_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_I_12_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_I_13_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_I_14_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_I_15_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_0_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_1_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_2_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_3_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_4_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_5_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_6_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_7_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_8_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_9_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_10_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_11_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_12_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_13_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_14_0_0; // @[Top.scala 103:20]
  wire [7:0] n1_O_15_0_0; // @[Top.scala 103:20]
  wire  n2_clock; // @[Top.scala 106:20]
  wire  n2_reset; // @[Top.scala 106:20]
  wire  n2_valid_up; // @[Top.scala 106:20]
  wire  n2_valid_down; // @[Top.scala 106:20]
  wire [7:0] n2_I_0_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_I_1_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_I_2_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_I_3_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_I_4_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_I_5_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_I_6_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_I_7_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_I_8_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_I_9_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_I_10_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_I_11_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_I_12_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_I_13_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_I_14_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_I_15_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_0_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_1_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_2_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_3_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_4_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_5_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_6_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_7_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_8_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_9_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_10_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_11_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_12_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_13_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_14_0_0; // @[Top.scala 106:20]
  wire [7:0] n2_O_15_0_0; // @[Top.scala 106:20]
  wire  n3_clock; // @[Top.scala 109:20]
  wire  n3_reset; // @[Top.scala 109:20]
  wire  n3_valid_up; // @[Top.scala 109:20]
  wire  n3_valid_down; // @[Top.scala 109:20]
  wire [7:0] n3_I_0_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_I_1_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_I_2_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_I_3_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_I_4_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_I_5_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_I_6_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_I_7_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_I_8_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_I_9_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_I_10_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_I_11_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_I_12_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_I_13_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_I_14_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_I_15_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_0_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_1_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_2_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_3_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_4_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_5_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_6_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_7_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_8_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_9_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_10_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_11_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_12_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_13_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_14_0_0; // @[Top.scala 109:20]
  wire [7:0] n3_O_15_0_0; // @[Top.scala 109:20]
  wire  n4_clock; // @[Top.scala 112:20]
  wire  n4_valid_up; // @[Top.scala 112:20]
  wire  n4_valid_down; // @[Top.scala 112:20]
  wire [7:0] n4_I_0_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_I_1_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_I_2_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_I_3_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_I_4_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_I_5_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_I_6_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_I_7_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_I_8_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_I_9_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_I_10_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_I_11_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_I_12_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_I_13_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_I_14_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_I_15_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_0_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_1_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_2_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_3_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_4_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_5_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_6_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_7_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_8_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_9_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_10_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_11_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_12_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_13_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_14_0_0; // @[Top.scala 112:20]
  wire [7:0] n4_O_15_0_0; // @[Top.scala 112:20]
  wire  n5_clock; // @[Top.scala 115:20]
  wire  n5_valid_up; // @[Top.scala 115:20]
  wire  n5_valid_down; // @[Top.scala 115:20]
  wire [7:0] n5_I_0_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_I_1_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_I_2_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_I_3_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_I_4_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_I_5_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_I_6_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_I_7_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_I_8_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_I_9_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_I_10_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_I_11_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_I_12_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_I_13_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_I_14_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_I_15_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_0_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_1_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_2_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_3_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_4_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_5_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_6_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_7_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_8_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_9_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_10_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_11_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_12_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_13_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_14_0_0; // @[Top.scala 115:20]
  wire [7:0] n5_O_15_0_0; // @[Top.scala 115:20]
  wire  n6_valid_up; // @[Top.scala 118:20]
  wire  n6_valid_down; // @[Top.scala 118:20]
  wire [7:0] n6_I0_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I0_1_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I0_2_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I0_3_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I0_4_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I0_5_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I0_6_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I0_7_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I0_8_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I0_9_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I0_10_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I0_11_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I0_12_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I0_13_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I0_14_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I0_15_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_1_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_2_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_3_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_4_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_5_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_6_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_7_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_8_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_9_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_10_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_11_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_12_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_13_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_14_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_I1_15_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_0_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_0_0_0_1; // @[Top.scala 118:20]
  wire [7:0] n6_O_1_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_1_0_0_1; // @[Top.scala 118:20]
  wire [7:0] n6_O_2_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_2_0_0_1; // @[Top.scala 118:20]
  wire [7:0] n6_O_3_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_3_0_0_1; // @[Top.scala 118:20]
  wire [7:0] n6_O_4_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_4_0_0_1; // @[Top.scala 118:20]
  wire [7:0] n6_O_5_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_5_0_0_1; // @[Top.scala 118:20]
  wire [7:0] n6_O_6_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_6_0_0_1; // @[Top.scala 118:20]
  wire [7:0] n6_O_7_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_7_0_0_1; // @[Top.scala 118:20]
  wire [7:0] n6_O_8_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_8_0_0_1; // @[Top.scala 118:20]
  wire [7:0] n6_O_9_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_9_0_0_1; // @[Top.scala 118:20]
  wire [7:0] n6_O_10_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_10_0_0_1; // @[Top.scala 118:20]
  wire [7:0] n6_O_11_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_11_0_0_1; // @[Top.scala 118:20]
  wire [7:0] n6_O_12_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_12_0_0_1; // @[Top.scala 118:20]
  wire [7:0] n6_O_13_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_13_0_0_1; // @[Top.scala 118:20]
  wire [7:0] n6_O_14_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_14_0_0_1; // @[Top.scala 118:20]
  wire [7:0] n6_O_15_0_0_0; // @[Top.scala 118:20]
  wire [7:0] n6_O_15_0_0_1; // @[Top.scala 118:20]
  wire  n19_valid_up; // @[Top.scala 122:21]
  wire  n19_valid_down; // @[Top.scala 122:21]
  wire [7:0] n19_I0_0_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_0_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I0_1_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_1_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I0_2_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_2_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I0_3_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_3_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I0_4_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_4_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I0_5_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_5_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I0_6_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_6_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I0_7_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_7_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I0_8_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_8_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I0_9_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_9_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I0_10_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_10_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I0_11_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_11_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I0_12_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_12_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I0_13_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_13_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I0_14_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_14_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I0_15_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I0_15_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_I1_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I1_1_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I1_2_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I1_3_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I1_4_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I1_5_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I1_6_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I1_7_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I1_8_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I1_9_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I1_10_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I1_11_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I1_12_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I1_13_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I1_14_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_I1_15_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_0_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_0_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_0_0_0_2; // @[Top.scala 122:21]
  wire [7:0] n19_O_1_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_1_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_1_0_0_2; // @[Top.scala 122:21]
  wire [7:0] n19_O_2_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_2_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_2_0_0_2; // @[Top.scala 122:21]
  wire [7:0] n19_O_3_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_3_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_3_0_0_2; // @[Top.scala 122:21]
  wire [7:0] n19_O_4_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_4_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_4_0_0_2; // @[Top.scala 122:21]
  wire [7:0] n19_O_5_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_5_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_5_0_0_2; // @[Top.scala 122:21]
  wire [7:0] n19_O_6_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_6_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_6_0_0_2; // @[Top.scala 122:21]
  wire [7:0] n19_O_7_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_7_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_7_0_0_2; // @[Top.scala 122:21]
  wire [7:0] n19_O_8_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_8_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_8_0_0_2; // @[Top.scala 122:21]
  wire [7:0] n19_O_9_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_9_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_9_0_0_2; // @[Top.scala 122:21]
  wire [7:0] n19_O_10_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_10_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_10_0_0_2; // @[Top.scala 122:21]
  wire [7:0] n19_O_11_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_11_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_11_0_0_2; // @[Top.scala 122:21]
  wire [7:0] n19_O_12_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_12_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_12_0_0_2; // @[Top.scala 122:21]
  wire [7:0] n19_O_13_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_13_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_13_0_0_2; // @[Top.scala 122:21]
  wire [7:0] n19_O_14_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_14_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_14_0_0_2; // @[Top.scala 122:21]
  wire [7:0] n19_O_15_0_0_0; // @[Top.scala 122:21]
  wire [7:0] n19_O_15_0_0_1; // @[Top.scala 122:21]
  wire [7:0] n19_O_15_0_0_2; // @[Top.scala 122:21]
  wire  n40_valid_up; // @[Top.scala 126:21]
  wire  n40_valid_down; // @[Top.scala 126:21]
  wire [7:0] n40_I_0_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_0_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_0_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_I_1_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_1_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_1_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_I_2_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_2_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_2_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_I_3_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_3_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_3_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_I_4_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_4_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_4_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_I_5_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_5_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_5_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_I_6_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_6_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_6_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_I_7_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_7_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_7_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_I_8_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_8_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_8_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_I_9_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_9_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_9_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_I_10_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_10_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_10_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_I_11_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_11_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_11_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_I_12_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_12_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_12_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_I_13_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_13_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_13_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_I_14_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_14_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_14_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_I_15_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_I_15_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_I_15_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_0_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_0_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_0_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_1_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_1_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_1_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_2_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_2_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_2_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_3_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_3_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_3_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_4_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_4_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_4_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_5_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_5_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_5_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_6_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_6_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_6_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_7_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_7_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_7_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_8_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_8_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_8_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_9_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_9_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_9_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_10_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_10_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_10_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_11_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_11_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_11_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_12_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_12_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_12_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_13_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_13_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_13_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_14_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_14_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_14_0_2; // @[Top.scala 126:21]
  wire [7:0] n40_O_15_0_0; // @[Top.scala 126:21]
  wire [7:0] n40_O_15_0_1; // @[Top.scala 126:21]
  wire [7:0] n40_O_15_0_2; // @[Top.scala 126:21]
  wire  n41_clock; // @[Top.scala 129:21]
  wire  n41_valid_up; // @[Top.scala 129:21]
  wire  n41_valid_down; // @[Top.scala 129:21]
  wire [7:0] n41_I_0_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_I_1_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_I_2_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_I_3_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_I_4_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_I_5_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_I_6_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_I_7_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_I_8_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_I_9_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_I_10_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_I_11_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_I_12_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_I_13_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_I_14_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_I_15_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_0_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_1_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_2_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_3_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_4_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_5_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_6_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_7_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_8_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_9_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_10_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_11_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_12_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_13_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_14_0_0; // @[Top.scala 129:21]
  wire [7:0] n41_O_15_0_0; // @[Top.scala 129:21]
  wire  n42_clock; // @[Top.scala 132:21]
  wire  n42_valid_up; // @[Top.scala 132:21]
  wire  n42_valid_down; // @[Top.scala 132:21]
  wire [7:0] n42_I_0_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_I_1_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_I_2_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_I_3_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_I_4_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_I_5_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_I_6_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_I_7_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_I_8_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_I_9_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_I_10_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_I_11_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_I_12_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_I_13_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_I_14_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_I_15_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_0_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_1_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_2_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_3_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_4_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_5_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_6_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_7_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_8_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_9_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_10_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_11_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_12_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_13_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_14_0_0; // @[Top.scala 132:21]
  wire [7:0] n42_O_15_0_0; // @[Top.scala 132:21]
  wire  n43_valid_up; // @[Top.scala 135:21]
  wire  n43_valid_down; // @[Top.scala 135:21]
  wire [7:0] n43_I0_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I0_1_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I0_2_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I0_3_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I0_4_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I0_5_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I0_6_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I0_7_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I0_8_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I0_9_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I0_10_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I0_11_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I0_12_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I0_13_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I0_14_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I0_15_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_1_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_2_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_3_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_4_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_5_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_6_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_7_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_8_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_9_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_10_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_11_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_12_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_13_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_14_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_I1_15_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_0_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_0_0_0_1; // @[Top.scala 135:21]
  wire [7:0] n43_O_1_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_1_0_0_1; // @[Top.scala 135:21]
  wire [7:0] n43_O_2_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_2_0_0_1; // @[Top.scala 135:21]
  wire [7:0] n43_O_3_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_3_0_0_1; // @[Top.scala 135:21]
  wire [7:0] n43_O_4_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_4_0_0_1; // @[Top.scala 135:21]
  wire [7:0] n43_O_5_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_5_0_0_1; // @[Top.scala 135:21]
  wire [7:0] n43_O_6_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_6_0_0_1; // @[Top.scala 135:21]
  wire [7:0] n43_O_7_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_7_0_0_1; // @[Top.scala 135:21]
  wire [7:0] n43_O_8_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_8_0_0_1; // @[Top.scala 135:21]
  wire [7:0] n43_O_9_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_9_0_0_1; // @[Top.scala 135:21]
  wire [7:0] n43_O_10_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_10_0_0_1; // @[Top.scala 135:21]
  wire [7:0] n43_O_11_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_11_0_0_1; // @[Top.scala 135:21]
  wire [7:0] n43_O_12_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_12_0_0_1; // @[Top.scala 135:21]
  wire [7:0] n43_O_13_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_13_0_0_1; // @[Top.scala 135:21]
  wire [7:0] n43_O_14_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_14_0_0_1; // @[Top.scala 135:21]
  wire [7:0] n43_O_15_0_0_0; // @[Top.scala 135:21]
  wire [7:0] n43_O_15_0_0_1; // @[Top.scala 135:21]
  wire  n56_valid_up; // @[Top.scala 139:21]
  wire  n56_valid_down; // @[Top.scala 139:21]
  wire [7:0] n56_I0_0_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_0_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I0_1_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_1_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I0_2_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_2_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I0_3_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_3_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I0_4_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_4_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I0_5_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_5_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I0_6_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_6_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I0_7_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_7_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I0_8_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_8_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I0_9_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_9_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I0_10_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_10_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I0_11_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_11_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I0_12_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_12_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I0_13_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_13_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I0_14_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_14_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I0_15_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I0_15_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_I1_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I1_1_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I1_2_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I1_3_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I1_4_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I1_5_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I1_6_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I1_7_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I1_8_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I1_9_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I1_10_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I1_11_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I1_12_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I1_13_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I1_14_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_I1_15_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_0_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_0_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_0_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n56_O_1_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_1_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_1_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n56_O_2_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_2_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_2_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n56_O_3_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_3_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_3_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n56_O_4_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_4_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_4_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n56_O_5_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_5_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_5_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n56_O_6_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_6_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_6_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n56_O_7_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_7_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_7_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n56_O_8_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_8_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_8_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n56_O_9_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_9_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_9_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n56_O_10_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_10_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_10_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n56_O_11_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_11_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_11_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n56_O_12_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_12_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_12_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n56_O_13_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_13_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_13_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n56_O_14_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_14_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_14_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n56_O_15_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n56_O_15_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n56_O_15_0_0_2; // @[Top.scala 139:21]
  wire  n77_valid_up; // @[Top.scala 143:21]
  wire  n77_valid_down; // @[Top.scala 143:21]
  wire [7:0] n77_I_0_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_0_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_0_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_I_1_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_1_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_1_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_I_2_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_2_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_2_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_I_3_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_3_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_3_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_I_4_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_4_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_4_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_I_5_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_5_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_5_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_I_6_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_6_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_6_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_I_7_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_7_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_7_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_I_8_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_8_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_8_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_I_9_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_9_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_9_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_I_10_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_10_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_10_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_I_11_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_11_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_11_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_I_12_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_12_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_12_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_I_13_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_13_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_13_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_I_14_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_14_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_14_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_I_15_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_I_15_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_I_15_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_0_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_0_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_0_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_1_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_1_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_1_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_2_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_2_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_2_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_3_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_3_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_3_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_4_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_4_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_4_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_5_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_5_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_5_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_6_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_6_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_6_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_7_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_7_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_7_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_8_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_8_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_8_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_9_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_9_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_9_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_10_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_10_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_10_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_11_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_11_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_11_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_12_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_12_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_12_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_13_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_13_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_13_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_14_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_14_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_14_0_2; // @[Top.scala 143:21]
  wire [7:0] n77_O_15_0_0; // @[Top.scala 143:21]
  wire [7:0] n77_O_15_0_1; // @[Top.scala 143:21]
  wire [7:0] n77_O_15_0_2; // @[Top.scala 143:21]
  wire  n78_valid_up; // @[Top.scala 146:21]
  wire  n78_valid_down; // @[Top.scala 146:21]
  wire [7:0] n78_I0_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I0_1_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_1_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_1_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I0_2_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_2_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_2_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I0_3_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_3_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_3_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I0_4_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_4_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_4_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I0_5_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_5_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_5_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I0_6_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_6_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_6_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I0_7_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_7_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_7_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I0_8_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_8_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_8_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I0_9_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_9_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_9_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I0_10_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_10_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_10_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I0_11_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_11_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_11_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I0_12_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_12_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_12_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I0_13_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_13_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_13_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I0_14_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_14_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_14_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I0_15_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I0_15_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I0_15_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_1_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_1_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_1_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_2_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_2_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_2_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_3_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_3_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_3_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_4_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_4_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_4_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_5_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_5_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_5_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_6_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_6_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_6_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_7_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_7_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_7_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_8_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_8_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_8_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_9_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_9_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_9_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_10_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_10_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_10_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_11_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_11_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_11_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_12_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_12_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_12_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_13_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_13_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_13_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_14_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_14_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_14_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_I1_15_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_I1_15_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_I1_15_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_0_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_0_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_0_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_0_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_0_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_0_0_1_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_1_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_1_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_1_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_1_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_1_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_1_0_1_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_2_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_2_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_2_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_2_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_2_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_2_0_1_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_3_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_3_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_3_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_3_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_3_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_3_0_1_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_4_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_4_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_4_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_4_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_4_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_4_0_1_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_5_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_5_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_5_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_5_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_5_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_5_0_1_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_6_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_6_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_6_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_6_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_6_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_6_0_1_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_7_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_7_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_7_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_7_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_7_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_7_0_1_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_8_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_8_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_8_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_8_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_8_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_8_0_1_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_9_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_9_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_9_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_9_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_9_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_9_0_1_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_10_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_10_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_10_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_10_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_10_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_10_0_1_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_11_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_11_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_11_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_11_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_11_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_11_0_1_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_12_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_12_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_12_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_12_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_12_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_12_0_1_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_13_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_13_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_13_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_13_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_13_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_13_0_1_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_14_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_14_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_14_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_14_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_14_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_14_0_1_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_15_0_0_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_15_0_0_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_15_0_0_2; // @[Top.scala 146:21]
  wire [7:0] n78_O_15_0_1_0; // @[Top.scala 146:21]
  wire [7:0] n78_O_15_0_1_1; // @[Top.scala 146:21]
  wire [7:0] n78_O_15_0_1_2; // @[Top.scala 146:21]
  wire  n88_clock; // @[Top.scala 150:21]
  wire  n88_valid_up; // @[Top.scala 150:21]
  wire  n88_valid_down; // @[Top.scala 150:21]
  wire [7:0] n88_I_0_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_I_1_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_I_2_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_I_3_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_I_4_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_I_5_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_I_6_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_I_7_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_I_8_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_I_9_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_I_10_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_I_11_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_I_12_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_I_13_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_I_14_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_I_15_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_0_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_1_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_2_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_3_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_4_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_5_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_6_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_7_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_8_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_9_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_10_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_11_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_12_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_13_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_14_0_0; // @[Top.scala 150:21]
  wire [7:0] n88_O_15_0_0; // @[Top.scala 150:21]
  wire  n89_clock; // @[Top.scala 153:21]
  wire  n89_valid_up; // @[Top.scala 153:21]
  wire  n89_valid_down; // @[Top.scala 153:21]
  wire [7:0] n89_I_0_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_I_1_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_I_2_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_I_3_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_I_4_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_I_5_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_I_6_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_I_7_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_I_8_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_I_9_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_I_10_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_I_11_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_I_12_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_I_13_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_I_14_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_I_15_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_0_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_1_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_2_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_3_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_4_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_5_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_6_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_7_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_8_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_9_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_10_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_11_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_12_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_13_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_14_0_0; // @[Top.scala 153:21]
  wire [7:0] n89_O_15_0_0; // @[Top.scala 153:21]
  wire  n90_valid_up; // @[Top.scala 156:21]
  wire  n90_valid_down; // @[Top.scala 156:21]
  wire [7:0] n90_I0_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I0_1_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I0_2_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I0_3_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I0_4_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I0_5_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I0_6_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I0_7_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I0_8_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I0_9_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I0_10_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I0_11_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I0_12_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I0_13_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I0_14_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I0_15_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_1_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_2_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_3_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_4_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_5_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_6_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_7_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_8_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_9_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_10_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_11_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_12_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_13_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_14_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_I1_15_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_0_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_0_0_0_1; // @[Top.scala 156:21]
  wire [7:0] n90_O_1_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_1_0_0_1; // @[Top.scala 156:21]
  wire [7:0] n90_O_2_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_2_0_0_1; // @[Top.scala 156:21]
  wire [7:0] n90_O_3_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_3_0_0_1; // @[Top.scala 156:21]
  wire [7:0] n90_O_4_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_4_0_0_1; // @[Top.scala 156:21]
  wire [7:0] n90_O_5_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_5_0_0_1; // @[Top.scala 156:21]
  wire [7:0] n90_O_6_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_6_0_0_1; // @[Top.scala 156:21]
  wire [7:0] n90_O_7_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_7_0_0_1; // @[Top.scala 156:21]
  wire [7:0] n90_O_8_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_8_0_0_1; // @[Top.scala 156:21]
  wire [7:0] n90_O_9_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_9_0_0_1; // @[Top.scala 156:21]
  wire [7:0] n90_O_10_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_10_0_0_1; // @[Top.scala 156:21]
  wire [7:0] n90_O_11_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_11_0_0_1; // @[Top.scala 156:21]
  wire [7:0] n90_O_12_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_12_0_0_1; // @[Top.scala 156:21]
  wire [7:0] n90_O_13_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_13_0_0_1; // @[Top.scala 156:21]
  wire [7:0] n90_O_14_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_14_0_0_1; // @[Top.scala 156:21]
  wire [7:0] n90_O_15_0_0_0; // @[Top.scala 156:21]
  wire [7:0] n90_O_15_0_0_1; // @[Top.scala 156:21]
  wire  n103_valid_up; // @[Top.scala 160:22]
  wire  n103_valid_down; // @[Top.scala 160:22]
  wire [7:0] n103_I0_0_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_0_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I0_1_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_1_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I0_2_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_2_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I0_3_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_3_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I0_4_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_4_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I0_5_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_5_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I0_6_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_6_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I0_7_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_7_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I0_8_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_8_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I0_9_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_9_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I0_10_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_10_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I0_11_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_11_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I0_12_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_12_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I0_13_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_13_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I0_14_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_14_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I0_15_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I0_15_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_I1_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I1_1_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I1_2_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I1_3_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I1_4_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I1_5_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I1_6_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I1_7_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I1_8_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I1_9_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I1_10_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I1_11_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I1_12_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I1_13_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I1_14_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_I1_15_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_0_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_0_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_0_0_0_2; // @[Top.scala 160:22]
  wire [7:0] n103_O_1_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_1_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_1_0_0_2; // @[Top.scala 160:22]
  wire [7:0] n103_O_2_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_2_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_2_0_0_2; // @[Top.scala 160:22]
  wire [7:0] n103_O_3_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_3_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_3_0_0_2; // @[Top.scala 160:22]
  wire [7:0] n103_O_4_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_4_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_4_0_0_2; // @[Top.scala 160:22]
  wire [7:0] n103_O_5_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_5_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_5_0_0_2; // @[Top.scala 160:22]
  wire [7:0] n103_O_6_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_6_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_6_0_0_2; // @[Top.scala 160:22]
  wire [7:0] n103_O_7_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_7_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_7_0_0_2; // @[Top.scala 160:22]
  wire [7:0] n103_O_8_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_8_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_8_0_0_2; // @[Top.scala 160:22]
  wire [7:0] n103_O_9_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_9_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_9_0_0_2; // @[Top.scala 160:22]
  wire [7:0] n103_O_10_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_10_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_10_0_0_2; // @[Top.scala 160:22]
  wire [7:0] n103_O_11_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_11_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_11_0_0_2; // @[Top.scala 160:22]
  wire [7:0] n103_O_12_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_12_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_12_0_0_2; // @[Top.scala 160:22]
  wire [7:0] n103_O_13_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_13_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_13_0_0_2; // @[Top.scala 160:22]
  wire [7:0] n103_O_14_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_14_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_14_0_0_2; // @[Top.scala 160:22]
  wire [7:0] n103_O_15_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n103_O_15_0_0_1; // @[Top.scala 160:22]
  wire [7:0] n103_O_15_0_0_2; // @[Top.scala 160:22]
  wire  n124_valid_up; // @[Top.scala 164:22]
  wire  n124_valid_down; // @[Top.scala 164:22]
  wire [7:0] n124_I_0_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_0_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_0_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_I_1_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_1_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_1_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_I_2_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_2_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_2_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_I_3_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_3_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_3_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_I_4_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_4_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_4_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_I_5_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_5_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_5_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_I_6_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_6_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_6_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_I_7_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_7_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_7_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_I_8_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_8_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_8_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_I_9_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_9_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_9_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_I_10_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_10_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_10_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_I_11_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_11_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_11_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_I_12_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_12_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_12_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_I_13_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_13_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_13_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_I_14_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_14_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_14_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_I_15_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_I_15_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_I_15_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_0_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_0_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_0_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_1_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_1_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_1_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_2_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_2_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_2_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_3_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_3_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_3_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_4_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_4_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_4_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_5_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_5_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_5_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_6_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_6_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_6_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_7_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_7_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_7_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_8_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_8_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_8_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_9_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_9_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_9_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_10_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_10_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_10_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_11_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_11_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_11_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_12_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_12_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_12_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_13_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_13_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_13_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_14_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_14_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_14_0_2; // @[Top.scala 164:22]
  wire [7:0] n124_O_15_0_0; // @[Top.scala 164:22]
  wire [7:0] n124_O_15_0_1; // @[Top.scala 164:22]
  wire [7:0] n124_O_15_0_2; // @[Top.scala 164:22]
  wire  n125_valid_up; // @[Top.scala 167:22]
  wire  n125_valid_down; // @[Top.scala 167:22]
  wire [7:0] n125_I0_0_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_0_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_0_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_0_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_0_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_0_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_1_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_1_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_1_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_1_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_1_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_1_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_2_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_2_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_2_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_2_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_2_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_2_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_3_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_3_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_3_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_3_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_3_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_3_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_4_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_4_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_4_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_4_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_4_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_4_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_5_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_5_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_5_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_5_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_5_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_5_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_6_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_6_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_6_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_6_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_6_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_6_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_7_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_7_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_7_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_7_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_7_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_7_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_8_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_8_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_8_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_8_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_8_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_8_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_9_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_9_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_9_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_9_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_9_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_9_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_10_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_10_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_10_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_10_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_10_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_10_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_11_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_11_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_11_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_11_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_11_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_11_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_12_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_12_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_12_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_12_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_12_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_12_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_13_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_13_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_13_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_13_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_13_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_13_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_14_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_14_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_14_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_14_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_14_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_14_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_15_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_15_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_15_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I0_15_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_I0_15_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_I0_15_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_1_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_1_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_1_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_2_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_2_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_2_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_3_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_3_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_3_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_4_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_4_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_4_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_5_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_5_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_5_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_6_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_6_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_6_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_7_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_7_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_7_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_8_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_8_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_8_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_9_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_9_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_9_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_10_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_10_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_10_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_11_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_11_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_11_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_12_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_12_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_12_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_13_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_13_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_13_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_14_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_14_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_14_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_I1_15_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_I1_15_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_I1_15_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_0_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_0_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_0_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_0_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_0_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_0_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_0_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_0_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_0_0_2_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_1_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_1_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_1_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_1_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_1_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_1_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_1_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_1_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_1_0_2_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_2_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_2_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_2_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_2_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_2_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_2_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_2_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_2_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_2_0_2_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_3_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_3_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_3_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_3_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_3_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_3_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_3_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_3_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_3_0_2_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_4_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_4_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_4_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_4_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_4_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_4_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_4_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_4_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_4_0_2_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_5_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_5_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_5_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_5_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_5_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_5_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_5_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_5_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_5_0_2_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_6_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_6_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_6_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_6_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_6_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_6_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_6_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_6_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_6_0_2_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_7_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_7_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_7_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_7_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_7_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_7_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_7_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_7_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_7_0_2_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_8_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_8_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_8_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_8_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_8_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_8_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_8_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_8_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_8_0_2_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_9_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_9_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_9_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_9_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_9_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_9_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_9_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_9_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_9_0_2_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_10_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_10_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_10_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_10_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_10_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_10_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_10_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_10_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_10_0_2_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_11_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_11_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_11_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_11_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_11_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_11_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_11_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_11_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_11_0_2_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_12_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_12_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_12_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_12_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_12_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_12_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_12_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_12_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_12_0_2_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_13_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_13_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_13_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_13_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_13_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_13_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_13_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_13_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_13_0_2_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_14_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_14_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_14_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_14_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_14_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_14_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_14_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_14_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_14_0_2_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_15_0_0_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_15_0_0_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_15_0_0_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_15_0_1_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_15_0_1_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_15_0_1_2; // @[Top.scala 167:22]
  wire [7:0] n125_O_15_0_2_0; // @[Top.scala 167:22]
  wire [7:0] n125_O_15_0_2_1; // @[Top.scala 167:22]
  wire [7:0] n125_O_15_0_2_2; // @[Top.scala 167:22]
  wire  n141_valid_up; // @[Top.scala 171:22]
  wire  n141_valid_down; // @[Top.scala 171:22]
  wire [7:0] n141_I_0_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_0_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_0_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_0_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_0_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_0_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_0_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_0_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_0_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_1_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_1_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_1_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_1_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_1_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_1_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_1_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_1_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_1_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_2_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_2_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_2_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_2_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_2_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_2_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_2_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_2_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_2_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_3_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_3_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_3_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_3_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_3_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_3_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_3_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_3_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_3_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_4_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_4_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_4_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_4_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_4_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_4_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_4_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_4_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_4_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_5_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_5_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_5_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_5_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_5_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_5_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_5_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_5_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_5_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_6_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_6_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_6_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_6_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_6_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_6_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_6_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_6_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_6_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_7_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_7_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_7_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_7_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_7_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_7_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_7_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_7_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_7_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_8_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_8_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_8_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_8_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_8_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_8_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_8_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_8_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_8_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_9_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_9_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_9_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_9_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_9_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_9_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_9_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_9_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_9_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_10_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_10_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_10_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_10_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_10_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_10_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_10_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_10_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_10_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_11_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_11_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_11_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_11_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_11_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_11_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_11_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_11_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_11_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_12_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_12_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_12_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_12_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_12_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_12_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_12_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_12_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_12_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_13_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_13_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_13_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_13_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_13_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_13_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_13_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_13_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_13_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_14_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_14_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_14_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_14_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_14_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_14_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_14_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_14_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_14_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_15_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_15_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_15_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_15_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_15_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_15_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_I_15_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_I_15_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_I_15_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_0_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_0_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_0_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_0_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_0_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_0_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_0_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_0_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_0_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_1_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_1_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_1_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_1_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_1_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_1_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_1_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_1_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_1_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_2_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_2_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_2_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_2_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_2_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_2_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_2_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_2_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_2_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_3_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_3_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_3_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_3_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_3_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_3_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_3_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_3_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_3_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_4_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_4_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_4_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_4_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_4_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_4_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_4_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_4_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_4_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_5_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_5_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_5_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_5_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_5_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_5_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_5_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_5_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_5_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_6_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_6_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_6_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_6_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_6_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_6_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_6_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_6_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_6_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_7_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_7_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_7_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_7_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_7_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_7_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_7_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_7_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_7_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_8_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_8_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_8_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_8_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_8_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_8_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_8_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_8_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_8_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_9_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_9_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_9_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_9_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_9_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_9_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_9_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_9_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_9_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_10_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_10_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_10_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_10_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_10_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_10_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_10_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_10_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_10_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_11_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_11_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_11_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_11_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_11_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_11_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_11_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_11_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_11_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_12_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_12_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_12_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_12_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_12_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_12_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_12_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_12_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_12_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_13_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_13_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_13_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_13_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_13_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_13_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_13_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_13_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_13_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_14_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_14_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_14_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_14_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_14_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_14_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_14_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_14_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_14_2_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_15_0_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_15_0_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_15_0_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_15_1_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_15_1_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_15_1_2; // @[Top.scala 171:22]
  wire [7:0] n141_O_15_2_0; // @[Top.scala 171:22]
  wire [7:0] n141_O_15_2_1; // @[Top.scala 171:22]
  wire [7:0] n141_O_15_2_2; // @[Top.scala 171:22]
  wire  n183_clock; // @[Top.scala 174:22]
  wire  n183_reset; // @[Top.scala 174:22]
  wire  n183_valid_up; // @[Top.scala 174:22]
  wire  n183_valid_down; // @[Top.scala 174:22]
  wire [7:0] n183_I_0_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_0_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_0_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_0_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_0_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_0_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_0_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_0_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_0_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_1_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_1_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_1_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_1_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_1_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_1_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_1_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_1_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_1_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_2_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_2_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_2_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_2_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_2_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_2_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_2_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_2_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_2_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_3_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_3_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_3_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_3_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_3_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_3_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_3_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_3_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_3_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_4_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_4_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_4_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_4_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_4_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_4_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_4_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_4_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_4_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_5_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_5_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_5_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_5_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_5_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_5_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_5_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_5_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_5_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_6_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_6_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_6_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_6_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_6_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_6_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_6_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_6_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_6_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_7_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_7_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_7_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_7_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_7_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_7_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_7_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_7_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_7_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_8_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_8_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_8_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_8_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_8_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_8_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_8_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_8_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_8_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_9_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_9_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_9_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_9_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_9_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_9_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_9_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_9_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_9_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_10_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_10_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_10_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_10_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_10_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_10_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_10_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_10_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_10_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_11_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_11_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_11_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_11_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_11_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_11_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_11_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_11_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_11_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_12_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_12_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_12_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_12_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_12_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_12_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_12_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_12_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_12_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_13_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_13_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_13_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_13_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_13_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_13_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_13_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_13_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_13_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_14_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_14_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_14_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_14_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_14_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_14_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_14_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_14_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_14_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_15_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_15_0_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_15_0_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_15_1_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_15_1_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_15_1_2; // @[Top.scala 174:22]
  wire [7:0] n183_I_15_2_0; // @[Top.scala 174:22]
  wire [7:0] n183_I_15_2_1; // @[Top.scala 174:22]
  wire [7:0] n183_I_15_2_2; // @[Top.scala 174:22]
  wire [7:0] n183_O_0_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_O_1_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_O_2_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_O_3_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_O_4_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_O_5_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_O_6_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_O_7_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_O_8_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_O_9_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_O_10_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_O_11_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_O_12_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_O_13_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_O_14_0_0; // @[Top.scala 174:22]
  wire [7:0] n183_O_15_0_0; // @[Top.scala 174:22]
  wire  n184_clock; // @[Top.scala 177:22]
  wire  n184_reset; // @[Top.scala 177:22]
  wire  n184_valid_up; // @[Top.scala 177:22]
  wire  n184_valid_down; // @[Top.scala 177:22]
  wire [7:0] n184_I_0_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_I_1_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_I_2_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_I_3_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_I_4_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_I_5_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_I_6_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_I_7_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_I_8_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_I_9_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_I_10_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_I_11_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_I_12_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_I_13_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_I_14_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_I_15_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_0_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_1_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_2_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_3_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_4_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_5_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_6_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_7_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_8_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_9_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_10_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_11_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_12_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_13_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_14_0_0; // @[Top.scala 177:22]
  wire [7:0] n184_O_15_0_0; // @[Top.scala 177:22]
  wire  n185_clock; // @[Top.scala 180:22]
  wire  n185_reset; // @[Top.scala 180:22]
  wire  n185_valid_up; // @[Top.scala 180:22]
  wire  n185_valid_down; // @[Top.scala 180:22]
  wire [7:0] n185_I0_0_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I0_1_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I0_2_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I0_3_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I0_4_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I0_5_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I0_6_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I0_7_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I0_8_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I0_9_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I0_10_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I0_11_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I0_12_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I0_13_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I0_14_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I0_15_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_0_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_1_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_2_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_3_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_4_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_5_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_6_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_7_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_8_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_9_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_10_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_11_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_12_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_13_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_14_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_I1_15_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_0_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_1_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_2_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_3_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_4_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_5_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_6_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_7_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_8_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_9_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_10_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_11_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_12_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_13_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_14_0_0; // @[Top.scala 180:22]
  wire [7:0] n185_O_15_0_0; // @[Top.scala 180:22]
  wire  n217_clock; // @[Top.scala 184:22]
  wire  n217_valid_up; // @[Top.scala 184:22]
  wire  n217_valid_down; // @[Top.scala 184:22]
  wire [7:0] n217_I_0_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_I_1_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_I_2_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_I_3_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_I_4_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_I_5_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_I_6_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_I_7_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_I_8_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_I_9_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_I_10_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_I_11_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_I_12_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_I_13_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_I_14_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_I_15_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_0_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_1_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_2_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_3_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_4_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_5_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_6_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_7_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_8_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_9_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_10_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_11_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_12_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_13_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_14_0_0; // @[Top.scala 184:22]
  wire [7:0] n217_O_15_0_0; // @[Top.scala 184:22]
  wire  n218_clock; // @[Top.scala 187:22]
  wire  n218_valid_up; // @[Top.scala 187:22]
  wire  n218_valid_down; // @[Top.scala 187:22]
  wire [7:0] n218_I_0_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_I_1_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_I_2_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_I_3_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_I_4_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_I_5_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_I_6_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_I_7_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_I_8_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_I_9_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_I_10_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_I_11_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_I_12_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_I_13_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_I_14_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_I_15_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_0_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_1_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_2_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_3_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_4_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_5_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_6_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_7_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_8_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_9_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_10_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_11_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_12_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_13_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_14_0_0; // @[Top.scala 187:22]
  wire [7:0] n218_O_15_0_0; // @[Top.scala 187:22]
  wire  n219_clock; // @[Top.scala 190:22]
  wire  n219_valid_up; // @[Top.scala 190:22]
  wire  n219_valid_down; // @[Top.scala 190:22]
  wire [7:0] n219_I_0_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_I_1_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_I_2_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_I_3_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_I_4_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_I_5_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_I_6_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_I_7_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_I_8_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_I_9_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_I_10_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_I_11_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_I_12_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_I_13_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_I_14_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_I_15_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_0_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_1_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_2_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_3_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_4_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_5_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_6_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_7_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_8_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_9_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_10_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_11_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_12_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_13_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_14_0_0; // @[Top.scala 190:22]
  wire [7:0] n219_O_15_0_0; // @[Top.scala 190:22]
  FIFO n1 ( // @[Top.scala 103:20]
    .clock(n1_clock),
    .valid_up(n1_valid_up),
    .valid_down(n1_valid_down),
    .I_0_0_0(n1_I_0_0_0),
    .I_1_0_0(n1_I_1_0_0),
    .I_2_0_0(n1_I_2_0_0),
    .I_3_0_0(n1_I_3_0_0),
    .I_4_0_0(n1_I_4_0_0),
    .I_5_0_0(n1_I_5_0_0),
    .I_6_0_0(n1_I_6_0_0),
    .I_7_0_0(n1_I_7_0_0),
    .I_8_0_0(n1_I_8_0_0),
    .I_9_0_0(n1_I_9_0_0),
    .I_10_0_0(n1_I_10_0_0),
    .I_11_0_0(n1_I_11_0_0),
    .I_12_0_0(n1_I_12_0_0),
    .I_13_0_0(n1_I_13_0_0),
    .I_14_0_0(n1_I_14_0_0),
    .I_15_0_0(n1_I_15_0_0),
    .O_0_0_0(n1_O_0_0_0),
    .O_1_0_0(n1_O_1_0_0),
    .O_2_0_0(n1_O_2_0_0),
    .O_3_0_0(n1_O_3_0_0),
    .O_4_0_0(n1_O_4_0_0),
    .O_5_0_0(n1_O_5_0_0),
    .O_6_0_0(n1_O_6_0_0),
    .O_7_0_0(n1_O_7_0_0),
    .O_8_0_0(n1_O_8_0_0),
    .O_9_0_0(n1_O_9_0_0),
    .O_10_0_0(n1_O_10_0_0),
    .O_11_0_0(n1_O_11_0_0),
    .O_12_0_0(n1_O_12_0_0),
    .O_13_0_0(n1_O_13_0_0),
    .O_14_0_0(n1_O_14_0_0),
    .O_15_0_0(n1_O_15_0_0)
  );
  ShiftTS n2 ( // @[Top.scala 106:20]
    .clock(n2_clock),
    .reset(n2_reset),
    .valid_up(n2_valid_up),
    .valid_down(n2_valid_down),
    .I_0_0_0(n2_I_0_0_0),
    .I_1_0_0(n2_I_1_0_0),
    .I_2_0_0(n2_I_2_0_0),
    .I_3_0_0(n2_I_3_0_0),
    .I_4_0_0(n2_I_4_0_0),
    .I_5_0_0(n2_I_5_0_0),
    .I_6_0_0(n2_I_6_0_0),
    .I_7_0_0(n2_I_7_0_0),
    .I_8_0_0(n2_I_8_0_0),
    .I_9_0_0(n2_I_9_0_0),
    .I_10_0_0(n2_I_10_0_0),
    .I_11_0_0(n2_I_11_0_0),
    .I_12_0_0(n2_I_12_0_0),
    .I_13_0_0(n2_I_13_0_0),
    .I_14_0_0(n2_I_14_0_0),
    .I_15_0_0(n2_I_15_0_0),
    .O_0_0_0(n2_O_0_0_0),
    .O_1_0_0(n2_O_1_0_0),
    .O_2_0_0(n2_O_2_0_0),
    .O_3_0_0(n2_O_3_0_0),
    .O_4_0_0(n2_O_4_0_0),
    .O_5_0_0(n2_O_5_0_0),
    .O_6_0_0(n2_O_6_0_0),
    .O_7_0_0(n2_O_7_0_0),
    .O_8_0_0(n2_O_8_0_0),
    .O_9_0_0(n2_O_9_0_0),
    .O_10_0_0(n2_O_10_0_0),
    .O_11_0_0(n2_O_11_0_0),
    .O_12_0_0(n2_O_12_0_0),
    .O_13_0_0(n2_O_13_0_0),
    .O_14_0_0(n2_O_14_0_0),
    .O_15_0_0(n2_O_15_0_0)
  );
  ShiftTS n3 ( // @[Top.scala 109:20]
    .clock(n3_clock),
    .reset(n3_reset),
    .valid_up(n3_valid_up),
    .valid_down(n3_valid_down),
    .I_0_0_0(n3_I_0_0_0),
    .I_1_0_0(n3_I_1_0_0),
    .I_2_0_0(n3_I_2_0_0),
    .I_3_0_0(n3_I_3_0_0),
    .I_4_0_0(n3_I_4_0_0),
    .I_5_0_0(n3_I_5_0_0),
    .I_6_0_0(n3_I_6_0_0),
    .I_7_0_0(n3_I_7_0_0),
    .I_8_0_0(n3_I_8_0_0),
    .I_9_0_0(n3_I_9_0_0),
    .I_10_0_0(n3_I_10_0_0),
    .I_11_0_0(n3_I_11_0_0),
    .I_12_0_0(n3_I_12_0_0),
    .I_13_0_0(n3_I_13_0_0),
    .I_14_0_0(n3_I_14_0_0),
    .I_15_0_0(n3_I_15_0_0),
    .O_0_0_0(n3_O_0_0_0),
    .O_1_0_0(n3_O_1_0_0),
    .O_2_0_0(n3_O_2_0_0),
    .O_3_0_0(n3_O_3_0_0),
    .O_4_0_0(n3_O_4_0_0),
    .O_5_0_0(n3_O_5_0_0),
    .O_6_0_0(n3_O_6_0_0),
    .O_7_0_0(n3_O_7_0_0),
    .O_8_0_0(n3_O_8_0_0),
    .O_9_0_0(n3_O_9_0_0),
    .O_10_0_0(n3_O_10_0_0),
    .O_11_0_0(n3_O_11_0_0),
    .O_12_0_0(n3_O_12_0_0),
    .O_13_0_0(n3_O_13_0_0),
    .O_14_0_0(n3_O_14_0_0),
    .O_15_0_0(n3_O_15_0_0)
  );
  ShiftTS_2 n4 ( // @[Top.scala 112:20]
    .clock(n4_clock),
    .valid_up(n4_valid_up),
    .valid_down(n4_valid_down),
    .I_0_0_0(n4_I_0_0_0),
    .I_1_0_0(n4_I_1_0_0),
    .I_2_0_0(n4_I_2_0_0),
    .I_3_0_0(n4_I_3_0_0),
    .I_4_0_0(n4_I_4_0_0),
    .I_5_0_0(n4_I_5_0_0),
    .I_6_0_0(n4_I_6_0_0),
    .I_7_0_0(n4_I_7_0_0),
    .I_8_0_0(n4_I_8_0_0),
    .I_9_0_0(n4_I_9_0_0),
    .I_10_0_0(n4_I_10_0_0),
    .I_11_0_0(n4_I_11_0_0),
    .I_12_0_0(n4_I_12_0_0),
    .I_13_0_0(n4_I_13_0_0),
    .I_14_0_0(n4_I_14_0_0),
    .I_15_0_0(n4_I_15_0_0),
    .O_0_0_0(n4_O_0_0_0),
    .O_1_0_0(n4_O_1_0_0),
    .O_2_0_0(n4_O_2_0_0),
    .O_3_0_0(n4_O_3_0_0),
    .O_4_0_0(n4_O_4_0_0),
    .O_5_0_0(n4_O_5_0_0),
    .O_6_0_0(n4_O_6_0_0),
    .O_7_0_0(n4_O_7_0_0),
    .O_8_0_0(n4_O_8_0_0),
    .O_9_0_0(n4_O_9_0_0),
    .O_10_0_0(n4_O_10_0_0),
    .O_11_0_0(n4_O_11_0_0),
    .O_12_0_0(n4_O_12_0_0),
    .O_13_0_0(n4_O_13_0_0),
    .O_14_0_0(n4_O_14_0_0),
    .O_15_0_0(n4_O_15_0_0)
  );
  ShiftTS_2 n5 ( // @[Top.scala 115:20]
    .clock(n5_clock),
    .valid_up(n5_valid_up),
    .valid_down(n5_valid_down),
    .I_0_0_0(n5_I_0_0_0),
    .I_1_0_0(n5_I_1_0_0),
    .I_2_0_0(n5_I_2_0_0),
    .I_3_0_0(n5_I_3_0_0),
    .I_4_0_0(n5_I_4_0_0),
    .I_5_0_0(n5_I_5_0_0),
    .I_6_0_0(n5_I_6_0_0),
    .I_7_0_0(n5_I_7_0_0),
    .I_8_0_0(n5_I_8_0_0),
    .I_9_0_0(n5_I_9_0_0),
    .I_10_0_0(n5_I_10_0_0),
    .I_11_0_0(n5_I_11_0_0),
    .I_12_0_0(n5_I_12_0_0),
    .I_13_0_0(n5_I_13_0_0),
    .I_14_0_0(n5_I_14_0_0),
    .I_15_0_0(n5_I_15_0_0),
    .O_0_0_0(n5_O_0_0_0),
    .O_1_0_0(n5_O_1_0_0),
    .O_2_0_0(n5_O_2_0_0),
    .O_3_0_0(n5_O_3_0_0),
    .O_4_0_0(n5_O_4_0_0),
    .O_5_0_0(n5_O_5_0_0),
    .O_6_0_0(n5_O_6_0_0),
    .O_7_0_0(n5_O_7_0_0),
    .O_8_0_0(n5_O_8_0_0),
    .O_9_0_0(n5_O_9_0_0),
    .O_10_0_0(n5_O_10_0_0),
    .O_11_0_0(n5_O_11_0_0),
    .O_12_0_0(n5_O_12_0_0),
    .O_13_0_0(n5_O_13_0_0),
    .O_14_0_0(n5_O_14_0_0),
    .O_15_0_0(n5_O_15_0_0)
  );
  Map2T n6 ( // @[Top.scala 118:20]
    .valid_up(n6_valid_up),
    .valid_down(n6_valid_down),
    .I0_0_0_0(n6_I0_0_0_0),
    .I0_1_0_0(n6_I0_1_0_0),
    .I0_2_0_0(n6_I0_2_0_0),
    .I0_3_0_0(n6_I0_3_0_0),
    .I0_4_0_0(n6_I0_4_0_0),
    .I0_5_0_0(n6_I0_5_0_0),
    .I0_6_0_0(n6_I0_6_0_0),
    .I0_7_0_0(n6_I0_7_0_0),
    .I0_8_0_0(n6_I0_8_0_0),
    .I0_9_0_0(n6_I0_9_0_0),
    .I0_10_0_0(n6_I0_10_0_0),
    .I0_11_0_0(n6_I0_11_0_0),
    .I0_12_0_0(n6_I0_12_0_0),
    .I0_13_0_0(n6_I0_13_0_0),
    .I0_14_0_0(n6_I0_14_0_0),
    .I0_15_0_0(n6_I0_15_0_0),
    .I1_0_0_0(n6_I1_0_0_0),
    .I1_1_0_0(n6_I1_1_0_0),
    .I1_2_0_0(n6_I1_2_0_0),
    .I1_3_0_0(n6_I1_3_0_0),
    .I1_4_0_0(n6_I1_4_0_0),
    .I1_5_0_0(n6_I1_5_0_0),
    .I1_6_0_0(n6_I1_6_0_0),
    .I1_7_0_0(n6_I1_7_0_0),
    .I1_8_0_0(n6_I1_8_0_0),
    .I1_9_0_0(n6_I1_9_0_0),
    .I1_10_0_0(n6_I1_10_0_0),
    .I1_11_0_0(n6_I1_11_0_0),
    .I1_12_0_0(n6_I1_12_0_0),
    .I1_13_0_0(n6_I1_13_0_0),
    .I1_14_0_0(n6_I1_14_0_0),
    .I1_15_0_0(n6_I1_15_0_0),
    .O_0_0_0_0(n6_O_0_0_0_0),
    .O_0_0_0_1(n6_O_0_0_0_1),
    .O_1_0_0_0(n6_O_1_0_0_0),
    .O_1_0_0_1(n6_O_1_0_0_1),
    .O_2_0_0_0(n6_O_2_0_0_0),
    .O_2_0_0_1(n6_O_2_0_0_1),
    .O_3_0_0_0(n6_O_3_0_0_0),
    .O_3_0_0_1(n6_O_3_0_0_1),
    .O_4_0_0_0(n6_O_4_0_0_0),
    .O_4_0_0_1(n6_O_4_0_0_1),
    .O_5_0_0_0(n6_O_5_0_0_0),
    .O_5_0_0_1(n6_O_5_0_0_1),
    .O_6_0_0_0(n6_O_6_0_0_0),
    .O_6_0_0_1(n6_O_6_0_0_1),
    .O_7_0_0_0(n6_O_7_0_0_0),
    .O_7_0_0_1(n6_O_7_0_0_1),
    .O_8_0_0_0(n6_O_8_0_0_0),
    .O_8_0_0_1(n6_O_8_0_0_1),
    .O_9_0_0_0(n6_O_9_0_0_0),
    .O_9_0_0_1(n6_O_9_0_0_1),
    .O_10_0_0_0(n6_O_10_0_0_0),
    .O_10_0_0_1(n6_O_10_0_0_1),
    .O_11_0_0_0(n6_O_11_0_0_0),
    .O_11_0_0_1(n6_O_11_0_0_1),
    .O_12_0_0_0(n6_O_12_0_0_0),
    .O_12_0_0_1(n6_O_12_0_0_1),
    .O_13_0_0_0(n6_O_13_0_0_0),
    .O_13_0_0_1(n6_O_13_0_0_1),
    .O_14_0_0_0(n6_O_14_0_0_0),
    .O_14_0_0_1(n6_O_14_0_0_1),
    .O_15_0_0_0(n6_O_15_0_0_0),
    .O_15_0_0_1(n6_O_15_0_0_1)
  );
  Map2T_1 n19 ( // @[Top.scala 122:21]
    .valid_up(n19_valid_up),
    .valid_down(n19_valid_down),
    .I0_0_0_0_0(n19_I0_0_0_0_0),
    .I0_0_0_0_1(n19_I0_0_0_0_1),
    .I0_1_0_0_0(n19_I0_1_0_0_0),
    .I0_1_0_0_1(n19_I0_1_0_0_1),
    .I0_2_0_0_0(n19_I0_2_0_0_0),
    .I0_2_0_0_1(n19_I0_2_0_0_1),
    .I0_3_0_0_0(n19_I0_3_0_0_0),
    .I0_3_0_0_1(n19_I0_3_0_0_1),
    .I0_4_0_0_0(n19_I0_4_0_0_0),
    .I0_4_0_0_1(n19_I0_4_0_0_1),
    .I0_5_0_0_0(n19_I0_5_0_0_0),
    .I0_5_0_0_1(n19_I0_5_0_0_1),
    .I0_6_0_0_0(n19_I0_6_0_0_0),
    .I0_6_0_0_1(n19_I0_6_0_0_1),
    .I0_7_0_0_0(n19_I0_7_0_0_0),
    .I0_7_0_0_1(n19_I0_7_0_0_1),
    .I0_8_0_0_0(n19_I0_8_0_0_0),
    .I0_8_0_0_1(n19_I0_8_0_0_1),
    .I0_9_0_0_0(n19_I0_9_0_0_0),
    .I0_9_0_0_1(n19_I0_9_0_0_1),
    .I0_10_0_0_0(n19_I0_10_0_0_0),
    .I0_10_0_0_1(n19_I0_10_0_0_1),
    .I0_11_0_0_0(n19_I0_11_0_0_0),
    .I0_11_0_0_1(n19_I0_11_0_0_1),
    .I0_12_0_0_0(n19_I0_12_0_0_0),
    .I0_12_0_0_1(n19_I0_12_0_0_1),
    .I0_13_0_0_0(n19_I0_13_0_0_0),
    .I0_13_0_0_1(n19_I0_13_0_0_1),
    .I0_14_0_0_0(n19_I0_14_0_0_0),
    .I0_14_0_0_1(n19_I0_14_0_0_1),
    .I0_15_0_0_0(n19_I0_15_0_0_0),
    .I0_15_0_0_1(n19_I0_15_0_0_1),
    .I1_0_0_0(n19_I1_0_0_0),
    .I1_1_0_0(n19_I1_1_0_0),
    .I1_2_0_0(n19_I1_2_0_0),
    .I1_3_0_0(n19_I1_3_0_0),
    .I1_4_0_0(n19_I1_4_0_0),
    .I1_5_0_0(n19_I1_5_0_0),
    .I1_6_0_0(n19_I1_6_0_0),
    .I1_7_0_0(n19_I1_7_0_0),
    .I1_8_0_0(n19_I1_8_0_0),
    .I1_9_0_0(n19_I1_9_0_0),
    .I1_10_0_0(n19_I1_10_0_0),
    .I1_11_0_0(n19_I1_11_0_0),
    .I1_12_0_0(n19_I1_12_0_0),
    .I1_13_0_0(n19_I1_13_0_0),
    .I1_14_0_0(n19_I1_14_0_0),
    .I1_15_0_0(n19_I1_15_0_0),
    .O_0_0_0_0(n19_O_0_0_0_0),
    .O_0_0_0_1(n19_O_0_0_0_1),
    .O_0_0_0_2(n19_O_0_0_0_2),
    .O_1_0_0_0(n19_O_1_0_0_0),
    .O_1_0_0_1(n19_O_1_0_0_1),
    .O_1_0_0_2(n19_O_1_0_0_2),
    .O_2_0_0_0(n19_O_2_0_0_0),
    .O_2_0_0_1(n19_O_2_0_0_1),
    .O_2_0_0_2(n19_O_2_0_0_2),
    .O_3_0_0_0(n19_O_3_0_0_0),
    .O_3_0_0_1(n19_O_3_0_0_1),
    .O_3_0_0_2(n19_O_3_0_0_2),
    .O_4_0_0_0(n19_O_4_0_0_0),
    .O_4_0_0_1(n19_O_4_0_0_1),
    .O_4_0_0_2(n19_O_4_0_0_2),
    .O_5_0_0_0(n19_O_5_0_0_0),
    .O_5_0_0_1(n19_O_5_0_0_1),
    .O_5_0_0_2(n19_O_5_0_0_2),
    .O_6_0_0_0(n19_O_6_0_0_0),
    .O_6_0_0_1(n19_O_6_0_0_1),
    .O_6_0_0_2(n19_O_6_0_0_2),
    .O_7_0_0_0(n19_O_7_0_0_0),
    .O_7_0_0_1(n19_O_7_0_0_1),
    .O_7_0_0_2(n19_O_7_0_0_2),
    .O_8_0_0_0(n19_O_8_0_0_0),
    .O_8_0_0_1(n19_O_8_0_0_1),
    .O_8_0_0_2(n19_O_8_0_0_2),
    .O_9_0_0_0(n19_O_9_0_0_0),
    .O_9_0_0_1(n19_O_9_0_0_1),
    .O_9_0_0_2(n19_O_9_0_0_2),
    .O_10_0_0_0(n19_O_10_0_0_0),
    .O_10_0_0_1(n19_O_10_0_0_1),
    .O_10_0_0_2(n19_O_10_0_0_2),
    .O_11_0_0_0(n19_O_11_0_0_0),
    .O_11_0_0_1(n19_O_11_0_0_1),
    .O_11_0_0_2(n19_O_11_0_0_2),
    .O_12_0_0_0(n19_O_12_0_0_0),
    .O_12_0_0_1(n19_O_12_0_0_1),
    .O_12_0_0_2(n19_O_12_0_0_2),
    .O_13_0_0_0(n19_O_13_0_0_0),
    .O_13_0_0_1(n19_O_13_0_0_1),
    .O_13_0_0_2(n19_O_13_0_0_2),
    .O_14_0_0_0(n19_O_14_0_0_0),
    .O_14_0_0_1(n19_O_14_0_0_1),
    .O_14_0_0_2(n19_O_14_0_0_2),
    .O_15_0_0_0(n19_O_15_0_0_0),
    .O_15_0_0_1(n19_O_15_0_0_1),
    .O_15_0_0_2(n19_O_15_0_0_2)
  );
  MapT n40 ( // @[Top.scala 126:21]
    .valid_up(n40_valid_up),
    .valid_down(n40_valid_down),
    .I_0_0_0_0(n40_I_0_0_0_0),
    .I_0_0_0_1(n40_I_0_0_0_1),
    .I_0_0_0_2(n40_I_0_0_0_2),
    .I_1_0_0_0(n40_I_1_0_0_0),
    .I_1_0_0_1(n40_I_1_0_0_1),
    .I_1_0_0_2(n40_I_1_0_0_2),
    .I_2_0_0_0(n40_I_2_0_0_0),
    .I_2_0_0_1(n40_I_2_0_0_1),
    .I_2_0_0_2(n40_I_2_0_0_2),
    .I_3_0_0_0(n40_I_3_0_0_0),
    .I_3_0_0_1(n40_I_3_0_0_1),
    .I_3_0_0_2(n40_I_3_0_0_2),
    .I_4_0_0_0(n40_I_4_0_0_0),
    .I_4_0_0_1(n40_I_4_0_0_1),
    .I_4_0_0_2(n40_I_4_0_0_2),
    .I_5_0_0_0(n40_I_5_0_0_0),
    .I_5_0_0_1(n40_I_5_0_0_1),
    .I_5_0_0_2(n40_I_5_0_0_2),
    .I_6_0_0_0(n40_I_6_0_0_0),
    .I_6_0_0_1(n40_I_6_0_0_1),
    .I_6_0_0_2(n40_I_6_0_0_2),
    .I_7_0_0_0(n40_I_7_0_0_0),
    .I_7_0_0_1(n40_I_7_0_0_1),
    .I_7_0_0_2(n40_I_7_0_0_2),
    .I_8_0_0_0(n40_I_8_0_0_0),
    .I_8_0_0_1(n40_I_8_0_0_1),
    .I_8_0_0_2(n40_I_8_0_0_2),
    .I_9_0_0_0(n40_I_9_0_0_0),
    .I_9_0_0_1(n40_I_9_0_0_1),
    .I_9_0_0_2(n40_I_9_0_0_2),
    .I_10_0_0_0(n40_I_10_0_0_0),
    .I_10_0_0_1(n40_I_10_0_0_1),
    .I_10_0_0_2(n40_I_10_0_0_2),
    .I_11_0_0_0(n40_I_11_0_0_0),
    .I_11_0_0_1(n40_I_11_0_0_1),
    .I_11_0_0_2(n40_I_11_0_0_2),
    .I_12_0_0_0(n40_I_12_0_0_0),
    .I_12_0_0_1(n40_I_12_0_0_1),
    .I_12_0_0_2(n40_I_12_0_0_2),
    .I_13_0_0_0(n40_I_13_0_0_0),
    .I_13_0_0_1(n40_I_13_0_0_1),
    .I_13_0_0_2(n40_I_13_0_0_2),
    .I_14_0_0_0(n40_I_14_0_0_0),
    .I_14_0_0_1(n40_I_14_0_0_1),
    .I_14_0_0_2(n40_I_14_0_0_2),
    .I_15_0_0_0(n40_I_15_0_0_0),
    .I_15_0_0_1(n40_I_15_0_0_1),
    .I_15_0_0_2(n40_I_15_0_0_2),
    .O_0_0_0(n40_O_0_0_0),
    .O_0_0_1(n40_O_0_0_1),
    .O_0_0_2(n40_O_0_0_2),
    .O_1_0_0(n40_O_1_0_0),
    .O_1_0_1(n40_O_1_0_1),
    .O_1_0_2(n40_O_1_0_2),
    .O_2_0_0(n40_O_2_0_0),
    .O_2_0_1(n40_O_2_0_1),
    .O_2_0_2(n40_O_2_0_2),
    .O_3_0_0(n40_O_3_0_0),
    .O_3_0_1(n40_O_3_0_1),
    .O_3_0_2(n40_O_3_0_2),
    .O_4_0_0(n40_O_4_0_0),
    .O_4_0_1(n40_O_4_0_1),
    .O_4_0_2(n40_O_4_0_2),
    .O_5_0_0(n40_O_5_0_0),
    .O_5_0_1(n40_O_5_0_1),
    .O_5_0_2(n40_O_5_0_2),
    .O_6_0_0(n40_O_6_0_0),
    .O_6_0_1(n40_O_6_0_1),
    .O_6_0_2(n40_O_6_0_2),
    .O_7_0_0(n40_O_7_0_0),
    .O_7_0_1(n40_O_7_0_1),
    .O_7_0_2(n40_O_7_0_2),
    .O_8_0_0(n40_O_8_0_0),
    .O_8_0_1(n40_O_8_0_1),
    .O_8_0_2(n40_O_8_0_2),
    .O_9_0_0(n40_O_9_0_0),
    .O_9_0_1(n40_O_9_0_1),
    .O_9_0_2(n40_O_9_0_2),
    .O_10_0_0(n40_O_10_0_0),
    .O_10_0_1(n40_O_10_0_1),
    .O_10_0_2(n40_O_10_0_2),
    .O_11_0_0(n40_O_11_0_0),
    .O_11_0_1(n40_O_11_0_1),
    .O_11_0_2(n40_O_11_0_2),
    .O_12_0_0(n40_O_12_0_0),
    .O_12_0_1(n40_O_12_0_1),
    .O_12_0_2(n40_O_12_0_2),
    .O_13_0_0(n40_O_13_0_0),
    .O_13_0_1(n40_O_13_0_1),
    .O_13_0_2(n40_O_13_0_2),
    .O_14_0_0(n40_O_14_0_0),
    .O_14_0_1(n40_O_14_0_1),
    .O_14_0_2(n40_O_14_0_2),
    .O_15_0_0(n40_O_15_0_0),
    .O_15_0_1(n40_O_15_0_1),
    .O_15_0_2(n40_O_15_0_2)
  );
  ShiftTS_2 n41 ( // @[Top.scala 129:21]
    .clock(n41_clock),
    .valid_up(n41_valid_up),
    .valid_down(n41_valid_down),
    .I_0_0_0(n41_I_0_0_0),
    .I_1_0_0(n41_I_1_0_0),
    .I_2_0_0(n41_I_2_0_0),
    .I_3_0_0(n41_I_3_0_0),
    .I_4_0_0(n41_I_4_0_0),
    .I_5_0_0(n41_I_5_0_0),
    .I_6_0_0(n41_I_6_0_0),
    .I_7_0_0(n41_I_7_0_0),
    .I_8_0_0(n41_I_8_0_0),
    .I_9_0_0(n41_I_9_0_0),
    .I_10_0_0(n41_I_10_0_0),
    .I_11_0_0(n41_I_11_0_0),
    .I_12_0_0(n41_I_12_0_0),
    .I_13_0_0(n41_I_13_0_0),
    .I_14_0_0(n41_I_14_0_0),
    .I_15_0_0(n41_I_15_0_0),
    .O_0_0_0(n41_O_0_0_0),
    .O_1_0_0(n41_O_1_0_0),
    .O_2_0_0(n41_O_2_0_0),
    .O_3_0_0(n41_O_3_0_0),
    .O_4_0_0(n41_O_4_0_0),
    .O_5_0_0(n41_O_5_0_0),
    .O_6_0_0(n41_O_6_0_0),
    .O_7_0_0(n41_O_7_0_0),
    .O_8_0_0(n41_O_8_0_0),
    .O_9_0_0(n41_O_9_0_0),
    .O_10_0_0(n41_O_10_0_0),
    .O_11_0_0(n41_O_11_0_0),
    .O_12_0_0(n41_O_12_0_0),
    .O_13_0_0(n41_O_13_0_0),
    .O_14_0_0(n41_O_14_0_0),
    .O_15_0_0(n41_O_15_0_0)
  );
  ShiftTS_2 n42 ( // @[Top.scala 132:21]
    .clock(n42_clock),
    .valid_up(n42_valid_up),
    .valid_down(n42_valid_down),
    .I_0_0_0(n42_I_0_0_0),
    .I_1_0_0(n42_I_1_0_0),
    .I_2_0_0(n42_I_2_0_0),
    .I_3_0_0(n42_I_3_0_0),
    .I_4_0_0(n42_I_4_0_0),
    .I_5_0_0(n42_I_5_0_0),
    .I_6_0_0(n42_I_6_0_0),
    .I_7_0_0(n42_I_7_0_0),
    .I_8_0_0(n42_I_8_0_0),
    .I_9_0_0(n42_I_9_0_0),
    .I_10_0_0(n42_I_10_0_0),
    .I_11_0_0(n42_I_11_0_0),
    .I_12_0_0(n42_I_12_0_0),
    .I_13_0_0(n42_I_13_0_0),
    .I_14_0_0(n42_I_14_0_0),
    .I_15_0_0(n42_I_15_0_0),
    .O_0_0_0(n42_O_0_0_0),
    .O_1_0_0(n42_O_1_0_0),
    .O_2_0_0(n42_O_2_0_0),
    .O_3_0_0(n42_O_3_0_0),
    .O_4_0_0(n42_O_4_0_0),
    .O_5_0_0(n42_O_5_0_0),
    .O_6_0_0(n42_O_6_0_0),
    .O_7_0_0(n42_O_7_0_0),
    .O_8_0_0(n42_O_8_0_0),
    .O_9_0_0(n42_O_9_0_0),
    .O_10_0_0(n42_O_10_0_0),
    .O_11_0_0(n42_O_11_0_0),
    .O_12_0_0(n42_O_12_0_0),
    .O_13_0_0(n42_O_13_0_0),
    .O_14_0_0(n42_O_14_0_0),
    .O_15_0_0(n42_O_15_0_0)
  );
  Map2T n43 ( // @[Top.scala 135:21]
    .valid_up(n43_valid_up),
    .valid_down(n43_valid_down),
    .I0_0_0_0(n43_I0_0_0_0),
    .I0_1_0_0(n43_I0_1_0_0),
    .I0_2_0_0(n43_I0_2_0_0),
    .I0_3_0_0(n43_I0_3_0_0),
    .I0_4_0_0(n43_I0_4_0_0),
    .I0_5_0_0(n43_I0_5_0_0),
    .I0_6_0_0(n43_I0_6_0_0),
    .I0_7_0_0(n43_I0_7_0_0),
    .I0_8_0_0(n43_I0_8_0_0),
    .I0_9_0_0(n43_I0_9_0_0),
    .I0_10_0_0(n43_I0_10_0_0),
    .I0_11_0_0(n43_I0_11_0_0),
    .I0_12_0_0(n43_I0_12_0_0),
    .I0_13_0_0(n43_I0_13_0_0),
    .I0_14_0_0(n43_I0_14_0_0),
    .I0_15_0_0(n43_I0_15_0_0),
    .I1_0_0_0(n43_I1_0_0_0),
    .I1_1_0_0(n43_I1_1_0_0),
    .I1_2_0_0(n43_I1_2_0_0),
    .I1_3_0_0(n43_I1_3_0_0),
    .I1_4_0_0(n43_I1_4_0_0),
    .I1_5_0_0(n43_I1_5_0_0),
    .I1_6_0_0(n43_I1_6_0_0),
    .I1_7_0_0(n43_I1_7_0_0),
    .I1_8_0_0(n43_I1_8_0_0),
    .I1_9_0_0(n43_I1_9_0_0),
    .I1_10_0_0(n43_I1_10_0_0),
    .I1_11_0_0(n43_I1_11_0_0),
    .I1_12_0_0(n43_I1_12_0_0),
    .I1_13_0_0(n43_I1_13_0_0),
    .I1_14_0_0(n43_I1_14_0_0),
    .I1_15_0_0(n43_I1_15_0_0),
    .O_0_0_0_0(n43_O_0_0_0_0),
    .O_0_0_0_1(n43_O_0_0_0_1),
    .O_1_0_0_0(n43_O_1_0_0_0),
    .O_1_0_0_1(n43_O_1_0_0_1),
    .O_2_0_0_0(n43_O_2_0_0_0),
    .O_2_0_0_1(n43_O_2_0_0_1),
    .O_3_0_0_0(n43_O_3_0_0_0),
    .O_3_0_0_1(n43_O_3_0_0_1),
    .O_4_0_0_0(n43_O_4_0_0_0),
    .O_4_0_0_1(n43_O_4_0_0_1),
    .O_5_0_0_0(n43_O_5_0_0_0),
    .O_5_0_0_1(n43_O_5_0_0_1),
    .O_6_0_0_0(n43_O_6_0_0_0),
    .O_6_0_0_1(n43_O_6_0_0_1),
    .O_7_0_0_0(n43_O_7_0_0_0),
    .O_7_0_0_1(n43_O_7_0_0_1),
    .O_8_0_0_0(n43_O_8_0_0_0),
    .O_8_0_0_1(n43_O_8_0_0_1),
    .O_9_0_0_0(n43_O_9_0_0_0),
    .O_9_0_0_1(n43_O_9_0_0_1),
    .O_10_0_0_0(n43_O_10_0_0_0),
    .O_10_0_0_1(n43_O_10_0_0_1),
    .O_11_0_0_0(n43_O_11_0_0_0),
    .O_11_0_0_1(n43_O_11_0_0_1),
    .O_12_0_0_0(n43_O_12_0_0_0),
    .O_12_0_0_1(n43_O_12_0_0_1),
    .O_13_0_0_0(n43_O_13_0_0_0),
    .O_13_0_0_1(n43_O_13_0_0_1),
    .O_14_0_0_0(n43_O_14_0_0_0),
    .O_14_0_0_1(n43_O_14_0_0_1),
    .O_15_0_0_0(n43_O_15_0_0_0),
    .O_15_0_0_1(n43_O_15_0_0_1)
  );
  Map2T_1 n56 ( // @[Top.scala 139:21]
    .valid_up(n56_valid_up),
    .valid_down(n56_valid_down),
    .I0_0_0_0_0(n56_I0_0_0_0_0),
    .I0_0_0_0_1(n56_I0_0_0_0_1),
    .I0_1_0_0_0(n56_I0_1_0_0_0),
    .I0_1_0_0_1(n56_I0_1_0_0_1),
    .I0_2_0_0_0(n56_I0_2_0_0_0),
    .I0_2_0_0_1(n56_I0_2_0_0_1),
    .I0_3_0_0_0(n56_I0_3_0_0_0),
    .I0_3_0_0_1(n56_I0_3_0_0_1),
    .I0_4_0_0_0(n56_I0_4_0_0_0),
    .I0_4_0_0_1(n56_I0_4_0_0_1),
    .I0_5_0_0_0(n56_I0_5_0_0_0),
    .I0_5_0_0_1(n56_I0_5_0_0_1),
    .I0_6_0_0_0(n56_I0_6_0_0_0),
    .I0_6_0_0_1(n56_I0_6_0_0_1),
    .I0_7_0_0_0(n56_I0_7_0_0_0),
    .I0_7_0_0_1(n56_I0_7_0_0_1),
    .I0_8_0_0_0(n56_I0_8_0_0_0),
    .I0_8_0_0_1(n56_I0_8_0_0_1),
    .I0_9_0_0_0(n56_I0_9_0_0_0),
    .I0_9_0_0_1(n56_I0_9_0_0_1),
    .I0_10_0_0_0(n56_I0_10_0_0_0),
    .I0_10_0_0_1(n56_I0_10_0_0_1),
    .I0_11_0_0_0(n56_I0_11_0_0_0),
    .I0_11_0_0_1(n56_I0_11_0_0_1),
    .I0_12_0_0_0(n56_I0_12_0_0_0),
    .I0_12_0_0_1(n56_I0_12_0_0_1),
    .I0_13_0_0_0(n56_I0_13_0_0_0),
    .I0_13_0_0_1(n56_I0_13_0_0_1),
    .I0_14_0_0_0(n56_I0_14_0_0_0),
    .I0_14_0_0_1(n56_I0_14_0_0_1),
    .I0_15_0_0_0(n56_I0_15_0_0_0),
    .I0_15_0_0_1(n56_I0_15_0_0_1),
    .I1_0_0_0(n56_I1_0_0_0),
    .I1_1_0_0(n56_I1_1_0_0),
    .I1_2_0_0(n56_I1_2_0_0),
    .I1_3_0_0(n56_I1_3_0_0),
    .I1_4_0_0(n56_I1_4_0_0),
    .I1_5_0_0(n56_I1_5_0_0),
    .I1_6_0_0(n56_I1_6_0_0),
    .I1_7_0_0(n56_I1_7_0_0),
    .I1_8_0_0(n56_I1_8_0_0),
    .I1_9_0_0(n56_I1_9_0_0),
    .I1_10_0_0(n56_I1_10_0_0),
    .I1_11_0_0(n56_I1_11_0_0),
    .I1_12_0_0(n56_I1_12_0_0),
    .I1_13_0_0(n56_I1_13_0_0),
    .I1_14_0_0(n56_I1_14_0_0),
    .I1_15_0_0(n56_I1_15_0_0),
    .O_0_0_0_0(n56_O_0_0_0_0),
    .O_0_0_0_1(n56_O_0_0_0_1),
    .O_0_0_0_2(n56_O_0_0_0_2),
    .O_1_0_0_0(n56_O_1_0_0_0),
    .O_1_0_0_1(n56_O_1_0_0_1),
    .O_1_0_0_2(n56_O_1_0_0_2),
    .O_2_0_0_0(n56_O_2_0_0_0),
    .O_2_0_0_1(n56_O_2_0_0_1),
    .O_2_0_0_2(n56_O_2_0_0_2),
    .O_3_0_0_0(n56_O_3_0_0_0),
    .O_3_0_0_1(n56_O_3_0_0_1),
    .O_3_0_0_2(n56_O_3_0_0_2),
    .O_4_0_0_0(n56_O_4_0_0_0),
    .O_4_0_0_1(n56_O_4_0_0_1),
    .O_4_0_0_2(n56_O_4_0_0_2),
    .O_5_0_0_0(n56_O_5_0_0_0),
    .O_5_0_0_1(n56_O_5_0_0_1),
    .O_5_0_0_2(n56_O_5_0_0_2),
    .O_6_0_0_0(n56_O_6_0_0_0),
    .O_6_0_0_1(n56_O_6_0_0_1),
    .O_6_0_0_2(n56_O_6_0_0_2),
    .O_7_0_0_0(n56_O_7_0_0_0),
    .O_7_0_0_1(n56_O_7_0_0_1),
    .O_7_0_0_2(n56_O_7_0_0_2),
    .O_8_0_0_0(n56_O_8_0_0_0),
    .O_8_0_0_1(n56_O_8_0_0_1),
    .O_8_0_0_2(n56_O_8_0_0_2),
    .O_9_0_0_0(n56_O_9_0_0_0),
    .O_9_0_0_1(n56_O_9_0_0_1),
    .O_9_0_0_2(n56_O_9_0_0_2),
    .O_10_0_0_0(n56_O_10_0_0_0),
    .O_10_0_0_1(n56_O_10_0_0_1),
    .O_10_0_0_2(n56_O_10_0_0_2),
    .O_11_0_0_0(n56_O_11_0_0_0),
    .O_11_0_0_1(n56_O_11_0_0_1),
    .O_11_0_0_2(n56_O_11_0_0_2),
    .O_12_0_0_0(n56_O_12_0_0_0),
    .O_12_0_0_1(n56_O_12_0_0_1),
    .O_12_0_0_2(n56_O_12_0_0_2),
    .O_13_0_0_0(n56_O_13_0_0_0),
    .O_13_0_0_1(n56_O_13_0_0_1),
    .O_13_0_0_2(n56_O_13_0_0_2),
    .O_14_0_0_0(n56_O_14_0_0_0),
    .O_14_0_0_1(n56_O_14_0_0_1),
    .O_14_0_0_2(n56_O_14_0_0_2),
    .O_15_0_0_0(n56_O_15_0_0_0),
    .O_15_0_0_1(n56_O_15_0_0_1),
    .O_15_0_0_2(n56_O_15_0_0_2)
  );
  MapT n77 ( // @[Top.scala 143:21]
    .valid_up(n77_valid_up),
    .valid_down(n77_valid_down),
    .I_0_0_0_0(n77_I_0_0_0_0),
    .I_0_0_0_1(n77_I_0_0_0_1),
    .I_0_0_0_2(n77_I_0_0_0_2),
    .I_1_0_0_0(n77_I_1_0_0_0),
    .I_1_0_0_1(n77_I_1_0_0_1),
    .I_1_0_0_2(n77_I_1_0_0_2),
    .I_2_0_0_0(n77_I_2_0_0_0),
    .I_2_0_0_1(n77_I_2_0_0_1),
    .I_2_0_0_2(n77_I_2_0_0_2),
    .I_3_0_0_0(n77_I_3_0_0_0),
    .I_3_0_0_1(n77_I_3_0_0_1),
    .I_3_0_0_2(n77_I_3_0_0_2),
    .I_4_0_0_0(n77_I_4_0_0_0),
    .I_4_0_0_1(n77_I_4_0_0_1),
    .I_4_0_0_2(n77_I_4_0_0_2),
    .I_5_0_0_0(n77_I_5_0_0_0),
    .I_5_0_0_1(n77_I_5_0_0_1),
    .I_5_0_0_2(n77_I_5_0_0_2),
    .I_6_0_0_0(n77_I_6_0_0_0),
    .I_6_0_0_1(n77_I_6_0_0_1),
    .I_6_0_0_2(n77_I_6_0_0_2),
    .I_7_0_0_0(n77_I_7_0_0_0),
    .I_7_0_0_1(n77_I_7_0_0_1),
    .I_7_0_0_2(n77_I_7_0_0_2),
    .I_8_0_0_0(n77_I_8_0_0_0),
    .I_8_0_0_1(n77_I_8_0_0_1),
    .I_8_0_0_2(n77_I_8_0_0_2),
    .I_9_0_0_0(n77_I_9_0_0_0),
    .I_9_0_0_1(n77_I_9_0_0_1),
    .I_9_0_0_2(n77_I_9_0_0_2),
    .I_10_0_0_0(n77_I_10_0_0_0),
    .I_10_0_0_1(n77_I_10_0_0_1),
    .I_10_0_0_2(n77_I_10_0_0_2),
    .I_11_0_0_0(n77_I_11_0_0_0),
    .I_11_0_0_1(n77_I_11_0_0_1),
    .I_11_0_0_2(n77_I_11_0_0_2),
    .I_12_0_0_0(n77_I_12_0_0_0),
    .I_12_0_0_1(n77_I_12_0_0_1),
    .I_12_0_0_2(n77_I_12_0_0_2),
    .I_13_0_0_0(n77_I_13_0_0_0),
    .I_13_0_0_1(n77_I_13_0_0_1),
    .I_13_0_0_2(n77_I_13_0_0_2),
    .I_14_0_0_0(n77_I_14_0_0_0),
    .I_14_0_0_1(n77_I_14_0_0_1),
    .I_14_0_0_2(n77_I_14_0_0_2),
    .I_15_0_0_0(n77_I_15_0_0_0),
    .I_15_0_0_1(n77_I_15_0_0_1),
    .I_15_0_0_2(n77_I_15_0_0_2),
    .O_0_0_0(n77_O_0_0_0),
    .O_0_0_1(n77_O_0_0_1),
    .O_0_0_2(n77_O_0_0_2),
    .O_1_0_0(n77_O_1_0_0),
    .O_1_0_1(n77_O_1_0_1),
    .O_1_0_2(n77_O_1_0_2),
    .O_2_0_0(n77_O_2_0_0),
    .O_2_0_1(n77_O_2_0_1),
    .O_2_0_2(n77_O_2_0_2),
    .O_3_0_0(n77_O_3_0_0),
    .O_3_0_1(n77_O_3_0_1),
    .O_3_0_2(n77_O_3_0_2),
    .O_4_0_0(n77_O_4_0_0),
    .O_4_0_1(n77_O_4_0_1),
    .O_4_0_2(n77_O_4_0_2),
    .O_5_0_0(n77_O_5_0_0),
    .O_5_0_1(n77_O_5_0_1),
    .O_5_0_2(n77_O_5_0_2),
    .O_6_0_0(n77_O_6_0_0),
    .O_6_0_1(n77_O_6_0_1),
    .O_6_0_2(n77_O_6_0_2),
    .O_7_0_0(n77_O_7_0_0),
    .O_7_0_1(n77_O_7_0_1),
    .O_7_0_2(n77_O_7_0_2),
    .O_8_0_0(n77_O_8_0_0),
    .O_8_0_1(n77_O_8_0_1),
    .O_8_0_2(n77_O_8_0_2),
    .O_9_0_0(n77_O_9_0_0),
    .O_9_0_1(n77_O_9_0_1),
    .O_9_0_2(n77_O_9_0_2),
    .O_10_0_0(n77_O_10_0_0),
    .O_10_0_1(n77_O_10_0_1),
    .O_10_0_2(n77_O_10_0_2),
    .O_11_0_0(n77_O_11_0_0),
    .O_11_0_1(n77_O_11_0_1),
    .O_11_0_2(n77_O_11_0_2),
    .O_12_0_0(n77_O_12_0_0),
    .O_12_0_1(n77_O_12_0_1),
    .O_12_0_2(n77_O_12_0_2),
    .O_13_0_0(n77_O_13_0_0),
    .O_13_0_1(n77_O_13_0_1),
    .O_13_0_2(n77_O_13_0_2),
    .O_14_0_0(n77_O_14_0_0),
    .O_14_0_1(n77_O_14_0_1),
    .O_14_0_2(n77_O_14_0_2),
    .O_15_0_0(n77_O_15_0_0),
    .O_15_0_1(n77_O_15_0_1),
    .O_15_0_2(n77_O_15_0_2)
  );
  Map2T_4 n78 ( // @[Top.scala 146:21]
    .valid_up(n78_valid_up),
    .valid_down(n78_valid_down),
    .I0_0_0_0(n78_I0_0_0_0),
    .I0_0_0_1(n78_I0_0_0_1),
    .I0_0_0_2(n78_I0_0_0_2),
    .I0_1_0_0(n78_I0_1_0_0),
    .I0_1_0_1(n78_I0_1_0_1),
    .I0_1_0_2(n78_I0_1_0_2),
    .I0_2_0_0(n78_I0_2_0_0),
    .I0_2_0_1(n78_I0_2_0_1),
    .I0_2_0_2(n78_I0_2_0_2),
    .I0_3_0_0(n78_I0_3_0_0),
    .I0_3_0_1(n78_I0_3_0_1),
    .I0_3_0_2(n78_I0_3_0_2),
    .I0_4_0_0(n78_I0_4_0_0),
    .I0_4_0_1(n78_I0_4_0_1),
    .I0_4_0_2(n78_I0_4_0_2),
    .I0_5_0_0(n78_I0_5_0_0),
    .I0_5_0_1(n78_I0_5_0_1),
    .I0_5_0_2(n78_I0_5_0_2),
    .I0_6_0_0(n78_I0_6_0_0),
    .I0_6_0_1(n78_I0_6_0_1),
    .I0_6_0_2(n78_I0_6_0_2),
    .I0_7_0_0(n78_I0_7_0_0),
    .I0_7_0_1(n78_I0_7_0_1),
    .I0_7_0_2(n78_I0_7_0_2),
    .I0_8_0_0(n78_I0_8_0_0),
    .I0_8_0_1(n78_I0_8_0_1),
    .I0_8_0_2(n78_I0_8_0_2),
    .I0_9_0_0(n78_I0_9_0_0),
    .I0_9_0_1(n78_I0_9_0_1),
    .I0_9_0_2(n78_I0_9_0_2),
    .I0_10_0_0(n78_I0_10_0_0),
    .I0_10_0_1(n78_I0_10_0_1),
    .I0_10_0_2(n78_I0_10_0_2),
    .I0_11_0_0(n78_I0_11_0_0),
    .I0_11_0_1(n78_I0_11_0_1),
    .I0_11_0_2(n78_I0_11_0_2),
    .I0_12_0_0(n78_I0_12_0_0),
    .I0_12_0_1(n78_I0_12_0_1),
    .I0_12_0_2(n78_I0_12_0_2),
    .I0_13_0_0(n78_I0_13_0_0),
    .I0_13_0_1(n78_I0_13_0_1),
    .I0_13_0_2(n78_I0_13_0_2),
    .I0_14_0_0(n78_I0_14_0_0),
    .I0_14_0_1(n78_I0_14_0_1),
    .I0_14_0_2(n78_I0_14_0_2),
    .I0_15_0_0(n78_I0_15_0_0),
    .I0_15_0_1(n78_I0_15_0_1),
    .I0_15_0_2(n78_I0_15_0_2),
    .I1_0_0_0(n78_I1_0_0_0),
    .I1_0_0_1(n78_I1_0_0_1),
    .I1_0_0_2(n78_I1_0_0_2),
    .I1_1_0_0(n78_I1_1_0_0),
    .I1_1_0_1(n78_I1_1_0_1),
    .I1_1_0_2(n78_I1_1_0_2),
    .I1_2_0_0(n78_I1_2_0_0),
    .I1_2_0_1(n78_I1_2_0_1),
    .I1_2_0_2(n78_I1_2_0_2),
    .I1_3_0_0(n78_I1_3_0_0),
    .I1_3_0_1(n78_I1_3_0_1),
    .I1_3_0_2(n78_I1_3_0_2),
    .I1_4_0_0(n78_I1_4_0_0),
    .I1_4_0_1(n78_I1_4_0_1),
    .I1_4_0_2(n78_I1_4_0_2),
    .I1_5_0_0(n78_I1_5_0_0),
    .I1_5_0_1(n78_I1_5_0_1),
    .I1_5_0_2(n78_I1_5_0_2),
    .I1_6_0_0(n78_I1_6_0_0),
    .I1_6_0_1(n78_I1_6_0_1),
    .I1_6_0_2(n78_I1_6_0_2),
    .I1_7_0_0(n78_I1_7_0_0),
    .I1_7_0_1(n78_I1_7_0_1),
    .I1_7_0_2(n78_I1_7_0_2),
    .I1_8_0_0(n78_I1_8_0_0),
    .I1_8_0_1(n78_I1_8_0_1),
    .I1_8_0_2(n78_I1_8_0_2),
    .I1_9_0_0(n78_I1_9_0_0),
    .I1_9_0_1(n78_I1_9_0_1),
    .I1_9_0_2(n78_I1_9_0_2),
    .I1_10_0_0(n78_I1_10_0_0),
    .I1_10_0_1(n78_I1_10_0_1),
    .I1_10_0_2(n78_I1_10_0_2),
    .I1_11_0_0(n78_I1_11_0_0),
    .I1_11_0_1(n78_I1_11_0_1),
    .I1_11_0_2(n78_I1_11_0_2),
    .I1_12_0_0(n78_I1_12_0_0),
    .I1_12_0_1(n78_I1_12_0_1),
    .I1_12_0_2(n78_I1_12_0_2),
    .I1_13_0_0(n78_I1_13_0_0),
    .I1_13_0_1(n78_I1_13_0_1),
    .I1_13_0_2(n78_I1_13_0_2),
    .I1_14_0_0(n78_I1_14_0_0),
    .I1_14_0_1(n78_I1_14_0_1),
    .I1_14_0_2(n78_I1_14_0_2),
    .I1_15_0_0(n78_I1_15_0_0),
    .I1_15_0_1(n78_I1_15_0_1),
    .I1_15_0_2(n78_I1_15_0_2),
    .O_0_0_0_0(n78_O_0_0_0_0),
    .O_0_0_0_1(n78_O_0_0_0_1),
    .O_0_0_0_2(n78_O_0_0_0_2),
    .O_0_0_1_0(n78_O_0_0_1_0),
    .O_0_0_1_1(n78_O_0_0_1_1),
    .O_0_0_1_2(n78_O_0_0_1_2),
    .O_1_0_0_0(n78_O_1_0_0_0),
    .O_1_0_0_1(n78_O_1_0_0_1),
    .O_1_0_0_2(n78_O_1_0_0_2),
    .O_1_0_1_0(n78_O_1_0_1_0),
    .O_1_0_1_1(n78_O_1_0_1_1),
    .O_1_0_1_2(n78_O_1_0_1_2),
    .O_2_0_0_0(n78_O_2_0_0_0),
    .O_2_0_0_1(n78_O_2_0_0_1),
    .O_2_0_0_2(n78_O_2_0_0_2),
    .O_2_0_1_0(n78_O_2_0_1_0),
    .O_2_0_1_1(n78_O_2_0_1_1),
    .O_2_0_1_2(n78_O_2_0_1_2),
    .O_3_0_0_0(n78_O_3_0_0_0),
    .O_3_0_0_1(n78_O_3_0_0_1),
    .O_3_0_0_2(n78_O_3_0_0_2),
    .O_3_0_1_0(n78_O_3_0_1_0),
    .O_3_0_1_1(n78_O_3_0_1_1),
    .O_3_0_1_2(n78_O_3_0_1_2),
    .O_4_0_0_0(n78_O_4_0_0_0),
    .O_4_0_0_1(n78_O_4_0_0_1),
    .O_4_0_0_2(n78_O_4_0_0_2),
    .O_4_0_1_0(n78_O_4_0_1_0),
    .O_4_0_1_1(n78_O_4_0_1_1),
    .O_4_0_1_2(n78_O_4_0_1_2),
    .O_5_0_0_0(n78_O_5_0_0_0),
    .O_5_0_0_1(n78_O_5_0_0_1),
    .O_5_0_0_2(n78_O_5_0_0_2),
    .O_5_0_1_0(n78_O_5_0_1_0),
    .O_5_0_1_1(n78_O_5_0_1_1),
    .O_5_0_1_2(n78_O_5_0_1_2),
    .O_6_0_0_0(n78_O_6_0_0_0),
    .O_6_0_0_1(n78_O_6_0_0_1),
    .O_6_0_0_2(n78_O_6_0_0_2),
    .O_6_0_1_0(n78_O_6_0_1_0),
    .O_6_0_1_1(n78_O_6_0_1_1),
    .O_6_0_1_2(n78_O_6_0_1_2),
    .O_7_0_0_0(n78_O_7_0_0_0),
    .O_7_0_0_1(n78_O_7_0_0_1),
    .O_7_0_0_2(n78_O_7_0_0_2),
    .O_7_0_1_0(n78_O_7_0_1_0),
    .O_7_0_1_1(n78_O_7_0_1_1),
    .O_7_0_1_2(n78_O_7_0_1_2),
    .O_8_0_0_0(n78_O_8_0_0_0),
    .O_8_0_0_1(n78_O_8_0_0_1),
    .O_8_0_0_2(n78_O_8_0_0_2),
    .O_8_0_1_0(n78_O_8_0_1_0),
    .O_8_0_1_1(n78_O_8_0_1_1),
    .O_8_0_1_2(n78_O_8_0_1_2),
    .O_9_0_0_0(n78_O_9_0_0_0),
    .O_9_0_0_1(n78_O_9_0_0_1),
    .O_9_0_0_2(n78_O_9_0_0_2),
    .O_9_0_1_0(n78_O_9_0_1_0),
    .O_9_0_1_1(n78_O_9_0_1_1),
    .O_9_0_1_2(n78_O_9_0_1_2),
    .O_10_0_0_0(n78_O_10_0_0_0),
    .O_10_0_0_1(n78_O_10_0_0_1),
    .O_10_0_0_2(n78_O_10_0_0_2),
    .O_10_0_1_0(n78_O_10_0_1_0),
    .O_10_0_1_1(n78_O_10_0_1_1),
    .O_10_0_1_2(n78_O_10_0_1_2),
    .O_11_0_0_0(n78_O_11_0_0_0),
    .O_11_0_0_1(n78_O_11_0_0_1),
    .O_11_0_0_2(n78_O_11_0_0_2),
    .O_11_0_1_0(n78_O_11_0_1_0),
    .O_11_0_1_1(n78_O_11_0_1_1),
    .O_11_0_1_2(n78_O_11_0_1_2),
    .O_12_0_0_0(n78_O_12_0_0_0),
    .O_12_0_0_1(n78_O_12_0_0_1),
    .O_12_0_0_2(n78_O_12_0_0_2),
    .O_12_0_1_0(n78_O_12_0_1_0),
    .O_12_0_1_1(n78_O_12_0_1_1),
    .O_12_0_1_2(n78_O_12_0_1_2),
    .O_13_0_0_0(n78_O_13_0_0_0),
    .O_13_0_0_1(n78_O_13_0_0_1),
    .O_13_0_0_2(n78_O_13_0_0_2),
    .O_13_0_1_0(n78_O_13_0_1_0),
    .O_13_0_1_1(n78_O_13_0_1_1),
    .O_13_0_1_2(n78_O_13_0_1_2),
    .O_14_0_0_0(n78_O_14_0_0_0),
    .O_14_0_0_1(n78_O_14_0_0_1),
    .O_14_0_0_2(n78_O_14_0_0_2),
    .O_14_0_1_0(n78_O_14_0_1_0),
    .O_14_0_1_1(n78_O_14_0_1_1),
    .O_14_0_1_2(n78_O_14_0_1_2),
    .O_15_0_0_0(n78_O_15_0_0_0),
    .O_15_0_0_1(n78_O_15_0_0_1),
    .O_15_0_0_2(n78_O_15_0_0_2),
    .O_15_0_1_0(n78_O_15_0_1_0),
    .O_15_0_1_1(n78_O_15_0_1_1),
    .O_15_0_1_2(n78_O_15_0_1_2)
  );
  ShiftTS_2 n88 ( // @[Top.scala 150:21]
    .clock(n88_clock),
    .valid_up(n88_valid_up),
    .valid_down(n88_valid_down),
    .I_0_0_0(n88_I_0_0_0),
    .I_1_0_0(n88_I_1_0_0),
    .I_2_0_0(n88_I_2_0_0),
    .I_3_0_0(n88_I_3_0_0),
    .I_4_0_0(n88_I_4_0_0),
    .I_5_0_0(n88_I_5_0_0),
    .I_6_0_0(n88_I_6_0_0),
    .I_7_0_0(n88_I_7_0_0),
    .I_8_0_0(n88_I_8_0_0),
    .I_9_0_0(n88_I_9_0_0),
    .I_10_0_0(n88_I_10_0_0),
    .I_11_0_0(n88_I_11_0_0),
    .I_12_0_0(n88_I_12_0_0),
    .I_13_0_0(n88_I_13_0_0),
    .I_14_0_0(n88_I_14_0_0),
    .I_15_0_0(n88_I_15_0_0),
    .O_0_0_0(n88_O_0_0_0),
    .O_1_0_0(n88_O_1_0_0),
    .O_2_0_0(n88_O_2_0_0),
    .O_3_0_0(n88_O_3_0_0),
    .O_4_0_0(n88_O_4_0_0),
    .O_5_0_0(n88_O_5_0_0),
    .O_6_0_0(n88_O_6_0_0),
    .O_7_0_0(n88_O_7_0_0),
    .O_8_0_0(n88_O_8_0_0),
    .O_9_0_0(n88_O_9_0_0),
    .O_10_0_0(n88_O_10_0_0),
    .O_11_0_0(n88_O_11_0_0),
    .O_12_0_0(n88_O_12_0_0),
    .O_13_0_0(n88_O_13_0_0),
    .O_14_0_0(n88_O_14_0_0),
    .O_15_0_0(n88_O_15_0_0)
  );
  ShiftTS_2 n89 ( // @[Top.scala 153:21]
    .clock(n89_clock),
    .valid_up(n89_valid_up),
    .valid_down(n89_valid_down),
    .I_0_0_0(n89_I_0_0_0),
    .I_1_0_0(n89_I_1_0_0),
    .I_2_0_0(n89_I_2_0_0),
    .I_3_0_0(n89_I_3_0_0),
    .I_4_0_0(n89_I_4_0_0),
    .I_5_0_0(n89_I_5_0_0),
    .I_6_0_0(n89_I_6_0_0),
    .I_7_0_0(n89_I_7_0_0),
    .I_8_0_0(n89_I_8_0_0),
    .I_9_0_0(n89_I_9_0_0),
    .I_10_0_0(n89_I_10_0_0),
    .I_11_0_0(n89_I_11_0_0),
    .I_12_0_0(n89_I_12_0_0),
    .I_13_0_0(n89_I_13_0_0),
    .I_14_0_0(n89_I_14_0_0),
    .I_15_0_0(n89_I_15_0_0),
    .O_0_0_0(n89_O_0_0_0),
    .O_1_0_0(n89_O_1_0_0),
    .O_2_0_0(n89_O_2_0_0),
    .O_3_0_0(n89_O_3_0_0),
    .O_4_0_0(n89_O_4_0_0),
    .O_5_0_0(n89_O_5_0_0),
    .O_6_0_0(n89_O_6_0_0),
    .O_7_0_0(n89_O_7_0_0),
    .O_8_0_0(n89_O_8_0_0),
    .O_9_0_0(n89_O_9_0_0),
    .O_10_0_0(n89_O_10_0_0),
    .O_11_0_0(n89_O_11_0_0),
    .O_12_0_0(n89_O_12_0_0),
    .O_13_0_0(n89_O_13_0_0),
    .O_14_0_0(n89_O_14_0_0),
    .O_15_0_0(n89_O_15_0_0)
  );
  Map2T n90 ( // @[Top.scala 156:21]
    .valid_up(n90_valid_up),
    .valid_down(n90_valid_down),
    .I0_0_0_0(n90_I0_0_0_0),
    .I0_1_0_0(n90_I0_1_0_0),
    .I0_2_0_0(n90_I0_2_0_0),
    .I0_3_0_0(n90_I0_3_0_0),
    .I0_4_0_0(n90_I0_4_0_0),
    .I0_5_0_0(n90_I0_5_0_0),
    .I0_6_0_0(n90_I0_6_0_0),
    .I0_7_0_0(n90_I0_7_0_0),
    .I0_8_0_0(n90_I0_8_0_0),
    .I0_9_0_0(n90_I0_9_0_0),
    .I0_10_0_0(n90_I0_10_0_0),
    .I0_11_0_0(n90_I0_11_0_0),
    .I0_12_0_0(n90_I0_12_0_0),
    .I0_13_0_0(n90_I0_13_0_0),
    .I0_14_0_0(n90_I0_14_0_0),
    .I0_15_0_0(n90_I0_15_0_0),
    .I1_0_0_0(n90_I1_0_0_0),
    .I1_1_0_0(n90_I1_1_0_0),
    .I1_2_0_0(n90_I1_2_0_0),
    .I1_3_0_0(n90_I1_3_0_0),
    .I1_4_0_0(n90_I1_4_0_0),
    .I1_5_0_0(n90_I1_5_0_0),
    .I1_6_0_0(n90_I1_6_0_0),
    .I1_7_0_0(n90_I1_7_0_0),
    .I1_8_0_0(n90_I1_8_0_0),
    .I1_9_0_0(n90_I1_9_0_0),
    .I1_10_0_0(n90_I1_10_0_0),
    .I1_11_0_0(n90_I1_11_0_0),
    .I1_12_0_0(n90_I1_12_0_0),
    .I1_13_0_0(n90_I1_13_0_0),
    .I1_14_0_0(n90_I1_14_0_0),
    .I1_15_0_0(n90_I1_15_0_0),
    .O_0_0_0_0(n90_O_0_0_0_0),
    .O_0_0_0_1(n90_O_0_0_0_1),
    .O_1_0_0_0(n90_O_1_0_0_0),
    .O_1_0_0_1(n90_O_1_0_0_1),
    .O_2_0_0_0(n90_O_2_0_0_0),
    .O_2_0_0_1(n90_O_2_0_0_1),
    .O_3_0_0_0(n90_O_3_0_0_0),
    .O_3_0_0_1(n90_O_3_0_0_1),
    .O_4_0_0_0(n90_O_4_0_0_0),
    .O_4_0_0_1(n90_O_4_0_0_1),
    .O_5_0_0_0(n90_O_5_0_0_0),
    .O_5_0_0_1(n90_O_5_0_0_1),
    .O_6_0_0_0(n90_O_6_0_0_0),
    .O_6_0_0_1(n90_O_6_0_0_1),
    .O_7_0_0_0(n90_O_7_0_0_0),
    .O_7_0_0_1(n90_O_7_0_0_1),
    .O_8_0_0_0(n90_O_8_0_0_0),
    .O_8_0_0_1(n90_O_8_0_0_1),
    .O_9_0_0_0(n90_O_9_0_0_0),
    .O_9_0_0_1(n90_O_9_0_0_1),
    .O_10_0_0_0(n90_O_10_0_0_0),
    .O_10_0_0_1(n90_O_10_0_0_1),
    .O_11_0_0_0(n90_O_11_0_0_0),
    .O_11_0_0_1(n90_O_11_0_0_1),
    .O_12_0_0_0(n90_O_12_0_0_0),
    .O_12_0_0_1(n90_O_12_0_0_1),
    .O_13_0_0_0(n90_O_13_0_0_0),
    .O_13_0_0_1(n90_O_13_0_0_1),
    .O_14_0_0_0(n90_O_14_0_0_0),
    .O_14_0_0_1(n90_O_14_0_0_1),
    .O_15_0_0_0(n90_O_15_0_0_0),
    .O_15_0_0_1(n90_O_15_0_0_1)
  );
  Map2T_1 n103 ( // @[Top.scala 160:22]
    .valid_up(n103_valid_up),
    .valid_down(n103_valid_down),
    .I0_0_0_0_0(n103_I0_0_0_0_0),
    .I0_0_0_0_1(n103_I0_0_0_0_1),
    .I0_1_0_0_0(n103_I0_1_0_0_0),
    .I0_1_0_0_1(n103_I0_1_0_0_1),
    .I0_2_0_0_0(n103_I0_2_0_0_0),
    .I0_2_0_0_1(n103_I0_2_0_0_1),
    .I0_3_0_0_0(n103_I0_3_0_0_0),
    .I0_3_0_0_1(n103_I0_3_0_0_1),
    .I0_4_0_0_0(n103_I0_4_0_0_0),
    .I0_4_0_0_1(n103_I0_4_0_0_1),
    .I0_5_0_0_0(n103_I0_5_0_0_0),
    .I0_5_0_0_1(n103_I0_5_0_0_1),
    .I0_6_0_0_0(n103_I0_6_0_0_0),
    .I0_6_0_0_1(n103_I0_6_0_0_1),
    .I0_7_0_0_0(n103_I0_7_0_0_0),
    .I0_7_0_0_1(n103_I0_7_0_0_1),
    .I0_8_0_0_0(n103_I0_8_0_0_0),
    .I0_8_0_0_1(n103_I0_8_0_0_1),
    .I0_9_0_0_0(n103_I0_9_0_0_0),
    .I0_9_0_0_1(n103_I0_9_0_0_1),
    .I0_10_0_0_0(n103_I0_10_0_0_0),
    .I0_10_0_0_1(n103_I0_10_0_0_1),
    .I0_11_0_0_0(n103_I0_11_0_0_0),
    .I0_11_0_0_1(n103_I0_11_0_0_1),
    .I0_12_0_0_0(n103_I0_12_0_0_0),
    .I0_12_0_0_1(n103_I0_12_0_0_1),
    .I0_13_0_0_0(n103_I0_13_0_0_0),
    .I0_13_0_0_1(n103_I0_13_0_0_1),
    .I0_14_0_0_0(n103_I0_14_0_0_0),
    .I0_14_0_0_1(n103_I0_14_0_0_1),
    .I0_15_0_0_0(n103_I0_15_0_0_0),
    .I0_15_0_0_1(n103_I0_15_0_0_1),
    .I1_0_0_0(n103_I1_0_0_0),
    .I1_1_0_0(n103_I1_1_0_0),
    .I1_2_0_0(n103_I1_2_0_0),
    .I1_3_0_0(n103_I1_3_0_0),
    .I1_4_0_0(n103_I1_4_0_0),
    .I1_5_0_0(n103_I1_5_0_0),
    .I1_6_0_0(n103_I1_6_0_0),
    .I1_7_0_0(n103_I1_7_0_0),
    .I1_8_0_0(n103_I1_8_0_0),
    .I1_9_0_0(n103_I1_9_0_0),
    .I1_10_0_0(n103_I1_10_0_0),
    .I1_11_0_0(n103_I1_11_0_0),
    .I1_12_0_0(n103_I1_12_0_0),
    .I1_13_0_0(n103_I1_13_0_0),
    .I1_14_0_0(n103_I1_14_0_0),
    .I1_15_0_0(n103_I1_15_0_0),
    .O_0_0_0_0(n103_O_0_0_0_0),
    .O_0_0_0_1(n103_O_0_0_0_1),
    .O_0_0_0_2(n103_O_0_0_0_2),
    .O_1_0_0_0(n103_O_1_0_0_0),
    .O_1_0_0_1(n103_O_1_0_0_1),
    .O_1_0_0_2(n103_O_1_0_0_2),
    .O_2_0_0_0(n103_O_2_0_0_0),
    .O_2_0_0_1(n103_O_2_0_0_1),
    .O_2_0_0_2(n103_O_2_0_0_2),
    .O_3_0_0_0(n103_O_3_0_0_0),
    .O_3_0_0_1(n103_O_3_0_0_1),
    .O_3_0_0_2(n103_O_3_0_0_2),
    .O_4_0_0_0(n103_O_4_0_0_0),
    .O_4_0_0_1(n103_O_4_0_0_1),
    .O_4_0_0_2(n103_O_4_0_0_2),
    .O_5_0_0_0(n103_O_5_0_0_0),
    .O_5_0_0_1(n103_O_5_0_0_1),
    .O_5_0_0_2(n103_O_5_0_0_2),
    .O_6_0_0_0(n103_O_6_0_0_0),
    .O_6_0_0_1(n103_O_6_0_0_1),
    .O_6_0_0_2(n103_O_6_0_0_2),
    .O_7_0_0_0(n103_O_7_0_0_0),
    .O_7_0_0_1(n103_O_7_0_0_1),
    .O_7_0_0_2(n103_O_7_0_0_2),
    .O_8_0_0_0(n103_O_8_0_0_0),
    .O_8_0_0_1(n103_O_8_0_0_1),
    .O_8_0_0_2(n103_O_8_0_0_2),
    .O_9_0_0_0(n103_O_9_0_0_0),
    .O_9_0_0_1(n103_O_9_0_0_1),
    .O_9_0_0_2(n103_O_9_0_0_2),
    .O_10_0_0_0(n103_O_10_0_0_0),
    .O_10_0_0_1(n103_O_10_0_0_1),
    .O_10_0_0_2(n103_O_10_0_0_2),
    .O_11_0_0_0(n103_O_11_0_0_0),
    .O_11_0_0_1(n103_O_11_0_0_1),
    .O_11_0_0_2(n103_O_11_0_0_2),
    .O_12_0_0_0(n103_O_12_0_0_0),
    .O_12_0_0_1(n103_O_12_0_0_1),
    .O_12_0_0_2(n103_O_12_0_0_2),
    .O_13_0_0_0(n103_O_13_0_0_0),
    .O_13_0_0_1(n103_O_13_0_0_1),
    .O_13_0_0_2(n103_O_13_0_0_2),
    .O_14_0_0_0(n103_O_14_0_0_0),
    .O_14_0_0_1(n103_O_14_0_0_1),
    .O_14_0_0_2(n103_O_14_0_0_2),
    .O_15_0_0_0(n103_O_15_0_0_0),
    .O_15_0_0_1(n103_O_15_0_0_1),
    .O_15_0_0_2(n103_O_15_0_0_2)
  );
  MapT n124 ( // @[Top.scala 164:22]
    .valid_up(n124_valid_up),
    .valid_down(n124_valid_down),
    .I_0_0_0_0(n124_I_0_0_0_0),
    .I_0_0_0_1(n124_I_0_0_0_1),
    .I_0_0_0_2(n124_I_0_0_0_2),
    .I_1_0_0_0(n124_I_1_0_0_0),
    .I_1_0_0_1(n124_I_1_0_0_1),
    .I_1_0_0_2(n124_I_1_0_0_2),
    .I_2_0_0_0(n124_I_2_0_0_0),
    .I_2_0_0_1(n124_I_2_0_0_1),
    .I_2_0_0_2(n124_I_2_0_0_2),
    .I_3_0_0_0(n124_I_3_0_0_0),
    .I_3_0_0_1(n124_I_3_0_0_1),
    .I_3_0_0_2(n124_I_3_0_0_2),
    .I_4_0_0_0(n124_I_4_0_0_0),
    .I_4_0_0_1(n124_I_4_0_0_1),
    .I_4_0_0_2(n124_I_4_0_0_2),
    .I_5_0_0_0(n124_I_5_0_0_0),
    .I_5_0_0_1(n124_I_5_0_0_1),
    .I_5_0_0_2(n124_I_5_0_0_2),
    .I_6_0_0_0(n124_I_6_0_0_0),
    .I_6_0_0_1(n124_I_6_0_0_1),
    .I_6_0_0_2(n124_I_6_0_0_2),
    .I_7_0_0_0(n124_I_7_0_0_0),
    .I_7_0_0_1(n124_I_7_0_0_1),
    .I_7_0_0_2(n124_I_7_0_0_2),
    .I_8_0_0_0(n124_I_8_0_0_0),
    .I_8_0_0_1(n124_I_8_0_0_1),
    .I_8_0_0_2(n124_I_8_0_0_2),
    .I_9_0_0_0(n124_I_9_0_0_0),
    .I_9_0_0_1(n124_I_9_0_0_1),
    .I_9_0_0_2(n124_I_9_0_0_2),
    .I_10_0_0_0(n124_I_10_0_0_0),
    .I_10_0_0_1(n124_I_10_0_0_1),
    .I_10_0_0_2(n124_I_10_0_0_2),
    .I_11_0_0_0(n124_I_11_0_0_0),
    .I_11_0_0_1(n124_I_11_0_0_1),
    .I_11_0_0_2(n124_I_11_0_0_2),
    .I_12_0_0_0(n124_I_12_0_0_0),
    .I_12_0_0_1(n124_I_12_0_0_1),
    .I_12_0_0_2(n124_I_12_0_0_2),
    .I_13_0_0_0(n124_I_13_0_0_0),
    .I_13_0_0_1(n124_I_13_0_0_1),
    .I_13_0_0_2(n124_I_13_0_0_2),
    .I_14_0_0_0(n124_I_14_0_0_0),
    .I_14_0_0_1(n124_I_14_0_0_1),
    .I_14_0_0_2(n124_I_14_0_0_2),
    .I_15_0_0_0(n124_I_15_0_0_0),
    .I_15_0_0_1(n124_I_15_0_0_1),
    .I_15_0_0_2(n124_I_15_0_0_2),
    .O_0_0_0(n124_O_0_0_0),
    .O_0_0_1(n124_O_0_0_1),
    .O_0_0_2(n124_O_0_0_2),
    .O_1_0_0(n124_O_1_0_0),
    .O_1_0_1(n124_O_1_0_1),
    .O_1_0_2(n124_O_1_0_2),
    .O_2_0_0(n124_O_2_0_0),
    .O_2_0_1(n124_O_2_0_1),
    .O_2_0_2(n124_O_2_0_2),
    .O_3_0_0(n124_O_3_0_0),
    .O_3_0_1(n124_O_3_0_1),
    .O_3_0_2(n124_O_3_0_2),
    .O_4_0_0(n124_O_4_0_0),
    .O_4_0_1(n124_O_4_0_1),
    .O_4_0_2(n124_O_4_0_2),
    .O_5_0_0(n124_O_5_0_0),
    .O_5_0_1(n124_O_5_0_1),
    .O_5_0_2(n124_O_5_0_2),
    .O_6_0_0(n124_O_6_0_0),
    .O_6_0_1(n124_O_6_0_1),
    .O_6_0_2(n124_O_6_0_2),
    .O_7_0_0(n124_O_7_0_0),
    .O_7_0_1(n124_O_7_0_1),
    .O_7_0_2(n124_O_7_0_2),
    .O_8_0_0(n124_O_8_0_0),
    .O_8_0_1(n124_O_8_0_1),
    .O_8_0_2(n124_O_8_0_2),
    .O_9_0_0(n124_O_9_0_0),
    .O_9_0_1(n124_O_9_0_1),
    .O_9_0_2(n124_O_9_0_2),
    .O_10_0_0(n124_O_10_0_0),
    .O_10_0_1(n124_O_10_0_1),
    .O_10_0_2(n124_O_10_0_2),
    .O_11_0_0(n124_O_11_0_0),
    .O_11_0_1(n124_O_11_0_1),
    .O_11_0_2(n124_O_11_0_2),
    .O_12_0_0(n124_O_12_0_0),
    .O_12_0_1(n124_O_12_0_1),
    .O_12_0_2(n124_O_12_0_2),
    .O_13_0_0(n124_O_13_0_0),
    .O_13_0_1(n124_O_13_0_1),
    .O_13_0_2(n124_O_13_0_2),
    .O_14_0_0(n124_O_14_0_0),
    .O_14_0_1(n124_O_14_0_1),
    .O_14_0_2(n124_O_14_0_2),
    .O_15_0_0(n124_O_15_0_0),
    .O_15_0_1(n124_O_15_0_1),
    .O_15_0_2(n124_O_15_0_2)
  );
  Map2T_7 n125 ( // @[Top.scala 167:22]
    .valid_up(n125_valid_up),
    .valid_down(n125_valid_down),
    .I0_0_0_0_0(n125_I0_0_0_0_0),
    .I0_0_0_0_1(n125_I0_0_0_0_1),
    .I0_0_0_0_2(n125_I0_0_0_0_2),
    .I0_0_0_1_0(n125_I0_0_0_1_0),
    .I0_0_0_1_1(n125_I0_0_0_1_1),
    .I0_0_0_1_2(n125_I0_0_0_1_2),
    .I0_1_0_0_0(n125_I0_1_0_0_0),
    .I0_1_0_0_1(n125_I0_1_0_0_1),
    .I0_1_0_0_2(n125_I0_1_0_0_2),
    .I0_1_0_1_0(n125_I0_1_0_1_0),
    .I0_1_0_1_1(n125_I0_1_0_1_1),
    .I0_1_0_1_2(n125_I0_1_0_1_2),
    .I0_2_0_0_0(n125_I0_2_0_0_0),
    .I0_2_0_0_1(n125_I0_2_0_0_1),
    .I0_2_0_0_2(n125_I0_2_0_0_2),
    .I0_2_0_1_0(n125_I0_2_0_1_0),
    .I0_2_0_1_1(n125_I0_2_0_1_1),
    .I0_2_0_1_2(n125_I0_2_0_1_2),
    .I0_3_0_0_0(n125_I0_3_0_0_0),
    .I0_3_0_0_1(n125_I0_3_0_0_1),
    .I0_3_0_0_2(n125_I0_3_0_0_2),
    .I0_3_0_1_0(n125_I0_3_0_1_0),
    .I0_3_0_1_1(n125_I0_3_0_1_1),
    .I0_3_0_1_2(n125_I0_3_0_1_2),
    .I0_4_0_0_0(n125_I0_4_0_0_0),
    .I0_4_0_0_1(n125_I0_4_0_0_1),
    .I0_4_0_0_2(n125_I0_4_0_0_2),
    .I0_4_0_1_0(n125_I0_4_0_1_0),
    .I0_4_0_1_1(n125_I0_4_0_1_1),
    .I0_4_0_1_2(n125_I0_4_0_1_2),
    .I0_5_0_0_0(n125_I0_5_0_0_0),
    .I0_5_0_0_1(n125_I0_5_0_0_1),
    .I0_5_0_0_2(n125_I0_5_0_0_2),
    .I0_5_0_1_0(n125_I0_5_0_1_0),
    .I0_5_0_1_1(n125_I0_5_0_1_1),
    .I0_5_0_1_2(n125_I0_5_0_1_2),
    .I0_6_0_0_0(n125_I0_6_0_0_0),
    .I0_6_0_0_1(n125_I0_6_0_0_1),
    .I0_6_0_0_2(n125_I0_6_0_0_2),
    .I0_6_0_1_0(n125_I0_6_0_1_0),
    .I0_6_0_1_1(n125_I0_6_0_1_1),
    .I0_6_0_1_2(n125_I0_6_0_1_2),
    .I0_7_0_0_0(n125_I0_7_0_0_0),
    .I0_7_0_0_1(n125_I0_7_0_0_1),
    .I0_7_0_0_2(n125_I0_7_0_0_2),
    .I0_7_0_1_0(n125_I0_7_0_1_0),
    .I0_7_0_1_1(n125_I0_7_0_1_1),
    .I0_7_0_1_2(n125_I0_7_0_1_2),
    .I0_8_0_0_0(n125_I0_8_0_0_0),
    .I0_8_0_0_1(n125_I0_8_0_0_1),
    .I0_8_0_0_2(n125_I0_8_0_0_2),
    .I0_8_0_1_0(n125_I0_8_0_1_0),
    .I0_8_0_1_1(n125_I0_8_0_1_1),
    .I0_8_0_1_2(n125_I0_8_0_1_2),
    .I0_9_0_0_0(n125_I0_9_0_0_0),
    .I0_9_0_0_1(n125_I0_9_0_0_1),
    .I0_9_0_0_2(n125_I0_9_0_0_2),
    .I0_9_0_1_0(n125_I0_9_0_1_0),
    .I0_9_0_1_1(n125_I0_9_0_1_1),
    .I0_9_0_1_2(n125_I0_9_0_1_2),
    .I0_10_0_0_0(n125_I0_10_0_0_0),
    .I0_10_0_0_1(n125_I0_10_0_0_1),
    .I0_10_0_0_2(n125_I0_10_0_0_2),
    .I0_10_0_1_0(n125_I0_10_0_1_0),
    .I0_10_0_1_1(n125_I0_10_0_1_1),
    .I0_10_0_1_2(n125_I0_10_0_1_2),
    .I0_11_0_0_0(n125_I0_11_0_0_0),
    .I0_11_0_0_1(n125_I0_11_0_0_1),
    .I0_11_0_0_2(n125_I0_11_0_0_2),
    .I0_11_0_1_0(n125_I0_11_0_1_0),
    .I0_11_0_1_1(n125_I0_11_0_1_1),
    .I0_11_0_1_2(n125_I0_11_0_1_2),
    .I0_12_0_0_0(n125_I0_12_0_0_0),
    .I0_12_0_0_1(n125_I0_12_0_0_1),
    .I0_12_0_0_2(n125_I0_12_0_0_2),
    .I0_12_0_1_0(n125_I0_12_0_1_0),
    .I0_12_0_1_1(n125_I0_12_0_1_1),
    .I0_12_0_1_2(n125_I0_12_0_1_2),
    .I0_13_0_0_0(n125_I0_13_0_0_0),
    .I0_13_0_0_1(n125_I0_13_0_0_1),
    .I0_13_0_0_2(n125_I0_13_0_0_2),
    .I0_13_0_1_0(n125_I0_13_0_1_0),
    .I0_13_0_1_1(n125_I0_13_0_1_1),
    .I0_13_0_1_2(n125_I0_13_0_1_2),
    .I0_14_0_0_0(n125_I0_14_0_0_0),
    .I0_14_0_0_1(n125_I0_14_0_0_1),
    .I0_14_0_0_2(n125_I0_14_0_0_2),
    .I0_14_0_1_0(n125_I0_14_0_1_0),
    .I0_14_0_1_1(n125_I0_14_0_1_1),
    .I0_14_0_1_2(n125_I0_14_0_1_2),
    .I0_15_0_0_0(n125_I0_15_0_0_0),
    .I0_15_0_0_1(n125_I0_15_0_0_1),
    .I0_15_0_0_2(n125_I0_15_0_0_2),
    .I0_15_0_1_0(n125_I0_15_0_1_0),
    .I0_15_0_1_1(n125_I0_15_0_1_1),
    .I0_15_0_1_2(n125_I0_15_0_1_2),
    .I1_0_0_0(n125_I1_0_0_0),
    .I1_0_0_1(n125_I1_0_0_1),
    .I1_0_0_2(n125_I1_0_0_2),
    .I1_1_0_0(n125_I1_1_0_0),
    .I1_1_0_1(n125_I1_1_0_1),
    .I1_1_0_2(n125_I1_1_0_2),
    .I1_2_0_0(n125_I1_2_0_0),
    .I1_2_0_1(n125_I1_2_0_1),
    .I1_2_0_2(n125_I1_2_0_2),
    .I1_3_0_0(n125_I1_3_0_0),
    .I1_3_0_1(n125_I1_3_0_1),
    .I1_3_0_2(n125_I1_3_0_2),
    .I1_4_0_0(n125_I1_4_0_0),
    .I1_4_0_1(n125_I1_4_0_1),
    .I1_4_0_2(n125_I1_4_0_2),
    .I1_5_0_0(n125_I1_5_0_0),
    .I1_5_0_1(n125_I1_5_0_1),
    .I1_5_0_2(n125_I1_5_0_2),
    .I1_6_0_0(n125_I1_6_0_0),
    .I1_6_0_1(n125_I1_6_0_1),
    .I1_6_0_2(n125_I1_6_0_2),
    .I1_7_0_0(n125_I1_7_0_0),
    .I1_7_0_1(n125_I1_7_0_1),
    .I1_7_0_2(n125_I1_7_0_2),
    .I1_8_0_0(n125_I1_8_0_0),
    .I1_8_0_1(n125_I1_8_0_1),
    .I1_8_0_2(n125_I1_8_0_2),
    .I1_9_0_0(n125_I1_9_0_0),
    .I1_9_0_1(n125_I1_9_0_1),
    .I1_9_0_2(n125_I1_9_0_2),
    .I1_10_0_0(n125_I1_10_0_0),
    .I1_10_0_1(n125_I1_10_0_1),
    .I1_10_0_2(n125_I1_10_0_2),
    .I1_11_0_0(n125_I1_11_0_0),
    .I1_11_0_1(n125_I1_11_0_1),
    .I1_11_0_2(n125_I1_11_0_2),
    .I1_12_0_0(n125_I1_12_0_0),
    .I1_12_0_1(n125_I1_12_0_1),
    .I1_12_0_2(n125_I1_12_0_2),
    .I1_13_0_0(n125_I1_13_0_0),
    .I1_13_0_1(n125_I1_13_0_1),
    .I1_13_0_2(n125_I1_13_0_2),
    .I1_14_0_0(n125_I1_14_0_0),
    .I1_14_0_1(n125_I1_14_0_1),
    .I1_14_0_2(n125_I1_14_0_2),
    .I1_15_0_0(n125_I1_15_0_0),
    .I1_15_0_1(n125_I1_15_0_1),
    .I1_15_0_2(n125_I1_15_0_2),
    .O_0_0_0_0(n125_O_0_0_0_0),
    .O_0_0_0_1(n125_O_0_0_0_1),
    .O_0_0_0_2(n125_O_0_0_0_2),
    .O_0_0_1_0(n125_O_0_0_1_0),
    .O_0_0_1_1(n125_O_0_0_1_1),
    .O_0_0_1_2(n125_O_0_0_1_2),
    .O_0_0_2_0(n125_O_0_0_2_0),
    .O_0_0_2_1(n125_O_0_0_2_1),
    .O_0_0_2_2(n125_O_0_0_2_2),
    .O_1_0_0_0(n125_O_1_0_0_0),
    .O_1_0_0_1(n125_O_1_0_0_1),
    .O_1_0_0_2(n125_O_1_0_0_2),
    .O_1_0_1_0(n125_O_1_0_1_0),
    .O_1_0_1_1(n125_O_1_0_1_1),
    .O_1_0_1_2(n125_O_1_0_1_2),
    .O_1_0_2_0(n125_O_1_0_2_0),
    .O_1_0_2_1(n125_O_1_0_2_1),
    .O_1_0_2_2(n125_O_1_0_2_2),
    .O_2_0_0_0(n125_O_2_0_0_0),
    .O_2_0_0_1(n125_O_2_0_0_1),
    .O_2_0_0_2(n125_O_2_0_0_2),
    .O_2_0_1_0(n125_O_2_0_1_0),
    .O_2_0_1_1(n125_O_2_0_1_1),
    .O_2_0_1_2(n125_O_2_0_1_2),
    .O_2_0_2_0(n125_O_2_0_2_0),
    .O_2_0_2_1(n125_O_2_0_2_1),
    .O_2_0_2_2(n125_O_2_0_2_2),
    .O_3_0_0_0(n125_O_3_0_0_0),
    .O_3_0_0_1(n125_O_3_0_0_1),
    .O_3_0_0_2(n125_O_3_0_0_2),
    .O_3_0_1_0(n125_O_3_0_1_0),
    .O_3_0_1_1(n125_O_3_0_1_1),
    .O_3_0_1_2(n125_O_3_0_1_2),
    .O_3_0_2_0(n125_O_3_0_2_0),
    .O_3_0_2_1(n125_O_3_0_2_1),
    .O_3_0_2_2(n125_O_3_0_2_2),
    .O_4_0_0_0(n125_O_4_0_0_0),
    .O_4_0_0_1(n125_O_4_0_0_1),
    .O_4_0_0_2(n125_O_4_0_0_2),
    .O_4_0_1_0(n125_O_4_0_1_0),
    .O_4_0_1_1(n125_O_4_0_1_1),
    .O_4_0_1_2(n125_O_4_0_1_2),
    .O_4_0_2_0(n125_O_4_0_2_0),
    .O_4_0_2_1(n125_O_4_0_2_1),
    .O_4_0_2_2(n125_O_4_0_2_2),
    .O_5_0_0_0(n125_O_5_0_0_0),
    .O_5_0_0_1(n125_O_5_0_0_1),
    .O_5_0_0_2(n125_O_5_0_0_2),
    .O_5_0_1_0(n125_O_5_0_1_0),
    .O_5_0_1_1(n125_O_5_0_1_1),
    .O_5_0_1_2(n125_O_5_0_1_2),
    .O_5_0_2_0(n125_O_5_0_2_0),
    .O_5_0_2_1(n125_O_5_0_2_1),
    .O_5_0_2_2(n125_O_5_0_2_2),
    .O_6_0_0_0(n125_O_6_0_0_0),
    .O_6_0_0_1(n125_O_6_0_0_1),
    .O_6_0_0_2(n125_O_6_0_0_2),
    .O_6_0_1_0(n125_O_6_0_1_0),
    .O_6_0_1_1(n125_O_6_0_1_1),
    .O_6_0_1_2(n125_O_6_0_1_2),
    .O_6_0_2_0(n125_O_6_0_2_0),
    .O_6_0_2_1(n125_O_6_0_2_1),
    .O_6_0_2_2(n125_O_6_0_2_2),
    .O_7_0_0_0(n125_O_7_0_0_0),
    .O_7_0_0_1(n125_O_7_0_0_1),
    .O_7_0_0_2(n125_O_7_0_0_2),
    .O_7_0_1_0(n125_O_7_0_1_0),
    .O_7_0_1_1(n125_O_7_0_1_1),
    .O_7_0_1_2(n125_O_7_0_1_2),
    .O_7_0_2_0(n125_O_7_0_2_0),
    .O_7_0_2_1(n125_O_7_0_2_1),
    .O_7_0_2_2(n125_O_7_0_2_2),
    .O_8_0_0_0(n125_O_8_0_0_0),
    .O_8_0_0_1(n125_O_8_0_0_1),
    .O_8_0_0_2(n125_O_8_0_0_2),
    .O_8_0_1_0(n125_O_8_0_1_0),
    .O_8_0_1_1(n125_O_8_0_1_1),
    .O_8_0_1_2(n125_O_8_0_1_2),
    .O_8_0_2_0(n125_O_8_0_2_0),
    .O_8_0_2_1(n125_O_8_0_2_1),
    .O_8_0_2_2(n125_O_8_0_2_2),
    .O_9_0_0_0(n125_O_9_0_0_0),
    .O_9_0_0_1(n125_O_9_0_0_1),
    .O_9_0_0_2(n125_O_9_0_0_2),
    .O_9_0_1_0(n125_O_9_0_1_0),
    .O_9_0_1_1(n125_O_9_0_1_1),
    .O_9_0_1_2(n125_O_9_0_1_2),
    .O_9_0_2_0(n125_O_9_0_2_0),
    .O_9_0_2_1(n125_O_9_0_2_1),
    .O_9_0_2_2(n125_O_9_0_2_2),
    .O_10_0_0_0(n125_O_10_0_0_0),
    .O_10_0_0_1(n125_O_10_0_0_1),
    .O_10_0_0_2(n125_O_10_0_0_2),
    .O_10_0_1_0(n125_O_10_0_1_0),
    .O_10_0_1_1(n125_O_10_0_1_1),
    .O_10_0_1_2(n125_O_10_0_1_2),
    .O_10_0_2_0(n125_O_10_0_2_0),
    .O_10_0_2_1(n125_O_10_0_2_1),
    .O_10_0_2_2(n125_O_10_0_2_2),
    .O_11_0_0_0(n125_O_11_0_0_0),
    .O_11_0_0_1(n125_O_11_0_0_1),
    .O_11_0_0_2(n125_O_11_0_0_2),
    .O_11_0_1_0(n125_O_11_0_1_0),
    .O_11_0_1_1(n125_O_11_0_1_1),
    .O_11_0_1_2(n125_O_11_0_1_2),
    .O_11_0_2_0(n125_O_11_0_2_0),
    .O_11_0_2_1(n125_O_11_0_2_1),
    .O_11_0_2_2(n125_O_11_0_2_2),
    .O_12_0_0_0(n125_O_12_0_0_0),
    .O_12_0_0_1(n125_O_12_0_0_1),
    .O_12_0_0_2(n125_O_12_0_0_2),
    .O_12_0_1_0(n125_O_12_0_1_0),
    .O_12_0_1_1(n125_O_12_0_1_1),
    .O_12_0_1_2(n125_O_12_0_1_2),
    .O_12_0_2_0(n125_O_12_0_2_0),
    .O_12_0_2_1(n125_O_12_0_2_1),
    .O_12_0_2_2(n125_O_12_0_2_2),
    .O_13_0_0_0(n125_O_13_0_0_0),
    .O_13_0_0_1(n125_O_13_0_0_1),
    .O_13_0_0_2(n125_O_13_0_0_2),
    .O_13_0_1_0(n125_O_13_0_1_0),
    .O_13_0_1_1(n125_O_13_0_1_1),
    .O_13_0_1_2(n125_O_13_0_1_2),
    .O_13_0_2_0(n125_O_13_0_2_0),
    .O_13_0_2_1(n125_O_13_0_2_1),
    .O_13_0_2_2(n125_O_13_0_2_2),
    .O_14_0_0_0(n125_O_14_0_0_0),
    .O_14_0_0_1(n125_O_14_0_0_1),
    .O_14_0_0_2(n125_O_14_0_0_2),
    .O_14_0_1_0(n125_O_14_0_1_0),
    .O_14_0_1_1(n125_O_14_0_1_1),
    .O_14_0_1_2(n125_O_14_0_1_2),
    .O_14_0_2_0(n125_O_14_0_2_0),
    .O_14_0_2_1(n125_O_14_0_2_1),
    .O_14_0_2_2(n125_O_14_0_2_2),
    .O_15_0_0_0(n125_O_15_0_0_0),
    .O_15_0_0_1(n125_O_15_0_0_1),
    .O_15_0_0_2(n125_O_15_0_0_2),
    .O_15_0_1_0(n125_O_15_0_1_0),
    .O_15_0_1_1(n125_O_15_0_1_1),
    .O_15_0_1_2(n125_O_15_0_1_2),
    .O_15_0_2_0(n125_O_15_0_2_0),
    .O_15_0_2_1(n125_O_15_0_2_1),
    .O_15_0_2_2(n125_O_15_0_2_2)
  );
  MapT_3 n141 ( // @[Top.scala 171:22]
    .valid_up(n141_valid_up),
    .valid_down(n141_valid_down),
    .I_0_0_0_0(n141_I_0_0_0_0),
    .I_0_0_0_1(n141_I_0_0_0_1),
    .I_0_0_0_2(n141_I_0_0_0_2),
    .I_0_0_1_0(n141_I_0_0_1_0),
    .I_0_0_1_1(n141_I_0_0_1_1),
    .I_0_0_1_2(n141_I_0_0_1_2),
    .I_0_0_2_0(n141_I_0_0_2_0),
    .I_0_0_2_1(n141_I_0_0_2_1),
    .I_0_0_2_2(n141_I_0_0_2_2),
    .I_1_0_0_0(n141_I_1_0_0_0),
    .I_1_0_0_1(n141_I_1_0_0_1),
    .I_1_0_0_2(n141_I_1_0_0_2),
    .I_1_0_1_0(n141_I_1_0_1_0),
    .I_1_0_1_1(n141_I_1_0_1_1),
    .I_1_0_1_2(n141_I_1_0_1_2),
    .I_1_0_2_0(n141_I_1_0_2_0),
    .I_1_0_2_1(n141_I_1_0_2_1),
    .I_1_0_2_2(n141_I_1_0_2_2),
    .I_2_0_0_0(n141_I_2_0_0_0),
    .I_2_0_0_1(n141_I_2_0_0_1),
    .I_2_0_0_2(n141_I_2_0_0_2),
    .I_2_0_1_0(n141_I_2_0_1_0),
    .I_2_0_1_1(n141_I_2_0_1_1),
    .I_2_0_1_2(n141_I_2_0_1_2),
    .I_2_0_2_0(n141_I_2_0_2_0),
    .I_2_0_2_1(n141_I_2_0_2_1),
    .I_2_0_2_2(n141_I_2_0_2_2),
    .I_3_0_0_0(n141_I_3_0_0_0),
    .I_3_0_0_1(n141_I_3_0_0_1),
    .I_3_0_0_2(n141_I_3_0_0_2),
    .I_3_0_1_0(n141_I_3_0_1_0),
    .I_3_0_1_1(n141_I_3_0_1_1),
    .I_3_0_1_2(n141_I_3_0_1_2),
    .I_3_0_2_0(n141_I_3_0_2_0),
    .I_3_0_2_1(n141_I_3_0_2_1),
    .I_3_0_2_2(n141_I_3_0_2_2),
    .I_4_0_0_0(n141_I_4_0_0_0),
    .I_4_0_0_1(n141_I_4_0_0_1),
    .I_4_0_0_2(n141_I_4_0_0_2),
    .I_4_0_1_0(n141_I_4_0_1_0),
    .I_4_0_1_1(n141_I_4_0_1_1),
    .I_4_0_1_2(n141_I_4_0_1_2),
    .I_4_0_2_0(n141_I_4_0_2_0),
    .I_4_0_2_1(n141_I_4_0_2_1),
    .I_4_0_2_2(n141_I_4_0_2_2),
    .I_5_0_0_0(n141_I_5_0_0_0),
    .I_5_0_0_1(n141_I_5_0_0_1),
    .I_5_0_0_2(n141_I_5_0_0_2),
    .I_5_0_1_0(n141_I_5_0_1_0),
    .I_5_0_1_1(n141_I_5_0_1_1),
    .I_5_0_1_2(n141_I_5_0_1_2),
    .I_5_0_2_0(n141_I_5_0_2_0),
    .I_5_0_2_1(n141_I_5_0_2_1),
    .I_5_0_2_2(n141_I_5_0_2_2),
    .I_6_0_0_0(n141_I_6_0_0_0),
    .I_6_0_0_1(n141_I_6_0_0_1),
    .I_6_0_0_2(n141_I_6_0_0_2),
    .I_6_0_1_0(n141_I_6_0_1_0),
    .I_6_0_1_1(n141_I_6_0_1_1),
    .I_6_0_1_2(n141_I_6_0_1_2),
    .I_6_0_2_0(n141_I_6_0_2_0),
    .I_6_0_2_1(n141_I_6_0_2_1),
    .I_6_0_2_2(n141_I_6_0_2_2),
    .I_7_0_0_0(n141_I_7_0_0_0),
    .I_7_0_0_1(n141_I_7_0_0_1),
    .I_7_0_0_2(n141_I_7_0_0_2),
    .I_7_0_1_0(n141_I_7_0_1_0),
    .I_7_0_1_1(n141_I_7_0_1_1),
    .I_7_0_1_2(n141_I_7_0_1_2),
    .I_7_0_2_0(n141_I_7_0_2_0),
    .I_7_0_2_1(n141_I_7_0_2_1),
    .I_7_0_2_2(n141_I_7_0_2_2),
    .I_8_0_0_0(n141_I_8_0_0_0),
    .I_8_0_0_1(n141_I_8_0_0_1),
    .I_8_0_0_2(n141_I_8_0_0_2),
    .I_8_0_1_0(n141_I_8_0_1_0),
    .I_8_0_1_1(n141_I_8_0_1_1),
    .I_8_0_1_2(n141_I_8_0_1_2),
    .I_8_0_2_0(n141_I_8_0_2_0),
    .I_8_0_2_1(n141_I_8_0_2_1),
    .I_8_0_2_2(n141_I_8_0_2_2),
    .I_9_0_0_0(n141_I_9_0_0_0),
    .I_9_0_0_1(n141_I_9_0_0_1),
    .I_9_0_0_2(n141_I_9_0_0_2),
    .I_9_0_1_0(n141_I_9_0_1_0),
    .I_9_0_1_1(n141_I_9_0_1_1),
    .I_9_0_1_2(n141_I_9_0_1_2),
    .I_9_0_2_0(n141_I_9_0_2_0),
    .I_9_0_2_1(n141_I_9_0_2_1),
    .I_9_0_2_2(n141_I_9_0_2_2),
    .I_10_0_0_0(n141_I_10_0_0_0),
    .I_10_0_0_1(n141_I_10_0_0_1),
    .I_10_0_0_2(n141_I_10_0_0_2),
    .I_10_0_1_0(n141_I_10_0_1_0),
    .I_10_0_1_1(n141_I_10_0_1_1),
    .I_10_0_1_2(n141_I_10_0_1_2),
    .I_10_0_2_0(n141_I_10_0_2_0),
    .I_10_0_2_1(n141_I_10_0_2_1),
    .I_10_0_2_2(n141_I_10_0_2_2),
    .I_11_0_0_0(n141_I_11_0_0_0),
    .I_11_0_0_1(n141_I_11_0_0_1),
    .I_11_0_0_2(n141_I_11_0_0_2),
    .I_11_0_1_0(n141_I_11_0_1_0),
    .I_11_0_1_1(n141_I_11_0_1_1),
    .I_11_0_1_2(n141_I_11_0_1_2),
    .I_11_0_2_0(n141_I_11_0_2_0),
    .I_11_0_2_1(n141_I_11_0_2_1),
    .I_11_0_2_2(n141_I_11_0_2_2),
    .I_12_0_0_0(n141_I_12_0_0_0),
    .I_12_0_0_1(n141_I_12_0_0_1),
    .I_12_0_0_2(n141_I_12_0_0_2),
    .I_12_0_1_0(n141_I_12_0_1_0),
    .I_12_0_1_1(n141_I_12_0_1_1),
    .I_12_0_1_2(n141_I_12_0_1_2),
    .I_12_0_2_0(n141_I_12_0_2_0),
    .I_12_0_2_1(n141_I_12_0_2_1),
    .I_12_0_2_2(n141_I_12_0_2_2),
    .I_13_0_0_0(n141_I_13_0_0_0),
    .I_13_0_0_1(n141_I_13_0_0_1),
    .I_13_0_0_2(n141_I_13_0_0_2),
    .I_13_0_1_0(n141_I_13_0_1_0),
    .I_13_0_1_1(n141_I_13_0_1_1),
    .I_13_0_1_2(n141_I_13_0_1_2),
    .I_13_0_2_0(n141_I_13_0_2_0),
    .I_13_0_2_1(n141_I_13_0_2_1),
    .I_13_0_2_2(n141_I_13_0_2_2),
    .I_14_0_0_0(n141_I_14_0_0_0),
    .I_14_0_0_1(n141_I_14_0_0_1),
    .I_14_0_0_2(n141_I_14_0_0_2),
    .I_14_0_1_0(n141_I_14_0_1_0),
    .I_14_0_1_1(n141_I_14_0_1_1),
    .I_14_0_1_2(n141_I_14_0_1_2),
    .I_14_0_2_0(n141_I_14_0_2_0),
    .I_14_0_2_1(n141_I_14_0_2_1),
    .I_14_0_2_2(n141_I_14_0_2_2),
    .I_15_0_0_0(n141_I_15_0_0_0),
    .I_15_0_0_1(n141_I_15_0_0_1),
    .I_15_0_0_2(n141_I_15_0_0_2),
    .I_15_0_1_0(n141_I_15_0_1_0),
    .I_15_0_1_1(n141_I_15_0_1_1),
    .I_15_0_1_2(n141_I_15_0_1_2),
    .I_15_0_2_0(n141_I_15_0_2_0),
    .I_15_0_2_1(n141_I_15_0_2_1),
    .I_15_0_2_2(n141_I_15_0_2_2),
    .O_0_0_0(n141_O_0_0_0),
    .O_0_0_1(n141_O_0_0_1),
    .O_0_0_2(n141_O_0_0_2),
    .O_0_1_0(n141_O_0_1_0),
    .O_0_1_1(n141_O_0_1_1),
    .O_0_1_2(n141_O_0_1_2),
    .O_0_2_0(n141_O_0_2_0),
    .O_0_2_1(n141_O_0_2_1),
    .O_0_2_2(n141_O_0_2_2),
    .O_1_0_0(n141_O_1_0_0),
    .O_1_0_1(n141_O_1_0_1),
    .O_1_0_2(n141_O_1_0_2),
    .O_1_1_0(n141_O_1_1_0),
    .O_1_1_1(n141_O_1_1_1),
    .O_1_1_2(n141_O_1_1_2),
    .O_1_2_0(n141_O_1_2_0),
    .O_1_2_1(n141_O_1_2_1),
    .O_1_2_2(n141_O_1_2_2),
    .O_2_0_0(n141_O_2_0_0),
    .O_2_0_1(n141_O_2_0_1),
    .O_2_0_2(n141_O_2_0_2),
    .O_2_1_0(n141_O_2_1_0),
    .O_2_1_1(n141_O_2_1_1),
    .O_2_1_2(n141_O_2_1_2),
    .O_2_2_0(n141_O_2_2_0),
    .O_2_2_1(n141_O_2_2_1),
    .O_2_2_2(n141_O_2_2_2),
    .O_3_0_0(n141_O_3_0_0),
    .O_3_0_1(n141_O_3_0_1),
    .O_3_0_2(n141_O_3_0_2),
    .O_3_1_0(n141_O_3_1_0),
    .O_3_1_1(n141_O_3_1_1),
    .O_3_1_2(n141_O_3_1_2),
    .O_3_2_0(n141_O_3_2_0),
    .O_3_2_1(n141_O_3_2_1),
    .O_3_2_2(n141_O_3_2_2),
    .O_4_0_0(n141_O_4_0_0),
    .O_4_0_1(n141_O_4_0_1),
    .O_4_0_2(n141_O_4_0_2),
    .O_4_1_0(n141_O_4_1_0),
    .O_4_1_1(n141_O_4_1_1),
    .O_4_1_2(n141_O_4_1_2),
    .O_4_2_0(n141_O_4_2_0),
    .O_4_2_1(n141_O_4_2_1),
    .O_4_2_2(n141_O_4_2_2),
    .O_5_0_0(n141_O_5_0_0),
    .O_5_0_1(n141_O_5_0_1),
    .O_5_0_2(n141_O_5_0_2),
    .O_5_1_0(n141_O_5_1_0),
    .O_5_1_1(n141_O_5_1_1),
    .O_5_1_2(n141_O_5_1_2),
    .O_5_2_0(n141_O_5_2_0),
    .O_5_2_1(n141_O_5_2_1),
    .O_5_2_2(n141_O_5_2_2),
    .O_6_0_0(n141_O_6_0_0),
    .O_6_0_1(n141_O_6_0_1),
    .O_6_0_2(n141_O_6_0_2),
    .O_6_1_0(n141_O_6_1_0),
    .O_6_1_1(n141_O_6_1_1),
    .O_6_1_2(n141_O_6_1_2),
    .O_6_2_0(n141_O_6_2_0),
    .O_6_2_1(n141_O_6_2_1),
    .O_6_2_2(n141_O_6_2_2),
    .O_7_0_0(n141_O_7_0_0),
    .O_7_0_1(n141_O_7_0_1),
    .O_7_0_2(n141_O_7_0_2),
    .O_7_1_0(n141_O_7_1_0),
    .O_7_1_1(n141_O_7_1_1),
    .O_7_1_2(n141_O_7_1_2),
    .O_7_2_0(n141_O_7_2_0),
    .O_7_2_1(n141_O_7_2_1),
    .O_7_2_2(n141_O_7_2_2),
    .O_8_0_0(n141_O_8_0_0),
    .O_8_0_1(n141_O_8_0_1),
    .O_8_0_2(n141_O_8_0_2),
    .O_8_1_0(n141_O_8_1_0),
    .O_8_1_1(n141_O_8_1_1),
    .O_8_1_2(n141_O_8_1_2),
    .O_8_2_0(n141_O_8_2_0),
    .O_8_2_1(n141_O_8_2_1),
    .O_8_2_2(n141_O_8_2_2),
    .O_9_0_0(n141_O_9_0_0),
    .O_9_0_1(n141_O_9_0_1),
    .O_9_0_2(n141_O_9_0_2),
    .O_9_1_0(n141_O_9_1_0),
    .O_9_1_1(n141_O_9_1_1),
    .O_9_1_2(n141_O_9_1_2),
    .O_9_2_0(n141_O_9_2_0),
    .O_9_2_1(n141_O_9_2_1),
    .O_9_2_2(n141_O_9_2_2),
    .O_10_0_0(n141_O_10_0_0),
    .O_10_0_1(n141_O_10_0_1),
    .O_10_0_2(n141_O_10_0_2),
    .O_10_1_0(n141_O_10_1_0),
    .O_10_1_1(n141_O_10_1_1),
    .O_10_1_2(n141_O_10_1_2),
    .O_10_2_0(n141_O_10_2_0),
    .O_10_2_1(n141_O_10_2_1),
    .O_10_2_2(n141_O_10_2_2),
    .O_11_0_0(n141_O_11_0_0),
    .O_11_0_1(n141_O_11_0_1),
    .O_11_0_2(n141_O_11_0_2),
    .O_11_1_0(n141_O_11_1_0),
    .O_11_1_1(n141_O_11_1_1),
    .O_11_1_2(n141_O_11_1_2),
    .O_11_2_0(n141_O_11_2_0),
    .O_11_2_1(n141_O_11_2_1),
    .O_11_2_2(n141_O_11_2_2),
    .O_12_0_0(n141_O_12_0_0),
    .O_12_0_1(n141_O_12_0_1),
    .O_12_0_2(n141_O_12_0_2),
    .O_12_1_0(n141_O_12_1_0),
    .O_12_1_1(n141_O_12_1_1),
    .O_12_1_2(n141_O_12_1_2),
    .O_12_2_0(n141_O_12_2_0),
    .O_12_2_1(n141_O_12_2_1),
    .O_12_2_2(n141_O_12_2_2),
    .O_13_0_0(n141_O_13_0_0),
    .O_13_0_1(n141_O_13_0_1),
    .O_13_0_2(n141_O_13_0_2),
    .O_13_1_0(n141_O_13_1_0),
    .O_13_1_1(n141_O_13_1_1),
    .O_13_1_2(n141_O_13_1_2),
    .O_13_2_0(n141_O_13_2_0),
    .O_13_2_1(n141_O_13_2_1),
    .O_13_2_2(n141_O_13_2_2),
    .O_14_0_0(n141_O_14_0_0),
    .O_14_0_1(n141_O_14_0_1),
    .O_14_0_2(n141_O_14_0_2),
    .O_14_1_0(n141_O_14_1_0),
    .O_14_1_1(n141_O_14_1_1),
    .O_14_1_2(n141_O_14_1_2),
    .O_14_2_0(n141_O_14_2_0),
    .O_14_2_1(n141_O_14_2_1),
    .O_14_2_2(n141_O_14_2_2),
    .O_15_0_0(n141_O_15_0_0),
    .O_15_0_1(n141_O_15_0_1),
    .O_15_0_2(n141_O_15_0_2),
    .O_15_1_0(n141_O_15_1_0),
    .O_15_1_1(n141_O_15_1_1),
    .O_15_1_2(n141_O_15_1_2),
    .O_15_2_0(n141_O_15_2_0),
    .O_15_2_1(n141_O_15_2_1),
    .O_15_2_2(n141_O_15_2_2)
  );
  MapT_4 n183 ( // @[Top.scala 174:22]
    .clock(n183_clock),
    .reset(n183_reset),
    .valid_up(n183_valid_up),
    .valid_down(n183_valid_down),
    .I_0_0_0(n183_I_0_0_0),
    .I_0_0_1(n183_I_0_0_1),
    .I_0_0_2(n183_I_0_0_2),
    .I_0_1_0(n183_I_0_1_0),
    .I_0_1_1(n183_I_0_1_1),
    .I_0_1_2(n183_I_0_1_2),
    .I_0_2_0(n183_I_0_2_0),
    .I_0_2_1(n183_I_0_2_1),
    .I_0_2_2(n183_I_0_2_2),
    .I_1_0_0(n183_I_1_0_0),
    .I_1_0_1(n183_I_1_0_1),
    .I_1_0_2(n183_I_1_0_2),
    .I_1_1_0(n183_I_1_1_0),
    .I_1_1_1(n183_I_1_1_1),
    .I_1_1_2(n183_I_1_1_2),
    .I_1_2_0(n183_I_1_2_0),
    .I_1_2_1(n183_I_1_2_1),
    .I_1_2_2(n183_I_1_2_2),
    .I_2_0_0(n183_I_2_0_0),
    .I_2_0_1(n183_I_2_0_1),
    .I_2_0_2(n183_I_2_0_2),
    .I_2_1_0(n183_I_2_1_0),
    .I_2_1_1(n183_I_2_1_1),
    .I_2_1_2(n183_I_2_1_2),
    .I_2_2_0(n183_I_2_2_0),
    .I_2_2_1(n183_I_2_2_1),
    .I_2_2_2(n183_I_2_2_2),
    .I_3_0_0(n183_I_3_0_0),
    .I_3_0_1(n183_I_3_0_1),
    .I_3_0_2(n183_I_3_0_2),
    .I_3_1_0(n183_I_3_1_0),
    .I_3_1_1(n183_I_3_1_1),
    .I_3_1_2(n183_I_3_1_2),
    .I_3_2_0(n183_I_3_2_0),
    .I_3_2_1(n183_I_3_2_1),
    .I_3_2_2(n183_I_3_2_2),
    .I_4_0_0(n183_I_4_0_0),
    .I_4_0_1(n183_I_4_0_1),
    .I_4_0_2(n183_I_4_0_2),
    .I_4_1_0(n183_I_4_1_0),
    .I_4_1_1(n183_I_4_1_1),
    .I_4_1_2(n183_I_4_1_2),
    .I_4_2_0(n183_I_4_2_0),
    .I_4_2_1(n183_I_4_2_1),
    .I_4_2_2(n183_I_4_2_2),
    .I_5_0_0(n183_I_5_0_0),
    .I_5_0_1(n183_I_5_0_1),
    .I_5_0_2(n183_I_5_0_2),
    .I_5_1_0(n183_I_5_1_0),
    .I_5_1_1(n183_I_5_1_1),
    .I_5_1_2(n183_I_5_1_2),
    .I_5_2_0(n183_I_5_2_0),
    .I_5_2_1(n183_I_5_2_1),
    .I_5_2_2(n183_I_5_2_2),
    .I_6_0_0(n183_I_6_0_0),
    .I_6_0_1(n183_I_6_0_1),
    .I_6_0_2(n183_I_6_0_2),
    .I_6_1_0(n183_I_6_1_0),
    .I_6_1_1(n183_I_6_1_1),
    .I_6_1_2(n183_I_6_1_2),
    .I_6_2_0(n183_I_6_2_0),
    .I_6_2_1(n183_I_6_2_1),
    .I_6_2_2(n183_I_6_2_2),
    .I_7_0_0(n183_I_7_0_0),
    .I_7_0_1(n183_I_7_0_1),
    .I_7_0_2(n183_I_7_0_2),
    .I_7_1_0(n183_I_7_1_0),
    .I_7_1_1(n183_I_7_1_1),
    .I_7_1_2(n183_I_7_1_2),
    .I_7_2_0(n183_I_7_2_0),
    .I_7_2_1(n183_I_7_2_1),
    .I_7_2_2(n183_I_7_2_2),
    .I_8_0_0(n183_I_8_0_0),
    .I_8_0_1(n183_I_8_0_1),
    .I_8_0_2(n183_I_8_0_2),
    .I_8_1_0(n183_I_8_1_0),
    .I_8_1_1(n183_I_8_1_1),
    .I_8_1_2(n183_I_8_1_2),
    .I_8_2_0(n183_I_8_2_0),
    .I_8_2_1(n183_I_8_2_1),
    .I_8_2_2(n183_I_8_2_2),
    .I_9_0_0(n183_I_9_0_0),
    .I_9_0_1(n183_I_9_0_1),
    .I_9_0_2(n183_I_9_0_2),
    .I_9_1_0(n183_I_9_1_0),
    .I_9_1_1(n183_I_9_1_1),
    .I_9_1_2(n183_I_9_1_2),
    .I_9_2_0(n183_I_9_2_0),
    .I_9_2_1(n183_I_9_2_1),
    .I_9_2_2(n183_I_9_2_2),
    .I_10_0_0(n183_I_10_0_0),
    .I_10_0_1(n183_I_10_0_1),
    .I_10_0_2(n183_I_10_0_2),
    .I_10_1_0(n183_I_10_1_0),
    .I_10_1_1(n183_I_10_1_1),
    .I_10_1_2(n183_I_10_1_2),
    .I_10_2_0(n183_I_10_2_0),
    .I_10_2_1(n183_I_10_2_1),
    .I_10_2_2(n183_I_10_2_2),
    .I_11_0_0(n183_I_11_0_0),
    .I_11_0_1(n183_I_11_0_1),
    .I_11_0_2(n183_I_11_0_2),
    .I_11_1_0(n183_I_11_1_0),
    .I_11_1_1(n183_I_11_1_1),
    .I_11_1_2(n183_I_11_1_2),
    .I_11_2_0(n183_I_11_2_0),
    .I_11_2_1(n183_I_11_2_1),
    .I_11_2_2(n183_I_11_2_2),
    .I_12_0_0(n183_I_12_0_0),
    .I_12_0_1(n183_I_12_0_1),
    .I_12_0_2(n183_I_12_0_2),
    .I_12_1_0(n183_I_12_1_0),
    .I_12_1_1(n183_I_12_1_1),
    .I_12_1_2(n183_I_12_1_2),
    .I_12_2_0(n183_I_12_2_0),
    .I_12_2_1(n183_I_12_2_1),
    .I_12_2_2(n183_I_12_2_2),
    .I_13_0_0(n183_I_13_0_0),
    .I_13_0_1(n183_I_13_0_1),
    .I_13_0_2(n183_I_13_0_2),
    .I_13_1_0(n183_I_13_1_0),
    .I_13_1_1(n183_I_13_1_1),
    .I_13_1_2(n183_I_13_1_2),
    .I_13_2_0(n183_I_13_2_0),
    .I_13_2_1(n183_I_13_2_1),
    .I_13_2_2(n183_I_13_2_2),
    .I_14_0_0(n183_I_14_0_0),
    .I_14_0_1(n183_I_14_0_1),
    .I_14_0_2(n183_I_14_0_2),
    .I_14_1_0(n183_I_14_1_0),
    .I_14_1_1(n183_I_14_1_1),
    .I_14_1_2(n183_I_14_1_2),
    .I_14_2_0(n183_I_14_2_0),
    .I_14_2_1(n183_I_14_2_1),
    .I_14_2_2(n183_I_14_2_2),
    .I_15_0_0(n183_I_15_0_0),
    .I_15_0_1(n183_I_15_0_1),
    .I_15_0_2(n183_I_15_0_2),
    .I_15_1_0(n183_I_15_1_0),
    .I_15_1_1(n183_I_15_1_1),
    .I_15_1_2(n183_I_15_1_2),
    .I_15_2_0(n183_I_15_2_0),
    .I_15_2_1(n183_I_15_2_1),
    .I_15_2_2(n183_I_15_2_2),
    .O_0_0_0(n183_O_0_0_0),
    .O_1_0_0(n183_O_1_0_0),
    .O_2_0_0(n183_O_2_0_0),
    .O_3_0_0(n183_O_3_0_0),
    .O_4_0_0(n183_O_4_0_0),
    .O_5_0_0(n183_O_5_0_0),
    .O_6_0_0(n183_O_6_0_0),
    .O_7_0_0(n183_O_7_0_0),
    .O_8_0_0(n183_O_8_0_0),
    .O_9_0_0(n183_O_9_0_0),
    .O_10_0_0(n183_O_10_0_0),
    .O_11_0_0(n183_O_11_0_0),
    .O_12_0_0(n183_O_12_0_0),
    .O_13_0_0(n183_O_13_0_0),
    .O_14_0_0(n183_O_14_0_0),
    .O_15_0_0(n183_O_15_0_0)
  );
  FIFO_1 n184 ( // @[Top.scala 177:22]
    .clock(n184_clock),
    .reset(n184_reset),
    .valid_up(n184_valid_up),
    .valid_down(n184_valid_down),
    .I_0_0_0(n184_I_0_0_0),
    .I_1_0_0(n184_I_1_0_0),
    .I_2_0_0(n184_I_2_0_0),
    .I_3_0_0(n184_I_3_0_0),
    .I_4_0_0(n184_I_4_0_0),
    .I_5_0_0(n184_I_5_0_0),
    .I_6_0_0(n184_I_6_0_0),
    .I_7_0_0(n184_I_7_0_0),
    .I_8_0_0(n184_I_8_0_0),
    .I_9_0_0(n184_I_9_0_0),
    .I_10_0_0(n184_I_10_0_0),
    .I_11_0_0(n184_I_11_0_0),
    .I_12_0_0(n184_I_12_0_0),
    .I_13_0_0(n184_I_13_0_0),
    .I_14_0_0(n184_I_14_0_0),
    .I_15_0_0(n184_I_15_0_0),
    .O_0_0_0(n184_O_0_0_0),
    .O_1_0_0(n184_O_1_0_0),
    .O_2_0_0(n184_O_2_0_0),
    .O_3_0_0(n184_O_3_0_0),
    .O_4_0_0(n184_O_4_0_0),
    .O_5_0_0(n184_O_5_0_0),
    .O_6_0_0(n184_O_6_0_0),
    .O_7_0_0(n184_O_7_0_0),
    .O_8_0_0(n184_O_8_0_0),
    .O_9_0_0(n184_O_9_0_0),
    .O_10_0_0(n184_O_10_0_0),
    .O_11_0_0(n184_O_11_0_0),
    .O_12_0_0(n184_O_12_0_0),
    .O_13_0_0(n184_O_13_0_0),
    .O_14_0_0(n184_O_14_0_0),
    .O_15_0_0(n184_O_15_0_0)
  );
  Map2T_8 n185 ( // @[Top.scala 180:22]
    .clock(n185_clock),
    .reset(n185_reset),
    .valid_up(n185_valid_up),
    .valid_down(n185_valid_down),
    .I0_0_0_0(n185_I0_0_0_0),
    .I0_1_0_0(n185_I0_1_0_0),
    .I0_2_0_0(n185_I0_2_0_0),
    .I0_3_0_0(n185_I0_3_0_0),
    .I0_4_0_0(n185_I0_4_0_0),
    .I0_5_0_0(n185_I0_5_0_0),
    .I0_6_0_0(n185_I0_6_0_0),
    .I0_7_0_0(n185_I0_7_0_0),
    .I0_8_0_0(n185_I0_8_0_0),
    .I0_9_0_0(n185_I0_9_0_0),
    .I0_10_0_0(n185_I0_10_0_0),
    .I0_11_0_0(n185_I0_11_0_0),
    .I0_12_0_0(n185_I0_12_0_0),
    .I0_13_0_0(n185_I0_13_0_0),
    .I0_14_0_0(n185_I0_14_0_0),
    .I0_15_0_0(n185_I0_15_0_0),
    .I1_0_0_0(n185_I1_0_0_0),
    .I1_1_0_0(n185_I1_1_0_0),
    .I1_2_0_0(n185_I1_2_0_0),
    .I1_3_0_0(n185_I1_3_0_0),
    .I1_4_0_0(n185_I1_4_0_0),
    .I1_5_0_0(n185_I1_5_0_0),
    .I1_6_0_0(n185_I1_6_0_0),
    .I1_7_0_0(n185_I1_7_0_0),
    .I1_8_0_0(n185_I1_8_0_0),
    .I1_9_0_0(n185_I1_9_0_0),
    .I1_10_0_0(n185_I1_10_0_0),
    .I1_11_0_0(n185_I1_11_0_0),
    .I1_12_0_0(n185_I1_12_0_0),
    .I1_13_0_0(n185_I1_13_0_0),
    .I1_14_0_0(n185_I1_14_0_0),
    .I1_15_0_0(n185_I1_15_0_0),
    .O_0_0_0(n185_O_0_0_0),
    .O_1_0_0(n185_O_1_0_0),
    .O_2_0_0(n185_O_2_0_0),
    .O_3_0_0(n185_O_3_0_0),
    .O_4_0_0(n185_O_4_0_0),
    .O_5_0_0(n185_O_5_0_0),
    .O_6_0_0(n185_O_6_0_0),
    .O_7_0_0(n185_O_7_0_0),
    .O_8_0_0(n185_O_8_0_0),
    .O_9_0_0(n185_O_9_0_0),
    .O_10_0_0(n185_O_10_0_0),
    .O_11_0_0(n185_O_11_0_0),
    .O_12_0_0(n185_O_12_0_0),
    .O_13_0_0(n185_O_13_0_0),
    .O_14_0_0(n185_O_14_0_0),
    .O_15_0_0(n185_O_15_0_0)
  );
  FIFO n217 ( // @[Top.scala 184:22]
    .clock(n217_clock),
    .valid_up(n217_valid_up),
    .valid_down(n217_valid_down),
    .I_0_0_0(n217_I_0_0_0),
    .I_1_0_0(n217_I_1_0_0),
    .I_2_0_0(n217_I_2_0_0),
    .I_3_0_0(n217_I_3_0_0),
    .I_4_0_0(n217_I_4_0_0),
    .I_5_0_0(n217_I_5_0_0),
    .I_6_0_0(n217_I_6_0_0),
    .I_7_0_0(n217_I_7_0_0),
    .I_8_0_0(n217_I_8_0_0),
    .I_9_0_0(n217_I_9_0_0),
    .I_10_0_0(n217_I_10_0_0),
    .I_11_0_0(n217_I_11_0_0),
    .I_12_0_0(n217_I_12_0_0),
    .I_13_0_0(n217_I_13_0_0),
    .I_14_0_0(n217_I_14_0_0),
    .I_15_0_0(n217_I_15_0_0),
    .O_0_0_0(n217_O_0_0_0),
    .O_1_0_0(n217_O_1_0_0),
    .O_2_0_0(n217_O_2_0_0),
    .O_3_0_0(n217_O_3_0_0),
    .O_4_0_0(n217_O_4_0_0),
    .O_5_0_0(n217_O_5_0_0),
    .O_6_0_0(n217_O_6_0_0),
    .O_7_0_0(n217_O_7_0_0),
    .O_8_0_0(n217_O_8_0_0),
    .O_9_0_0(n217_O_9_0_0),
    .O_10_0_0(n217_O_10_0_0),
    .O_11_0_0(n217_O_11_0_0),
    .O_12_0_0(n217_O_12_0_0),
    .O_13_0_0(n217_O_13_0_0),
    .O_14_0_0(n217_O_14_0_0),
    .O_15_0_0(n217_O_15_0_0)
  );
  FIFO n218 ( // @[Top.scala 187:22]
    .clock(n218_clock),
    .valid_up(n218_valid_up),
    .valid_down(n218_valid_down),
    .I_0_0_0(n218_I_0_0_0),
    .I_1_0_0(n218_I_1_0_0),
    .I_2_0_0(n218_I_2_0_0),
    .I_3_0_0(n218_I_3_0_0),
    .I_4_0_0(n218_I_4_0_0),
    .I_5_0_0(n218_I_5_0_0),
    .I_6_0_0(n218_I_6_0_0),
    .I_7_0_0(n218_I_7_0_0),
    .I_8_0_0(n218_I_8_0_0),
    .I_9_0_0(n218_I_9_0_0),
    .I_10_0_0(n218_I_10_0_0),
    .I_11_0_0(n218_I_11_0_0),
    .I_12_0_0(n218_I_12_0_0),
    .I_13_0_0(n218_I_13_0_0),
    .I_14_0_0(n218_I_14_0_0),
    .I_15_0_0(n218_I_15_0_0),
    .O_0_0_0(n218_O_0_0_0),
    .O_1_0_0(n218_O_1_0_0),
    .O_2_0_0(n218_O_2_0_0),
    .O_3_0_0(n218_O_3_0_0),
    .O_4_0_0(n218_O_4_0_0),
    .O_5_0_0(n218_O_5_0_0),
    .O_6_0_0(n218_O_6_0_0),
    .O_7_0_0(n218_O_7_0_0),
    .O_8_0_0(n218_O_8_0_0),
    .O_9_0_0(n218_O_9_0_0),
    .O_10_0_0(n218_O_10_0_0),
    .O_11_0_0(n218_O_11_0_0),
    .O_12_0_0(n218_O_12_0_0),
    .O_13_0_0(n218_O_13_0_0),
    .O_14_0_0(n218_O_14_0_0),
    .O_15_0_0(n218_O_15_0_0)
  );
  FIFO n219 ( // @[Top.scala 190:22]
    .clock(n219_clock),
    .valid_up(n219_valid_up),
    .valid_down(n219_valid_down),
    .I_0_0_0(n219_I_0_0_0),
    .I_1_0_0(n219_I_1_0_0),
    .I_2_0_0(n219_I_2_0_0),
    .I_3_0_0(n219_I_3_0_0),
    .I_4_0_0(n219_I_4_0_0),
    .I_5_0_0(n219_I_5_0_0),
    .I_6_0_0(n219_I_6_0_0),
    .I_7_0_0(n219_I_7_0_0),
    .I_8_0_0(n219_I_8_0_0),
    .I_9_0_0(n219_I_9_0_0),
    .I_10_0_0(n219_I_10_0_0),
    .I_11_0_0(n219_I_11_0_0),
    .I_12_0_0(n219_I_12_0_0),
    .I_13_0_0(n219_I_13_0_0),
    .I_14_0_0(n219_I_14_0_0),
    .I_15_0_0(n219_I_15_0_0),
    .O_0_0_0(n219_O_0_0_0),
    .O_1_0_0(n219_O_1_0_0),
    .O_2_0_0(n219_O_2_0_0),
    .O_3_0_0(n219_O_3_0_0),
    .O_4_0_0(n219_O_4_0_0),
    .O_5_0_0(n219_O_5_0_0),
    .O_6_0_0(n219_O_6_0_0),
    .O_7_0_0(n219_O_7_0_0),
    .O_8_0_0(n219_O_8_0_0),
    .O_9_0_0(n219_O_9_0_0),
    .O_10_0_0(n219_O_10_0_0),
    .O_11_0_0(n219_O_11_0_0),
    .O_12_0_0(n219_O_12_0_0),
    .O_13_0_0(n219_O_13_0_0),
    .O_14_0_0(n219_O_14_0_0),
    .O_15_0_0(n219_O_15_0_0)
  );
  assign valid_down = n219_valid_down; // @[Top.scala 194:16]
  assign O_0_0_0 = n219_O_0_0_0; // @[Top.scala 193:7]
  assign O_1_0_0 = n219_O_1_0_0; // @[Top.scala 193:7]
  assign O_2_0_0 = n219_O_2_0_0; // @[Top.scala 193:7]
  assign O_3_0_0 = n219_O_3_0_0; // @[Top.scala 193:7]
  assign O_4_0_0 = n219_O_4_0_0; // @[Top.scala 193:7]
  assign O_5_0_0 = n219_O_5_0_0; // @[Top.scala 193:7]
  assign O_6_0_0 = n219_O_6_0_0; // @[Top.scala 193:7]
  assign O_7_0_0 = n219_O_7_0_0; // @[Top.scala 193:7]
  assign O_8_0_0 = n219_O_8_0_0; // @[Top.scala 193:7]
  assign O_9_0_0 = n219_O_9_0_0; // @[Top.scala 193:7]
  assign O_10_0_0 = n219_O_10_0_0; // @[Top.scala 193:7]
  assign O_11_0_0 = n219_O_11_0_0; // @[Top.scala 193:7]
  assign O_12_0_0 = n219_O_12_0_0; // @[Top.scala 193:7]
  assign O_13_0_0 = n219_O_13_0_0; // @[Top.scala 193:7]
  assign O_14_0_0 = n219_O_14_0_0; // @[Top.scala 193:7]
  assign O_15_0_0 = n219_O_15_0_0; // @[Top.scala 193:7]
  assign n1_clock = clock;
  assign n1_valid_up = valid_up; // @[Top.scala 105:17]
  assign n1_I_0_0_0 = I_0_0_0; // @[Top.scala 104:10]
  assign n1_I_1_0_0 = I_1_0_0; // @[Top.scala 104:10]
  assign n1_I_2_0_0 = I_2_0_0; // @[Top.scala 104:10]
  assign n1_I_3_0_0 = I_3_0_0; // @[Top.scala 104:10]
  assign n1_I_4_0_0 = I_4_0_0; // @[Top.scala 104:10]
  assign n1_I_5_0_0 = I_5_0_0; // @[Top.scala 104:10]
  assign n1_I_6_0_0 = I_6_0_0; // @[Top.scala 104:10]
  assign n1_I_7_0_0 = I_7_0_0; // @[Top.scala 104:10]
  assign n1_I_8_0_0 = I_8_0_0; // @[Top.scala 104:10]
  assign n1_I_9_0_0 = I_9_0_0; // @[Top.scala 104:10]
  assign n1_I_10_0_0 = I_10_0_0; // @[Top.scala 104:10]
  assign n1_I_11_0_0 = I_11_0_0; // @[Top.scala 104:10]
  assign n1_I_12_0_0 = I_12_0_0; // @[Top.scala 104:10]
  assign n1_I_13_0_0 = I_13_0_0; // @[Top.scala 104:10]
  assign n1_I_14_0_0 = I_14_0_0; // @[Top.scala 104:10]
  assign n1_I_15_0_0 = I_15_0_0; // @[Top.scala 104:10]
  assign n2_clock = clock;
  assign n2_reset = reset;
  assign n2_valid_up = n1_valid_down; // @[Top.scala 108:17]
  assign n2_I_0_0_0 = n1_O_0_0_0; // @[Top.scala 107:10]
  assign n2_I_1_0_0 = n1_O_1_0_0; // @[Top.scala 107:10]
  assign n2_I_2_0_0 = n1_O_2_0_0; // @[Top.scala 107:10]
  assign n2_I_3_0_0 = n1_O_3_0_0; // @[Top.scala 107:10]
  assign n2_I_4_0_0 = n1_O_4_0_0; // @[Top.scala 107:10]
  assign n2_I_5_0_0 = n1_O_5_0_0; // @[Top.scala 107:10]
  assign n2_I_6_0_0 = n1_O_6_0_0; // @[Top.scala 107:10]
  assign n2_I_7_0_0 = n1_O_7_0_0; // @[Top.scala 107:10]
  assign n2_I_8_0_0 = n1_O_8_0_0; // @[Top.scala 107:10]
  assign n2_I_9_0_0 = n1_O_9_0_0; // @[Top.scala 107:10]
  assign n2_I_10_0_0 = n1_O_10_0_0; // @[Top.scala 107:10]
  assign n2_I_11_0_0 = n1_O_11_0_0; // @[Top.scala 107:10]
  assign n2_I_12_0_0 = n1_O_12_0_0; // @[Top.scala 107:10]
  assign n2_I_13_0_0 = n1_O_13_0_0; // @[Top.scala 107:10]
  assign n2_I_14_0_0 = n1_O_14_0_0; // @[Top.scala 107:10]
  assign n2_I_15_0_0 = n1_O_15_0_0; // @[Top.scala 107:10]
  assign n3_clock = clock;
  assign n3_reset = reset;
  assign n3_valid_up = n2_valid_down; // @[Top.scala 111:17]
  assign n3_I_0_0_0 = n2_O_0_0_0; // @[Top.scala 110:10]
  assign n3_I_1_0_0 = n2_O_1_0_0; // @[Top.scala 110:10]
  assign n3_I_2_0_0 = n2_O_2_0_0; // @[Top.scala 110:10]
  assign n3_I_3_0_0 = n2_O_3_0_0; // @[Top.scala 110:10]
  assign n3_I_4_0_0 = n2_O_4_0_0; // @[Top.scala 110:10]
  assign n3_I_5_0_0 = n2_O_5_0_0; // @[Top.scala 110:10]
  assign n3_I_6_0_0 = n2_O_6_0_0; // @[Top.scala 110:10]
  assign n3_I_7_0_0 = n2_O_7_0_0; // @[Top.scala 110:10]
  assign n3_I_8_0_0 = n2_O_8_0_0; // @[Top.scala 110:10]
  assign n3_I_9_0_0 = n2_O_9_0_0; // @[Top.scala 110:10]
  assign n3_I_10_0_0 = n2_O_10_0_0; // @[Top.scala 110:10]
  assign n3_I_11_0_0 = n2_O_11_0_0; // @[Top.scala 110:10]
  assign n3_I_12_0_0 = n2_O_12_0_0; // @[Top.scala 110:10]
  assign n3_I_13_0_0 = n2_O_13_0_0; // @[Top.scala 110:10]
  assign n3_I_14_0_0 = n2_O_14_0_0; // @[Top.scala 110:10]
  assign n3_I_15_0_0 = n2_O_15_0_0; // @[Top.scala 110:10]
  assign n4_clock = clock;
  assign n4_valid_up = n3_valid_down; // @[Top.scala 114:17]
  assign n4_I_0_0_0 = n3_O_0_0_0; // @[Top.scala 113:10]
  assign n4_I_1_0_0 = n3_O_1_0_0; // @[Top.scala 113:10]
  assign n4_I_2_0_0 = n3_O_2_0_0; // @[Top.scala 113:10]
  assign n4_I_3_0_0 = n3_O_3_0_0; // @[Top.scala 113:10]
  assign n4_I_4_0_0 = n3_O_4_0_0; // @[Top.scala 113:10]
  assign n4_I_5_0_0 = n3_O_5_0_0; // @[Top.scala 113:10]
  assign n4_I_6_0_0 = n3_O_6_0_0; // @[Top.scala 113:10]
  assign n4_I_7_0_0 = n3_O_7_0_0; // @[Top.scala 113:10]
  assign n4_I_8_0_0 = n3_O_8_0_0; // @[Top.scala 113:10]
  assign n4_I_9_0_0 = n3_O_9_0_0; // @[Top.scala 113:10]
  assign n4_I_10_0_0 = n3_O_10_0_0; // @[Top.scala 113:10]
  assign n4_I_11_0_0 = n3_O_11_0_0; // @[Top.scala 113:10]
  assign n4_I_12_0_0 = n3_O_12_0_0; // @[Top.scala 113:10]
  assign n4_I_13_0_0 = n3_O_13_0_0; // @[Top.scala 113:10]
  assign n4_I_14_0_0 = n3_O_14_0_0; // @[Top.scala 113:10]
  assign n4_I_15_0_0 = n3_O_15_0_0; // @[Top.scala 113:10]
  assign n5_clock = clock;
  assign n5_valid_up = n4_valid_down; // @[Top.scala 117:17]
  assign n5_I_0_0_0 = n4_O_0_0_0; // @[Top.scala 116:10]
  assign n5_I_1_0_0 = n4_O_1_0_0; // @[Top.scala 116:10]
  assign n5_I_2_0_0 = n4_O_2_0_0; // @[Top.scala 116:10]
  assign n5_I_3_0_0 = n4_O_3_0_0; // @[Top.scala 116:10]
  assign n5_I_4_0_0 = n4_O_4_0_0; // @[Top.scala 116:10]
  assign n5_I_5_0_0 = n4_O_5_0_0; // @[Top.scala 116:10]
  assign n5_I_6_0_0 = n4_O_6_0_0; // @[Top.scala 116:10]
  assign n5_I_7_0_0 = n4_O_7_0_0; // @[Top.scala 116:10]
  assign n5_I_8_0_0 = n4_O_8_0_0; // @[Top.scala 116:10]
  assign n5_I_9_0_0 = n4_O_9_0_0; // @[Top.scala 116:10]
  assign n5_I_10_0_0 = n4_O_10_0_0; // @[Top.scala 116:10]
  assign n5_I_11_0_0 = n4_O_11_0_0; // @[Top.scala 116:10]
  assign n5_I_12_0_0 = n4_O_12_0_0; // @[Top.scala 116:10]
  assign n5_I_13_0_0 = n4_O_13_0_0; // @[Top.scala 116:10]
  assign n5_I_14_0_0 = n4_O_14_0_0; // @[Top.scala 116:10]
  assign n5_I_15_0_0 = n4_O_15_0_0; // @[Top.scala 116:10]
  assign n6_valid_up = n5_valid_down & n4_valid_down; // @[Top.scala 121:17]
  assign n6_I0_0_0_0 = n5_O_0_0_0; // @[Top.scala 119:11]
  assign n6_I0_1_0_0 = n5_O_1_0_0; // @[Top.scala 119:11]
  assign n6_I0_2_0_0 = n5_O_2_0_0; // @[Top.scala 119:11]
  assign n6_I0_3_0_0 = n5_O_3_0_0; // @[Top.scala 119:11]
  assign n6_I0_4_0_0 = n5_O_4_0_0; // @[Top.scala 119:11]
  assign n6_I0_5_0_0 = n5_O_5_0_0; // @[Top.scala 119:11]
  assign n6_I0_6_0_0 = n5_O_6_0_0; // @[Top.scala 119:11]
  assign n6_I0_7_0_0 = n5_O_7_0_0; // @[Top.scala 119:11]
  assign n6_I0_8_0_0 = n5_O_8_0_0; // @[Top.scala 119:11]
  assign n6_I0_9_0_0 = n5_O_9_0_0; // @[Top.scala 119:11]
  assign n6_I0_10_0_0 = n5_O_10_0_0; // @[Top.scala 119:11]
  assign n6_I0_11_0_0 = n5_O_11_0_0; // @[Top.scala 119:11]
  assign n6_I0_12_0_0 = n5_O_12_0_0; // @[Top.scala 119:11]
  assign n6_I0_13_0_0 = n5_O_13_0_0; // @[Top.scala 119:11]
  assign n6_I0_14_0_0 = n5_O_14_0_0; // @[Top.scala 119:11]
  assign n6_I0_15_0_0 = n5_O_15_0_0; // @[Top.scala 119:11]
  assign n6_I1_0_0_0 = n4_O_0_0_0; // @[Top.scala 120:11]
  assign n6_I1_1_0_0 = n4_O_1_0_0; // @[Top.scala 120:11]
  assign n6_I1_2_0_0 = n4_O_2_0_0; // @[Top.scala 120:11]
  assign n6_I1_3_0_0 = n4_O_3_0_0; // @[Top.scala 120:11]
  assign n6_I1_4_0_0 = n4_O_4_0_0; // @[Top.scala 120:11]
  assign n6_I1_5_0_0 = n4_O_5_0_0; // @[Top.scala 120:11]
  assign n6_I1_6_0_0 = n4_O_6_0_0; // @[Top.scala 120:11]
  assign n6_I1_7_0_0 = n4_O_7_0_0; // @[Top.scala 120:11]
  assign n6_I1_8_0_0 = n4_O_8_0_0; // @[Top.scala 120:11]
  assign n6_I1_9_0_0 = n4_O_9_0_0; // @[Top.scala 120:11]
  assign n6_I1_10_0_0 = n4_O_10_0_0; // @[Top.scala 120:11]
  assign n6_I1_11_0_0 = n4_O_11_0_0; // @[Top.scala 120:11]
  assign n6_I1_12_0_0 = n4_O_12_0_0; // @[Top.scala 120:11]
  assign n6_I1_13_0_0 = n4_O_13_0_0; // @[Top.scala 120:11]
  assign n6_I1_14_0_0 = n4_O_14_0_0; // @[Top.scala 120:11]
  assign n6_I1_15_0_0 = n4_O_15_0_0; // @[Top.scala 120:11]
  assign n19_valid_up = n6_valid_down & n3_valid_down; // @[Top.scala 125:18]
  assign n19_I0_0_0_0_0 = n6_O_0_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_0_0_0_1 = n6_O_0_0_0_1; // @[Top.scala 123:12]
  assign n19_I0_1_0_0_0 = n6_O_1_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_1_0_0_1 = n6_O_1_0_0_1; // @[Top.scala 123:12]
  assign n19_I0_2_0_0_0 = n6_O_2_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_2_0_0_1 = n6_O_2_0_0_1; // @[Top.scala 123:12]
  assign n19_I0_3_0_0_0 = n6_O_3_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_3_0_0_1 = n6_O_3_0_0_1; // @[Top.scala 123:12]
  assign n19_I0_4_0_0_0 = n6_O_4_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_4_0_0_1 = n6_O_4_0_0_1; // @[Top.scala 123:12]
  assign n19_I0_5_0_0_0 = n6_O_5_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_5_0_0_1 = n6_O_5_0_0_1; // @[Top.scala 123:12]
  assign n19_I0_6_0_0_0 = n6_O_6_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_6_0_0_1 = n6_O_6_0_0_1; // @[Top.scala 123:12]
  assign n19_I0_7_0_0_0 = n6_O_7_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_7_0_0_1 = n6_O_7_0_0_1; // @[Top.scala 123:12]
  assign n19_I0_8_0_0_0 = n6_O_8_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_8_0_0_1 = n6_O_8_0_0_1; // @[Top.scala 123:12]
  assign n19_I0_9_0_0_0 = n6_O_9_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_9_0_0_1 = n6_O_9_0_0_1; // @[Top.scala 123:12]
  assign n19_I0_10_0_0_0 = n6_O_10_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_10_0_0_1 = n6_O_10_0_0_1; // @[Top.scala 123:12]
  assign n19_I0_11_0_0_0 = n6_O_11_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_11_0_0_1 = n6_O_11_0_0_1; // @[Top.scala 123:12]
  assign n19_I0_12_0_0_0 = n6_O_12_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_12_0_0_1 = n6_O_12_0_0_1; // @[Top.scala 123:12]
  assign n19_I0_13_0_0_0 = n6_O_13_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_13_0_0_1 = n6_O_13_0_0_1; // @[Top.scala 123:12]
  assign n19_I0_14_0_0_0 = n6_O_14_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_14_0_0_1 = n6_O_14_0_0_1; // @[Top.scala 123:12]
  assign n19_I0_15_0_0_0 = n6_O_15_0_0_0; // @[Top.scala 123:12]
  assign n19_I0_15_0_0_1 = n6_O_15_0_0_1; // @[Top.scala 123:12]
  assign n19_I1_0_0_0 = n3_O_0_0_0; // @[Top.scala 124:12]
  assign n19_I1_1_0_0 = n3_O_1_0_0; // @[Top.scala 124:12]
  assign n19_I1_2_0_0 = n3_O_2_0_0; // @[Top.scala 124:12]
  assign n19_I1_3_0_0 = n3_O_3_0_0; // @[Top.scala 124:12]
  assign n19_I1_4_0_0 = n3_O_4_0_0; // @[Top.scala 124:12]
  assign n19_I1_5_0_0 = n3_O_5_0_0; // @[Top.scala 124:12]
  assign n19_I1_6_0_0 = n3_O_6_0_0; // @[Top.scala 124:12]
  assign n19_I1_7_0_0 = n3_O_7_0_0; // @[Top.scala 124:12]
  assign n19_I1_8_0_0 = n3_O_8_0_0; // @[Top.scala 124:12]
  assign n19_I1_9_0_0 = n3_O_9_0_0; // @[Top.scala 124:12]
  assign n19_I1_10_0_0 = n3_O_10_0_0; // @[Top.scala 124:12]
  assign n19_I1_11_0_0 = n3_O_11_0_0; // @[Top.scala 124:12]
  assign n19_I1_12_0_0 = n3_O_12_0_0; // @[Top.scala 124:12]
  assign n19_I1_13_0_0 = n3_O_13_0_0; // @[Top.scala 124:12]
  assign n19_I1_14_0_0 = n3_O_14_0_0; // @[Top.scala 124:12]
  assign n19_I1_15_0_0 = n3_O_15_0_0; // @[Top.scala 124:12]
  assign n40_valid_up = n19_valid_down; // @[Top.scala 128:18]
  assign n40_I_0_0_0_0 = n19_O_0_0_0_0; // @[Top.scala 127:11]
  assign n40_I_0_0_0_1 = n19_O_0_0_0_1; // @[Top.scala 127:11]
  assign n40_I_0_0_0_2 = n19_O_0_0_0_2; // @[Top.scala 127:11]
  assign n40_I_1_0_0_0 = n19_O_1_0_0_0; // @[Top.scala 127:11]
  assign n40_I_1_0_0_1 = n19_O_1_0_0_1; // @[Top.scala 127:11]
  assign n40_I_1_0_0_2 = n19_O_1_0_0_2; // @[Top.scala 127:11]
  assign n40_I_2_0_0_0 = n19_O_2_0_0_0; // @[Top.scala 127:11]
  assign n40_I_2_0_0_1 = n19_O_2_0_0_1; // @[Top.scala 127:11]
  assign n40_I_2_0_0_2 = n19_O_2_0_0_2; // @[Top.scala 127:11]
  assign n40_I_3_0_0_0 = n19_O_3_0_0_0; // @[Top.scala 127:11]
  assign n40_I_3_0_0_1 = n19_O_3_0_0_1; // @[Top.scala 127:11]
  assign n40_I_3_0_0_2 = n19_O_3_0_0_2; // @[Top.scala 127:11]
  assign n40_I_4_0_0_0 = n19_O_4_0_0_0; // @[Top.scala 127:11]
  assign n40_I_4_0_0_1 = n19_O_4_0_0_1; // @[Top.scala 127:11]
  assign n40_I_4_0_0_2 = n19_O_4_0_0_2; // @[Top.scala 127:11]
  assign n40_I_5_0_0_0 = n19_O_5_0_0_0; // @[Top.scala 127:11]
  assign n40_I_5_0_0_1 = n19_O_5_0_0_1; // @[Top.scala 127:11]
  assign n40_I_5_0_0_2 = n19_O_5_0_0_2; // @[Top.scala 127:11]
  assign n40_I_6_0_0_0 = n19_O_6_0_0_0; // @[Top.scala 127:11]
  assign n40_I_6_0_0_1 = n19_O_6_0_0_1; // @[Top.scala 127:11]
  assign n40_I_6_0_0_2 = n19_O_6_0_0_2; // @[Top.scala 127:11]
  assign n40_I_7_0_0_0 = n19_O_7_0_0_0; // @[Top.scala 127:11]
  assign n40_I_7_0_0_1 = n19_O_7_0_0_1; // @[Top.scala 127:11]
  assign n40_I_7_0_0_2 = n19_O_7_0_0_2; // @[Top.scala 127:11]
  assign n40_I_8_0_0_0 = n19_O_8_0_0_0; // @[Top.scala 127:11]
  assign n40_I_8_0_0_1 = n19_O_8_0_0_1; // @[Top.scala 127:11]
  assign n40_I_8_0_0_2 = n19_O_8_0_0_2; // @[Top.scala 127:11]
  assign n40_I_9_0_0_0 = n19_O_9_0_0_0; // @[Top.scala 127:11]
  assign n40_I_9_0_0_1 = n19_O_9_0_0_1; // @[Top.scala 127:11]
  assign n40_I_9_0_0_2 = n19_O_9_0_0_2; // @[Top.scala 127:11]
  assign n40_I_10_0_0_0 = n19_O_10_0_0_0; // @[Top.scala 127:11]
  assign n40_I_10_0_0_1 = n19_O_10_0_0_1; // @[Top.scala 127:11]
  assign n40_I_10_0_0_2 = n19_O_10_0_0_2; // @[Top.scala 127:11]
  assign n40_I_11_0_0_0 = n19_O_11_0_0_0; // @[Top.scala 127:11]
  assign n40_I_11_0_0_1 = n19_O_11_0_0_1; // @[Top.scala 127:11]
  assign n40_I_11_0_0_2 = n19_O_11_0_0_2; // @[Top.scala 127:11]
  assign n40_I_12_0_0_0 = n19_O_12_0_0_0; // @[Top.scala 127:11]
  assign n40_I_12_0_0_1 = n19_O_12_0_0_1; // @[Top.scala 127:11]
  assign n40_I_12_0_0_2 = n19_O_12_0_0_2; // @[Top.scala 127:11]
  assign n40_I_13_0_0_0 = n19_O_13_0_0_0; // @[Top.scala 127:11]
  assign n40_I_13_0_0_1 = n19_O_13_0_0_1; // @[Top.scala 127:11]
  assign n40_I_13_0_0_2 = n19_O_13_0_0_2; // @[Top.scala 127:11]
  assign n40_I_14_0_0_0 = n19_O_14_0_0_0; // @[Top.scala 127:11]
  assign n40_I_14_0_0_1 = n19_O_14_0_0_1; // @[Top.scala 127:11]
  assign n40_I_14_0_0_2 = n19_O_14_0_0_2; // @[Top.scala 127:11]
  assign n40_I_15_0_0_0 = n19_O_15_0_0_0; // @[Top.scala 127:11]
  assign n40_I_15_0_0_1 = n19_O_15_0_0_1; // @[Top.scala 127:11]
  assign n40_I_15_0_0_2 = n19_O_15_0_0_2; // @[Top.scala 127:11]
  assign n41_clock = clock;
  assign n41_valid_up = n2_valid_down; // @[Top.scala 131:18]
  assign n41_I_0_0_0 = n2_O_0_0_0; // @[Top.scala 130:11]
  assign n41_I_1_0_0 = n2_O_1_0_0; // @[Top.scala 130:11]
  assign n41_I_2_0_0 = n2_O_2_0_0; // @[Top.scala 130:11]
  assign n41_I_3_0_0 = n2_O_3_0_0; // @[Top.scala 130:11]
  assign n41_I_4_0_0 = n2_O_4_0_0; // @[Top.scala 130:11]
  assign n41_I_5_0_0 = n2_O_5_0_0; // @[Top.scala 130:11]
  assign n41_I_6_0_0 = n2_O_6_0_0; // @[Top.scala 130:11]
  assign n41_I_7_0_0 = n2_O_7_0_0; // @[Top.scala 130:11]
  assign n41_I_8_0_0 = n2_O_8_0_0; // @[Top.scala 130:11]
  assign n41_I_9_0_0 = n2_O_9_0_0; // @[Top.scala 130:11]
  assign n41_I_10_0_0 = n2_O_10_0_0; // @[Top.scala 130:11]
  assign n41_I_11_0_0 = n2_O_11_0_0; // @[Top.scala 130:11]
  assign n41_I_12_0_0 = n2_O_12_0_0; // @[Top.scala 130:11]
  assign n41_I_13_0_0 = n2_O_13_0_0; // @[Top.scala 130:11]
  assign n41_I_14_0_0 = n2_O_14_0_0; // @[Top.scala 130:11]
  assign n41_I_15_0_0 = n2_O_15_0_0; // @[Top.scala 130:11]
  assign n42_clock = clock;
  assign n42_valid_up = n41_valid_down; // @[Top.scala 134:18]
  assign n42_I_0_0_0 = n41_O_0_0_0; // @[Top.scala 133:11]
  assign n42_I_1_0_0 = n41_O_1_0_0; // @[Top.scala 133:11]
  assign n42_I_2_0_0 = n41_O_2_0_0; // @[Top.scala 133:11]
  assign n42_I_3_0_0 = n41_O_3_0_0; // @[Top.scala 133:11]
  assign n42_I_4_0_0 = n41_O_4_0_0; // @[Top.scala 133:11]
  assign n42_I_5_0_0 = n41_O_5_0_0; // @[Top.scala 133:11]
  assign n42_I_6_0_0 = n41_O_6_0_0; // @[Top.scala 133:11]
  assign n42_I_7_0_0 = n41_O_7_0_0; // @[Top.scala 133:11]
  assign n42_I_8_0_0 = n41_O_8_0_0; // @[Top.scala 133:11]
  assign n42_I_9_0_0 = n41_O_9_0_0; // @[Top.scala 133:11]
  assign n42_I_10_0_0 = n41_O_10_0_0; // @[Top.scala 133:11]
  assign n42_I_11_0_0 = n41_O_11_0_0; // @[Top.scala 133:11]
  assign n42_I_12_0_0 = n41_O_12_0_0; // @[Top.scala 133:11]
  assign n42_I_13_0_0 = n41_O_13_0_0; // @[Top.scala 133:11]
  assign n42_I_14_0_0 = n41_O_14_0_0; // @[Top.scala 133:11]
  assign n42_I_15_0_0 = n41_O_15_0_0; // @[Top.scala 133:11]
  assign n43_valid_up = n42_valid_down & n41_valid_down; // @[Top.scala 138:18]
  assign n43_I0_0_0_0 = n42_O_0_0_0; // @[Top.scala 136:12]
  assign n43_I0_1_0_0 = n42_O_1_0_0; // @[Top.scala 136:12]
  assign n43_I0_2_0_0 = n42_O_2_0_0; // @[Top.scala 136:12]
  assign n43_I0_3_0_0 = n42_O_3_0_0; // @[Top.scala 136:12]
  assign n43_I0_4_0_0 = n42_O_4_0_0; // @[Top.scala 136:12]
  assign n43_I0_5_0_0 = n42_O_5_0_0; // @[Top.scala 136:12]
  assign n43_I0_6_0_0 = n42_O_6_0_0; // @[Top.scala 136:12]
  assign n43_I0_7_0_0 = n42_O_7_0_0; // @[Top.scala 136:12]
  assign n43_I0_8_0_0 = n42_O_8_0_0; // @[Top.scala 136:12]
  assign n43_I0_9_0_0 = n42_O_9_0_0; // @[Top.scala 136:12]
  assign n43_I0_10_0_0 = n42_O_10_0_0; // @[Top.scala 136:12]
  assign n43_I0_11_0_0 = n42_O_11_0_0; // @[Top.scala 136:12]
  assign n43_I0_12_0_0 = n42_O_12_0_0; // @[Top.scala 136:12]
  assign n43_I0_13_0_0 = n42_O_13_0_0; // @[Top.scala 136:12]
  assign n43_I0_14_0_0 = n42_O_14_0_0; // @[Top.scala 136:12]
  assign n43_I0_15_0_0 = n42_O_15_0_0; // @[Top.scala 136:12]
  assign n43_I1_0_0_0 = n41_O_0_0_0; // @[Top.scala 137:12]
  assign n43_I1_1_0_0 = n41_O_1_0_0; // @[Top.scala 137:12]
  assign n43_I1_2_0_0 = n41_O_2_0_0; // @[Top.scala 137:12]
  assign n43_I1_3_0_0 = n41_O_3_0_0; // @[Top.scala 137:12]
  assign n43_I1_4_0_0 = n41_O_4_0_0; // @[Top.scala 137:12]
  assign n43_I1_5_0_0 = n41_O_5_0_0; // @[Top.scala 137:12]
  assign n43_I1_6_0_0 = n41_O_6_0_0; // @[Top.scala 137:12]
  assign n43_I1_7_0_0 = n41_O_7_0_0; // @[Top.scala 137:12]
  assign n43_I1_8_0_0 = n41_O_8_0_0; // @[Top.scala 137:12]
  assign n43_I1_9_0_0 = n41_O_9_0_0; // @[Top.scala 137:12]
  assign n43_I1_10_0_0 = n41_O_10_0_0; // @[Top.scala 137:12]
  assign n43_I1_11_0_0 = n41_O_11_0_0; // @[Top.scala 137:12]
  assign n43_I1_12_0_0 = n41_O_12_0_0; // @[Top.scala 137:12]
  assign n43_I1_13_0_0 = n41_O_13_0_0; // @[Top.scala 137:12]
  assign n43_I1_14_0_0 = n41_O_14_0_0; // @[Top.scala 137:12]
  assign n43_I1_15_0_0 = n41_O_15_0_0; // @[Top.scala 137:12]
  assign n56_valid_up = n43_valid_down & n2_valid_down; // @[Top.scala 142:18]
  assign n56_I0_0_0_0_0 = n43_O_0_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_0_0_0_1 = n43_O_0_0_0_1; // @[Top.scala 140:12]
  assign n56_I0_1_0_0_0 = n43_O_1_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_1_0_0_1 = n43_O_1_0_0_1; // @[Top.scala 140:12]
  assign n56_I0_2_0_0_0 = n43_O_2_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_2_0_0_1 = n43_O_2_0_0_1; // @[Top.scala 140:12]
  assign n56_I0_3_0_0_0 = n43_O_3_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_3_0_0_1 = n43_O_3_0_0_1; // @[Top.scala 140:12]
  assign n56_I0_4_0_0_0 = n43_O_4_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_4_0_0_1 = n43_O_4_0_0_1; // @[Top.scala 140:12]
  assign n56_I0_5_0_0_0 = n43_O_5_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_5_0_0_1 = n43_O_5_0_0_1; // @[Top.scala 140:12]
  assign n56_I0_6_0_0_0 = n43_O_6_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_6_0_0_1 = n43_O_6_0_0_1; // @[Top.scala 140:12]
  assign n56_I0_7_0_0_0 = n43_O_7_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_7_0_0_1 = n43_O_7_0_0_1; // @[Top.scala 140:12]
  assign n56_I0_8_0_0_0 = n43_O_8_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_8_0_0_1 = n43_O_8_0_0_1; // @[Top.scala 140:12]
  assign n56_I0_9_0_0_0 = n43_O_9_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_9_0_0_1 = n43_O_9_0_0_1; // @[Top.scala 140:12]
  assign n56_I0_10_0_0_0 = n43_O_10_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_10_0_0_1 = n43_O_10_0_0_1; // @[Top.scala 140:12]
  assign n56_I0_11_0_0_0 = n43_O_11_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_11_0_0_1 = n43_O_11_0_0_1; // @[Top.scala 140:12]
  assign n56_I0_12_0_0_0 = n43_O_12_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_12_0_0_1 = n43_O_12_0_0_1; // @[Top.scala 140:12]
  assign n56_I0_13_0_0_0 = n43_O_13_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_13_0_0_1 = n43_O_13_0_0_1; // @[Top.scala 140:12]
  assign n56_I0_14_0_0_0 = n43_O_14_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_14_0_0_1 = n43_O_14_0_0_1; // @[Top.scala 140:12]
  assign n56_I0_15_0_0_0 = n43_O_15_0_0_0; // @[Top.scala 140:12]
  assign n56_I0_15_0_0_1 = n43_O_15_0_0_1; // @[Top.scala 140:12]
  assign n56_I1_0_0_0 = n2_O_0_0_0; // @[Top.scala 141:12]
  assign n56_I1_1_0_0 = n2_O_1_0_0; // @[Top.scala 141:12]
  assign n56_I1_2_0_0 = n2_O_2_0_0; // @[Top.scala 141:12]
  assign n56_I1_3_0_0 = n2_O_3_0_0; // @[Top.scala 141:12]
  assign n56_I1_4_0_0 = n2_O_4_0_0; // @[Top.scala 141:12]
  assign n56_I1_5_0_0 = n2_O_5_0_0; // @[Top.scala 141:12]
  assign n56_I1_6_0_0 = n2_O_6_0_0; // @[Top.scala 141:12]
  assign n56_I1_7_0_0 = n2_O_7_0_0; // @[Top.scala 141:12]
  assign n56_I1_8_0_0 = n2_O_8_0_0; // @[Top.scala 141:12]
  assign n56_I1_9_0_0 = n2_O_9_0_0; // @[Top.scala 141:12]
  assign n56_I1_10_0_0 = n2_O_10_0_0; // @[Top.scala 141:12]
  assign n56_I1_11_0_0 = n2_O_11_0_0; // @[Top.scala 141:12]
  assign n56_I1_12_0_0 = n2_O_12_0_0; // @[Top.scala 141:12]
  assign n56_I1_13_0_0 = n2_O_13_0_0; // @[Top.scala 141:12]
  assign n56_I1_14_0_0 = n2_O_14_0_0; // @[Top.scala 141:12]
  assign n56_I1_15_0_0 = n2_O_15_0_0; // @[Top.scala 141:12]
  assign n77_valid_up = n56_valid_down; // @[Top.scala 145:18]
  assign n77_I_0_0_0_0 = n56_O_0_0_0_0; // @[Top.scala 144:11]
  assign n77_I_0_0_0_1 = n56_O_0_0_0_1; // @[Top.scala 144:11]
  assign n77_I_0_0_0_2 = n56_O_0_0_0_2; // @[Top.scala 144:11]
  assign n77_I_1_0_0_0 = n56_O_1_0_0_0; // @[Top.scala 144:11]
  assign n77_I_1_0_0_1 = n56_O_1_0_0_1; // @[Top.scala 144:11]
  assign n77_I_1_0_0_2 = n56_O_1_0_0_2; // @[Top.scala 144:11]
  assign n77_I_2_0_0_0 = n56_O_2_0_0_0; // @[Top.scala 144:11]
  assign n77_I_2_0_0_1 = n56_O_2_0_0_1; // @[Top.scala 144:11]
  assign n77_I_2_0_0_2 = n56_O_2_0_0_2; // @[Top.scala 144:11]
  assign n77_I_3_0_0_0 = n56_O_3_0_0_0; // @[Top.scala 144:11]
  assign n77_I_3_0_0_1 = n56_O_3_0_0_1; // @[Top.scala 144:11]
  assign n77_I_3_0_0_2 = n56_O_3_0_0_2; // @[Top.scala 144:11]
  assign n77_I_4_0_0_0 = n56_O_4_0_0_0; // @[Top.scala 144:11]
  assign n77_I_4_0_0_1 = n56_O_4_0_0_1; // @[Top.scala 144:11]
  assign n77_I_4_0_0_2 = n56_O_4_0_0_2; // @[Top.scala 144:11]
  assign n77_I_5_0_0_0 = n56_O_5_0_0_0; // @[Top.scala 144:11]
  assign n77_I_5_0_0_1 = n56_O_5_0_0_1; // @[Top.scala 144:11]
  assign n77_I_5_0_0_2 = n56_O_5_0_0_2; // @[Top.scala 144:11]
  assign n77_I_6_0_0_0 = n56_O_6_0_0_0; // @[Top.scala 144:11]
  assign n77_I_6_0_0_1 = n56_O_6_0_0_1; // @[Top.scala 144:11]
  assign n77_I_6_0_0_2 = n56_O_6_0_0_2; // @[Top.scala 144:11]
  assign n77_I_7_0_0_0 = n56_O_7_0_0_0; // @[Top.scala 144:11]
  assign n77_I_7_0_0_1 = n56_O_7_0_0_1; // @[Top.scala 144:11]
  assign n77_I_7_0_0_2 = n56_O_7_0_0_2; // @[Top.scala 144:11]
  assign n77_I_8_0_0_0 = n56_O_8_0_0_0; // @[Top.scala 144:11]
  assign n77_I_8_0_0_1 = n56_O_8_0_0_1; // @[Top.scala 144:11]
  assign n77_I_8_0_0_2 = n56_O_8_0_0_2; // @[Top.scala 144:11]
  assign n77_I_9_0_0_0 = n56_O_9_0_0_0; // @[Top.scala 144:11]
  assign n77_I_9_0_0_1 = n56_O_9_0_0_1; // @[Top.scala 144:11]
  assign n77_I_9_0_0_2 = n56_O_9_0_0_2; // @[Top.scala 144:11]
  assign n77_I_10_0_0_0 = n56_O_10_0_0_0; // @[Top.scala 144:11]
  assign n77_I_10_0_0_1 = n56_O_10_0_0_1; // @[Top.scala 144:11]
  assign n77_I_10_0_0_2 = n56_O_10_0_0_2; // @[Top.scala 144:11]
  assign n77_I_11_0_0_0 = n56_O_11_0_0_0; // @[Top.scala 144:11]
  assign n77_I_11_0_0_1 = n56_O_11_0_0_1; // @[Top.scala 144:11]
  assign n77_I_11_0_0_2 = n56_O_11_0_0_2; // @[Top.scala 144:11]
  assign n77_I_12_0_0_0 = n56_O_12_0_0_0; // @[Top.scala 144:11]
  assign n77_I_12_0_0_1 = n56_O_12_0_0_1; // @[Top.scala 144:11]
  assign n77_I_12_0_0_2 = n56_O_12_0_0_2; // @[Top.scala 144:11]
  assign n77_I_13_0_0_0 = n56_O_13_0_0_0; // @[Top.scala 144:11]
  assign n77_I_13_0_0_1 = n56_O_13_0_0_1; // @[Top.scala 144:11]
  assign n77_I_13_0_0_2 = n56_O_13_0_0_2; // @[Top.scala 144:11]
  assign n77_I_14_0_0_0 = n56_O_14_0_0_0; // @[Top.scala 144:11]
  assign n77_I_14_0_0_1 = n56_O_14_0_0_1; // @[Top.scala 144:11]
  assign n77_I_14_0_0_2 = n56_O_14_0_0_2; // @[Top.scala 144:11]
  assign n77_I_15_0_0_0 = n56_O_15_0_0_0; // @[Top.scala 144:11]
  assign n77_I_15_0_0_1 = n56_O_15_0_0_1; // @[Top.scala 144:11]
  assign n77_I_15_0_0_2 = n56_O_15_0_0_2; // @[Top.scala 144:11]
  assign n78_valid_up = n40_valid_down & n77_valid_down; // @[Top.scala 149:18]
  assign n78_I0_0_0_0 = n40_O_0_0_0; // @[Top.scala 147:12]
  assign n78_I0_0_0_1 = n40_O_0_0_1; // @[Top.scala 147:12]
  assign n78_I0_0_0_2 = n40_O_0_0_2; // @[Top.scala 147:12]
  assign n78_I0_1_0_0 = n40_O_1_0_0; // @[Top.scala 147:12]
  assign n78_I0_1_0_1 = n40_O_1_0_1; // @[Top.scala 147:12]
  assign n78_I0_1_0_2 = n40_O_1_0_2; // @[Top.scala 147:12]
  assign n78_I0_2_0_0 = n40_O_2_0_0; // @[Top.scala 147:12]
  assign n78_I0_2_0_1 = n40_O_2_0_1; // @[Top.scala 147:12]
  assign n78_I0_2_0_2 = n40_O_2_0_2; // @[Top.scala 147:12]
  assign n78_I0_3_0_0 = n40_O_3_0_0; // @[Top.scala 147:12]
  assign n78_I0_3_0_1 = n40_O_3_0_1; // @[Top.scala 147:12]
  assign n78_I0_3_0_2 = n40_O_3_0_2; // @[Top.scala 147:12]
  assign n78_I0_4_0_0 = n40_O_4_0_0; // @[Top.scala 147:12]
  assign n78_I0_4_0_1 = n40_O_4_0_1; // @[Top.scala 147:12]
  assign n78_I0_4_0_2 = n40_O_4_0_2; // @[Top.scala 147:12]
  assign n78_I0_5_0_0 = n40_O_5_0_0; // @[Top.scala 147:12]
  assign n78_I0_5_0_1 = n40_O_5_0_1; // @[Top.scala 147:12]
  assign n78_I0_5_0_2 = n40_O_5_0_2; // @[Top.scala 147:12]
  assign n78_I0_6_0_0 = n40_O_6_0_0; // @[Top.scala 147:12]
  assign n78_I0_6_0_1 = n40_O_6_0_1; // @[Top.scala 147:12]
  assign n78_I0_6_0_2 = n40_O_6_0_2; // @[Top.scala 147:12]
  assign n78_I0_7_0_0 = n40_O_7_0_0; // @[Top.scala 147:12]
  assign n78_I0_7_0_1 = n40_O_7_0_1; // @[Top.scala 147:12]
  assign n78_I0_7_0_2 = n40_O_7_0_2; // @[Top.scala 147:12]
  assign n78_I0_8_0_0 = n40_O_8_0_0; // @[Top.scala 147:12]
  assign n78_I0_8_0_1 = n40_O_8_0_1; // @[Top.scala 147:12]
  assign n78_I0_8_0_2 = n40_O_8_0_2; // @[Top.scala 147:12]
  assign n78_I0_9_0_0 = n40_O_9_0_0; // @[Top.scala 147:12]
  assign n78_I0_9_0_1 = n40_O_9_0_1; // @[Top.scala 147:12]
  assign n78_I0_9_0_2 = n40_O_9_0_2; // @[Top.scala 147:12]
  assign n78_I0_10_0_0 = n40_O_10_0_0; // @[Top.scala 147:12]
  assign n78_I0_10_0_1 = n40_O_10_0_1; // @[Top.scala 147:12]
  assign n78_I0_10_0_2 = n40_O_10_0_2; // @[Top.scala 147:12]
  assign n78_I0_11_0_0 = n40_O_11_0_0; // @[Top.scala 147:12]
  assign n78_I0_11_0_1 = n40_O_11_0_1; // @[Top.scala 147:12]
  assign n78_I0_11_0_2 = n40_O_11_0_2; // @[Top.scala 147:12]
  assign n78_I0_12_0_0 = n40_O_12_0_0; // @[Top.scala 147:12]
  assign n78_I0_12_0_1 = n40_O_12_0_1; // @[Top.scala 147:12]
  assign n78_I0_12_0_2 = n40_O_12_0_2; // @[Top.scala 147:12]
  assign n78_I0_13_0_0 = n40_O_13_0_0; // @[Top.scala 147:12]
  assign n78_I0_13_0_1 = n40_O_13_0_1; // @[Top.scala 147:12]
  assign n78_I0_13_0_2 = n40_O_13_0_2; // @[Top.scala 147:12]
  assign n78_I0_14_0_0 = n40_O_14_0_0; // @[Top.scala 147:12]
  assign n78_I0_14_0_1 = n40_O_14_0_1; // @[Top.scala 147:12]
  assign n78_I0_14_0_2 = n40_O_14_0_2; // @[Top.scala 147:12]
  assign n78_I0_15_0_0 = n40_O_15_0_0; // @[Top.scala 147:12]
  assign n78_I0_15_0_1 = n40_O_15_0_1; // @[Top.scala 147:12]
  assign n78_I0_15_0_2 = n40_O_15_0_2; // @[Top.scala 147:12]
  assign n78_I1_0_0_0 = n77_O_0_0_0; // @[Top.scala 148:12]
  assign n78_I1_0_0_1 = n77_O_0_0_1; // @[Top.scala 148:12]
  assign n78_I1_0_0_2 = n77_O_0_0_2; // @[Top.scala 148:12]
  assign n78_I1_1_0_0 = n77_O_1_0_0; // @[Top.scala 148:12]
  assign n78_I1_1_0_1 = n77_O_1_0_1; // @[Top.scala 148:12]
  assign n78_I1_1_0_2 = n77_O_1_0_2; // @[Top.scala 148:12]
  assign n78_I1_2_0_0 = n77_O_2_0_0; // @[Top.scala 148:12]
  assign n78_I1_2_0_1 = n77_O_2_0_1; // @[Top.scala 148:12]
  assign n78_I1_2_0_2 = n77_O_2_0_2; // @[Top.scala 148:12]
  assign n78_I1_3_0_0 = n77_O_3_0_0; // @[Top.scala 148:12]
  assign n78_I1_3_0_1 = n77_O_3_0_1; // @[Top.scala 148:12]
  assign n78_I1_3_0_2 = n77_O_3_0_2; // @[Top.scala 148:12]
  assign n78_I1_4_0_0 = n77_O_4_0_0; // @[Top.scala 148:12]
  assign n78_I1_4_0_1 = n77_O_4_0_1; // @[Top.scala 148:12]
  assign n78_I1_4_0_2 = n77_O_4_0_2; // @[Top.scala 148:12]
  assign n78_I1_5_0_0 = n77_O_5_0_0; // @[Top.scala 148:12]
  assign n78_I1_5_0_1 = n77_O_5_0_1; // @[Top.scala 148:12]
  assign n78_I1_5_0_2 = n77_O_5_0_2; // @[Top.scala 148:12]
  assign n78_I1_6_0_0 = n77_O_6_0_0; // @[Top.scala 148:12]
  assign n78_I1_6_0_1 = n77_O_6_0_1; // @[Top.scala 148:12]
  assign n78_I1_6_0_2 = n77_O_6_0_2; // @[Top.scala 148:12]
  assign n78_I1_7_0_0 = n77_O_7_0_0; // @[Top.scala 148:12]
  assign n78_I1_7_0_1 = n77_O_7_0_1; // @[Top.scala 148:12]
  assign n78_I1_7_0_2 = n77_O_7_0_2; // @[Top.scala 148:12]
  assign n78_I1_8_0_0 = n77_O_8_0_0; // @[Top.scala 148:12]
  assign n78_I1_8_0_1 = n77_O_8_0_1; // @[Top.scala 148:12]
  assign n78_I1_8_0_2 = n77_O_8_0_2; // @[Top.scala 148:12]
  assign n78_I1_9_0_0 = n77_O_9_0_0; // @[Top.scala 148:12]
  assign n78_I1_9_0_1 = n77_O_9_0_1; // @[Top.scala 148:12]
  assign n78_I1_9_0_2 = n77_O_9_0_2; // @[Top.scala 148:12]
  assign n78_I1_10_0_0 = n77_O_10_0_0; // @[Top.scala 148:12]
  assign n78_I1_10_0_1 = n77_O_10_0_1; // @[Top.scala 148:12]
  assign n78_I1_10_0_2 = n77_O_10_0_2; // @[Top.scala 148:12]
  assign n78_I1_11_0_0 = n77_O_11_0_0; // @[Top.scala 148:12]
  assign n78_I1_11_0_1 = n77_O_11_0_1; // @[Top.scala 148:12]
  assign n78_I1_11_0_2 = n77_O_11_0_2; // @[Top.scala 148:12]
  assign n78_I1_12_0_0 = n77_O_12_0_0; // @[Top.scala 148:12]
  assign n78_I1_12_0_1 = n77_O_12_0_1; // @[Top.scala 148:12]
  assign n78_I1_12_0_2 = n77_O_12_0_2; // @[Top.scala 148:12]
  assign n78_I1_13_0_0 = n77_O_13_0_0; // @[Top.scala 148:12]
  assign n78_I1_13_0_1 = n77_O_13_0_1; // @[Top.scala 148:12]
  assign n78_I1_13_0_2 = n77_O_13_0_2; // @[Top.scala 148:12]
  assign n78_I1_14_0_0 = n77_O_14_0_0; // @[Top.scala 148:12]
  assign n78_I1_14_0_1 = n77_O_14_0_1; // @[Top.scala 148:12]
  assign n78_I1_14_0_2 = n77_O_14_0_2; // @[Top.scala 148:12]
  assign n78_I1_15_0_0 = n77_O_15_0_0; // @[Top.scala 148:12]
  assign n78_I1_15_0_1 = n77_O_15_0_1; // @[Top.scala 148:12]
  assign n78_I1_15_0_2 = n77_O_15_0_2; // @[Top.scala 148:12]
  assign n88_clock = clock;
  assign n88_valid_up = n1_valid_down; // @[Top.scala 152:18]
  assign n88_I_0_0_0 = n1_O_0_0_0; // @[Top.scala 151:11]
  assign n88_I_1_0_0 = n1_O_1_0_0; // @[Top.scala 151:11]
  assign n88_I_2_0_0 = n1_O_2_0_0; // @[Top.scala 151:11]
  assign n88_I_3_0_0 = n1_O_3_0_0; // @[Top.scala 151:11]
  assign n88_I_4_0_0 = n1_O_4_0_0; // @[Top.scala 151:11]
  assign n88_I_5_0_0 = n1_O_5_0_0; // @[Top.scala 151:11]
  assign n88_I_6_0_0 = n1_O_6_0_0; // @[Top.scala 151:11]
  assign n88_I_7_0_0 = n1_O_7_0_0; // @[Top.scala 151:11]
  assign n88_I_8_0_0 = n1_O_8_0_0; // @[Top.scala 151:11]
  assign n88_I_9_0_0 = n1_O_9_0_0; // @[Top.scala 151:11]
  assign n88_I_10_0_0 = n1_O_10_0_0; // @[Top.scala 151:11]
  assign n88_I_11_0_0 = n1_O_11_0_0; // @[Top.scala 151:11]
  assign n88_I_12_0_0 = n1_O_12_0_0; // @[Top.scala 151:11]
  assign n88_I_13_0_0 = n1_O_13_0_0; // @[Top.scala 151:11]
  assign n88_I_14_0_0 = n1_O_14_0_0; // @[Top.scala 151:11]
  assign n88_I_15_0_0 = n1_O_15_0_0; // @[Top.scala 151:11]
  assign n89_clock = clock;
  assign n89_valid_up = n88_valid_down; // @[Top.scala 155:18]
  assign n89_I_0_0_0 = n88_O_0_0_0; // @[Top.scala 154:11]
  assign n89_I_1_0_0 = n88_O_1_0_0; // @[Top.scala 154:11]
  assign n89_I_2_0_0 = n88_O_2_0_0; // @[Top.scala 154:11]
  assign n89_I_3_0_0 = n88_O_3_0_0; // @[Top.scala 154:11]
  assign n89_I_4_0_0 = n88_O_4_0_0; // @[Top.scala 154:11]
  assign n89_I_5_0_0 = n88_O_5_0_0; // @[Top.scala 154:11]
  assign n89_I_6_0_0 = n88_O_6_0_0; // @[Top.scala 154:11]
  assign n89_I_7_0_0 = n88_O_7_0_0; // @[Top.scala 154:11]
  assign n89_I_8_0_0 = n88_O_8_0_0; // @[Top.scala 154:11]
  assign n89_I_9_0_0 = n88_O_9_0_0; // @[Top.scala 154:11]
  assign n89_I_10_0_0 = n88_O_10_0_0; // @[Top.scala 154:11]
  assign n89_I_11_0_0 = n88_O_11_0_0; // @[Top.scala 154:11]
  assign n89_I_12_0_0 = n88_O_12_0_0; // @[Top.scala 154:11]
  assign n89_I_13_0_0 = n88_O_13_0_0; // @[Top.scala 154:11]
  assign n89_I_14_0_0 = n88_O_14_0_0; // @[Top.scala 154:11]
  assign n89_I_15_0_0 = n88_O_15_0_0; // @[Top.scala 154:11]
  assign n90_valid_up = n89_valid_down & n88_valid_down; // @[Top.scala 159:18]
  assign n90_I0_0_0_0 = n89_O_0_0_0; // @[Top.scala 157:12]
  assign n90_I0_1_0_0 = n89_O_1_0_0; // @[Top.scala 157:12]
  assign n90_I0_2_0_0 = n89_O_2_0_0; // @[Top.scala 157:12]
  assign n90_I0_3_0_0 = n89_O_3_0_0; // @[Top.scala 157:12]
  assign n90_I0_4_0_0 = n89_O_4_0_0; // @[Top.scala 157:12]
  assign n90_I0_5_0_0 = n89_O_5_0_0; // @[Top.scala 157:12]
  assign n90_I0_6_0_0 = n89_O_6_0_0; // @[Top.scala 157:12]
  assign n90_I0_7_0_0 = n89_O_7_0_0; // @[Top.scala 157:12]
  assign n90_I0_8_0_0 = n89_O_8_0_0; // @[Top.scala 157:12]
  assign n90_I0_9_0_0 = n89_O_9_0_0; // @[Top.scala 157:12]
  assign n90_I0_10_0_0 = n89_O_10_0_0; // @[Top.scala 157:12]
  assign n90_I0_11_0_0 = n89_O_11_0_0; // @[Top.scala 157:12]
  assign n90_I0_12_0_0 = n89_O_12_0_0; // @[Top.scala 157:12]
  assign n90_I0_13_0_0 = n89_O_13_0_0; // @[Top.scala 157:12]
  assign n90_I0_14_0_0 = n89_O_14_0_0; // @[Top.scala 157:12]
  assign n90_I0_15_0_0 = n89_O_15_0_0; // @[Top.scala 157:12]
  assign n90_I1_0_0_0 = n88_O_0_0_0; // @[Top.scala 158:12]
  assign n90_I1_1_0_0 = n88_O_1_0_0; // @[Top.scala 158:12]
  assign n90_I1_2_0_0 = n88_O_2_0_0; // @[Top.scala 158:12]
  assign n90_I1_3_0_0 = n88_O_3_0_0; // @[Top.scala 158:12]
  assign n90_I1_4_0_0 = n88_O_4_0_0; // @[Top.scala 158:12]
  assign n90_I1_5_0_0 = n88_O_5_0_0; // @[Top.scala 158:12]
  assign n90_I1_6_0_0 = n88_O_6_0_0; // @[Top.scala 158:12]
  assign n90_I1_7_0_0 = n88_O_7_0_0; // @[Top.scala 158:12]
  assign n90_I1_8_0_0 = n88_O_8_0_0; // @[Top.scala 158:12]
  assign n90_I1_9_0_0 = n88_O_9_0_0; // @[Top.scala 158:12]
  assign n90_I1_10_0_0 = n88_O_10_0_0; // @[Top.scala 158:12]
  assign n90_I1_11_0_0 = n88_O_11_0_0; // @[Top.scala 158:12]
  assign n90_I1_12_0_0 = n88_O_12_0_0; // @[Top.scala 158:12]
  assign n90_I1_13_0_0 = n88_O_13_0_0; // @[Top.scala 158:12]
  assign n90_I1_14_0_0 = n88_O_14_0_0; // @[Top.scala 158:12]
  assign n90_I1_15_0_0 = n88_O_15_0_0; // @[Top.scala 158:12]
  assign n103_valid_up = n90_valid_down & n1_valid_down; // @[Top.scala 163:19]
  assign n103_I0_0_0_0_0 = n90_O_0_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_0_0_0_1 = n90_O_0_0_0_1; // @[Top.scala 161:13]
  assign n103_I0_1_0_0_0 = n90_O_1_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_1_0_0_1 = n90_O_1_0_0_1; // @[Top.scala 161:13]
  assign n103_I0_2_0_0_0 = n90_O_2_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_2_0_0_1 = n90_O_2_0_0_1; // @[Top.scala 161:13]
  assign n103_I0_3_0_0_0 = n90_O_3_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_3_0_0_1 = n90_O_3_0_0_1; // @[Top.scala 161:13]
  assign n103_I0_4_0_0_0 = n90_O_4_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_4_0_0_1 = n90_O_4_0_0_1; // @[Top.scala 161:13]
  assign n103_I0_5_0_0_0 = n90_O_5_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_5_0_0_1 = n90_O_5_0_0_1; // @[Top.scala 161:13]
  assign n103_I0_6_0_0_0 = n90_O_6_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_6_0_0_1 = n90_O_6_0_0_1; // @[Top.scala 161:13]
  assign n103_I0_7_0_0_0 = n90_O_7_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_7_0_0_1 = n90_O_7_0_0_1; // @[Top.scala 161:13]
  assign n103_I0_8_0_0_0 = n90_O_8_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_8_0_0_1 = n90_O_8_0_0_1; // @[Top.scala 161:13]
  assign n103_I0_9_0_0_0 = n90_O_9_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_9_0_0_1 = n90_O_9_0_0_1; // @[Top.scala 161:13]
  assign n103_I0_10_0_0_0 = n90_O_10_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_10_0_0_1 = n90_O_10_0_0_1; // @[Top.scala 161:13]
  assign n103_I0_11_0_0_0 = n90_O_11_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_11_0_0_1 = n90_O_11_0_0_1; // @[Top.scala 161:13]
  assign n103_I0_12_0_0_0 = n90_O_12_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_12_0_0_1 = n90_O_12_0_0_1; // @[Top.scala 161:13]
  assign n103_I0_13_0_0_0 = n90_O_13_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_13_0_0_1 = n90_O_13_0_0_1; // @[Top.scala 161:13]
  assign n103_I0_14_0_0_0 = n90_O_14_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_14_0_0_1 = n90_O_14_0_0_1; // @[Top.scala 161:13]
  assign n103_I0_15_0_0_0 = n90_O_15_0_0_0; // @[Top.scala 161:13]
  assign n103_I0_15_0_0_1 = n90_O_15_0_0_1; // @[Top.scala 161:13]
  assign n103_I1_0_0_0 = n1_O_0_0_0; // @[Top.scala 162:13]
  assign n103_I1_1_0_0 = n1_O_1_0_0; // @[Top.scala 162:13]
  assign n103_I1_2_0_0 = n1_O_2_0_0; // @[Top.scala 162:13]
  assign n103_I1_3_0_0 = n1_O_3_0_0; // @[Top.scala 162:13]
  assign n103_I1_4_0_0 = n1_O_4_0_0; // @[Top.scala 162:13]
  assign n103_I1_5_0_0 = n1_O_5_0_0; // @[Top.scala 162:13]
  assign n103_I1_6_0_0 = n1_O_6_0_0; // @[Top.scala 162:13]
  assign n103_I1_7_0_0 = n1_O_7_0_0; // @[Top.scala 162:13]
  assign n103_I1_8_0_0 = n1_O_8_0_0; // @[Top.scala 162:13]
  assign n103_I1_9_0_0 = n1_O_9_0_0; // @[Top.scala 162:13]
  assign n103_I1_10_0_0 = n1_O_10_0_0; // @[Top.scala 162:13]
  assign n103_I1_11_0_0 = n1_O_11_0_0; // @[Top.scala 162:13]
  assign n103_I1_12_0_0 = n1_O_12_0_0; // @[Top.scala 162:13]
  assign n103_I1_13_0_0 = n1_O_13_0_0; // @[Top.scala 162:13]
  assign n103_I1_14_0_0 = n1_O_14_0_0; // @[Top.scala 162:13]
  assign n103_I1_15_0_0 = n1_O_15_0_0; // @[Top.scala 162:13]
  assign n124_valid_up = n103_valid_down; // @[Top.scala 166:19]
  assign n124_I_0_0_0_0 = n103_O_0_0_0_0; // @[Top.scala 165:12]
  assign n124_I_0_0_0_1 = n103_O_0_0_0_1; // @[Top.scala 165:12]
  assign n124_I_0_0_0_2 = n103_O_0_0_0_2; // @[Top.scala 165:12]
  assign n124_I_1_0_0_0 = n103_O_1_0_0_0; // @[Top.scala 165:12]
  assign n124_I_1_0_0_1 = n103_O_1_0_0_1; // @[Top.scala 165:12]
  assign n124_I_1_0_0_2 = n103_O_1_0_0_2; // @[Top.scala 165:12]
  assign n124_I_2_0_0_0 = n103_O_2_0_0_0; // @[Top.scala 165:12]
  assign n124_I_2_0_0_1 = n103_O_2_0_0_1; // @[Top.scala 165:12]
  assign n124_I_2_0_0_2 = n103_O_2_0_0_2; // @[Top.scala 165:12]
  assign n124_I_3_0_0_0 = n103_O_3_0_0_0; // @[Top.scala 165:12]
  assign n124_I_3_0_0_1 = n103_O_3_0_0_1; // @[Top.scala 165:12]
  assign n124_I_3_0_0_2 = n103_O_3_0_0_2; // @[Top.scala 165:12]
  assign n124_I_4_0_0_0 = n103_O_4_0_0_0; // @[Top.scala 165:12]
  assign n124_I_4_0_0_1 = n103_O_4_0_0_1; // @[Top.scala 165:12]
  assign n124_I_4_0_0_2 = n103_O_4_0_0_2; // @[Top.scala 165:12]
  assign n124_I_5_0_0_0 = n103_O_5_0_0_0; // @[Top.scala 165:12]
  assign n124_I_5_0_0_1 = n103_O_5_0_0_1; // @[Top.scala 165:12]
  assign n124_I_5_0_0_2 = n103_O_5_0_0_2; // @[Top.scala 165:12]
  assign n124_I_6_0_0_0 = n103_O_6_0_0_0; // @[Top.scala 165:12]
  assign n124_I_6_0_0_1 = n103_O_6_0_0_1; // @[Top.scala 165:12]
  assign n124_I_6_0_0_2 = n103_O_6_0_0_2; // @[Top.scala 165:12]
  assign n124_I_7_0_0_0 = n103_O_7_0_0_0; // @[Top.scala 165:12]
  assign n124_I_7_0_0_1 = n103_O_7_0_0_1; // @[Top.scala 165:12]
  assign n124_I_7_0_0_2 = n103_O_7_0_0_2; // @[Top.scala 165:12]
  assign n124_I_8_0_0_0 = n103_O_8_0_0_0; // @[Top.scala 165:12]
  assign n124_I_8_0_0_1 = n103_O_8_0_0_1; // @[Top.scala 165:12]
  assign n124_I_8_0_0_2 = n103_O_8_0_0_2; // @[Top.scala 165:12]
  assign n124_I_9_0_0_0 = n103_O_9_0_0_0; // @[Top.scala 165:12]
  assign n124_I_9_0_0_1 = n103_O_9_0_0_1; // @[Top.scala 165:12]
  assign n124_I_9_0_0_2 = n103_O_9_0_0_2; // @[Top.scala 165:12]
  assign n124_I_10_0_0_0 = n103_O_10_0_0_0; // @[Top.scala 165:12]
  assign n124_I_10_0_0_1 = n103_O_10_0_0_1; // @[Top.scala 165:12]
  assign n124_I_10_0_0_2 = n103_O_10_0_0_2; // @[Top.scala 165:12]
  assign n124_I_11_0_0_0 = n103_O_11_0_0_0; // @[Top.scala 165:12]
  assign n124_I_11_0_0_1 = n103_O_11_0_0_1; // @[Top.scala 165:12]
  assign n124_I_11_0_0_2 = n103_O_11_0_0_2; // @[Top.scala 165:12]
  assign n124_I_12_0_0_0 = n103_O_12_0_0_0; // @[Top.scala 165:12]
  assign n124_I_12_0_0_1 = n103_O_12_0_0_1; // @[Top.scala 165:12]
  assign n124_I_12_0_0_2 = n103_O_12_0_0_2; // @[Top.scala 165:12]
  assign n124_I_13_0_0_0 = n103_O_13_0_0_0; // @[Top.scala 165:12]
  assign n124_I_13_0_0_1 = n103_O_13_0_0_1; // @[Top.scala 165:12]
  assign n124_I_13_0_0_2 = n103_O_13_0_0_2; // @[Top.scala 165:12]
  assign n124_I_14_0_0_0 = n103_O_14_0_0_0; // @[Top.scala 165:12]
  assign n124_I_14_0_0_1 = n103_O_14_0_0_1; // @[Top.scala 165:12]
  assign n124_I_14_0_0_2 = n103_O_14_0_0_2; // @[Top.scala 165:12]
  assign n124_I_15_0_0_0 = n103_O_15_0_0_0; // @[Top.scala 165:12]
  assign n124_I_15_0_0_1 = n103_O_15_0_0_1; // @[Top.scala 165:12]
  assign n124_I_15_0_0_2 = n103_O_15_0_0_2; // @[Top.scala 165:12]
  assign n125_valid_up = n78_valid_down & n124_valid_down; // @[Top.scala 170:19]
  assign n125_I0_0_0_0_0 = n78_O_0_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_0_0_0_1 = n78_O_0_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_0_0_0_2 = n78_O_0_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_0_0_1_0 = n78_O_0_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_0_0_1_1 = n78_O_0_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_0_0_1_2 = n78_O_0_0_1_2; // @[Top.scala 168:13]
  assign n125_I0_1_0_0_0 = n78_O_1_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_1_0_0_1 = n78_O_1_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_1_0_0_2 = n78_O_1_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_1_0_1_0 = n78_O_1_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_1_0_1_1 = n78_O_1_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_1_0_1_2 = n78_O_1_0_1_2; // @[Top.scala 168:13]
  assign n125_I0_2_0_0_0 = n78_O_2_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_2_0_0_1 = n78_O_2_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_2_0_0_2 = n78_O_2_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_2_0_1_0 = n78_O_2_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_2_0_1_1 = n78_O_2_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_2_0_1_2 = n78_O_2_0_1_2; // @[Top.scala 168:13]
  assign n125_I0_3_0_0_0 = n78_O_3_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_3_0_0_1 = n78_O_3_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_3_0_0_2 = n78_O_3_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_3_0_1_0 = n78_O_3_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_3_0_1_1 = n78_O_3_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_3_0_1_2 = n78_O_3_0_1_2; // @[Top.scala 168:13]
  assign n125_I0_4_0_0_0 = n78_O_4_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_4_0_0_1 = n78_O_4_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_4_0_0_2 = n78_O_4_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_4_0_1_0 = n78_O_4_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_4_0_1_1 = n78_O_4_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_4_0_1_2 = n78_O_4_0_1_2; // @[Top.scala 168:13]
  assign n125_I0_5_0_0_0 = n78_O_5_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_5_0_0_1 = n78_O_5_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_5_0_0_2 = n78_O_5_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_5_0_1_0 = n78_O_5_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_5_0_1_1 = n78_O_5_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_5_0_1_2 = n78_O_5_0_1_2; // @[Top.scala 168:13]
  assign n125_I0_6_0_0_0 = n78_O_6_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_6_0_0_1 = n78_O_6_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_6_0_0_2 = n78_O_6_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_6_0_1_0 = n78_O_6_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_6_0_1_1 = n78_O_6_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_6_0_1_2 = n78_O_6_0_1_2; // @[Top.scala 168:13]
  assign n125_I0_7_0_0_0 = n78_O_7_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_7_0_0_1 = n78_O_7_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_7_0_0_2 = n78_O_7_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_7_0_1_0 = n78_O_7_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_7_0_1_1 = n78_O_7_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_7_0_1_2 = n78_O_7_0_1_2; // @[Top.scala 168:13]
  assign n125_I0_8_0_0_0 = n78_O_8_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_8_0_0_1 = n78_O_8_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_8_0_0_2 = n78_O_8_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_8_0_1_0 = n78_O_8_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_8_0_1_1 = n78_O_8_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_8_0_1_2 = n78_O_8_0_1_2; // @[Top.scala 168:13]
  assign n125_I0_9_0_0_0 = n78_O_9_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_9_0_0_1 = n78_O_9_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_9_0_0_2 = n78_O_9_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_9_0_1_0 = n78_O_9_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_9_0_1_1 = n78_O_9_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_9_0_1_2 = n78_O_9_0_1_2; // @[Top.scala 168:13]
  assign n125_I0_10_0_0_0 = n78_O_10_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_10_0_0_1 = n78_O_10_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_10_0_0_2 = n78_O_10_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_10_0_1_0 = n78_O_10_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_10_0_1_1 = n78_O_10_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_10_0_1_2 = n78_O_10_0_1_2; // @[Top.scala 168:13]
  assign n125_I0_11_0_0_0 = n78_O_11_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_11_0_0_1 = n78_O_11_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_11_0_0_2 = n78_O_11_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_11_0_1_0 = n78_O_11_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_11_0_1_1 = n78_O_11_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_11_0_1_2 = n78_O_11_0_1_2; // @[Top.scala 168:13]
  assign n125_I0_12_0_0_0 = n78_O_12_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_12_0_0_1 = n78_O_12_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_12_0_0_2 = n78_O_12_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_12_0_1_0 = n78_O_12_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_12_0_1_1 = n78_O_12_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_12_0_1_2 = n78_O_12_0_1_2; // @[Top.scala 168:13]
  assign n125_I0_13_0_0_0 = n78_O_13_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_13_0_0_1 = n78_O_13_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_13_0_0_2 = n78_O_13_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_13_0_1_0 = n78_O_13_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_13_0_1_1 = n78_O_13_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_13_0_1_2 = n78_O_13_0_1_2; // @[Top.scala 168:13]
  assign n125_I0_14_0_0_0 = n78_O_14_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_14_0_0_1 = n78_O_14_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_14_0_0_2 = n78_O_14_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_14_0_1_0 = n78_O_14_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_14_0_1_1 = n78_O_14_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_14_0_1_2 = n78_O_14_0_1_2; // @[Top.scala 168:13]
  assign n125_I0_15_0_0_0 = n78_O_15_0_0_0; // @[Top.scala 168:13]
  assign n125_I0_15_0_0_1 = n78_O_15_0_0_1; // @[Top.scala 168:13]
  assign n125_I0_15_0_0_2 = n78_O_15_0_0_2; // @[Top.scala 168:13]
  assign n125_I0_15_0_1_0 = n78_O_15_0_1_0; // @[Top.scala 168:13]
  assign n125_I0_15_0_1_1 = n78_O_15_0_1_1; // @[Top.scala 168:13]
  assign n125_I0_15_0_1_2 = n78_O_15_0_1_2; // @[Top.scala 168:13]
  assign n125_I1_0_0_0 = n124_O_0_0_0; // @[Top.scala 169:13]
  assign n125_I1_0_0_1 = n124_O_0_0_1; // @[Top.scala 169:13]
  assign n125_I1_0_0_2 = n124_O_0_0_2; // @[Top.scala 169:13]
  assign n125_I1_1_0_0 = n124_O_1_0_0; // @[Top.scala 169:13]
  assign n125_I1_1_0_1 = n124_O_1_0_1; // @[Top.scala 169:13]
  assign n125_I1_1_0_2 = n124_O_1_0_2; // @[Top.scala 169:13]
  assign n125_I1_2_0_0 = n124_O_2_0_0; // @[Top.scala 169:13]
  assign n125_I1_2_0_1 = n124_O_2_0_1; // @[Top.scala 169:13]
  assign n125_I1_2_0_2 = n124_O_2_0_2; // @[Top.scala 169:13]
  assign n125_I1_3_0_0 = n124_O_3_0_0; // @[Top.scala 169:13]
  assign n125_I1_3_0_1 = n124_O_3_0_1; // @[Top.scala 169:13]
  assign n125_I1_3_0_2 = n124_O_3_0_2; // @[Top.scala 169:13]
  assign n125_I1_4_0_0 = n124_O_4_0_0; // @[Top.scala 169:13]
  assign n125_I1_4_0_1 = n124_O_4_0_1; // @[Top.scala 169:13]
  assign n125_I1_4_0_2 = n124_O_4_0_2; // @[Top.scala 169:13]
  assign n125_I1_5_0_0 = n124_O_5_0_0; // @[Top.scala 169:13]
  assign n125_I1_5_0_1 = n124_O_5_0_1; // @[Top.scala 169:13]
  assign n125_I1_5_0_2 = n124_O_5_0_2; // @[Top.scala 169:13]
  assign n125_I1_6_0_0 = n124_O_6_0_0; // @[Top.scala 169:13]
  assign n125_I1_6_0_1 = n124_O_6_0_1; // @[Top.scala 169:13]
  assign n125_I1_6_0_2 = n124_O_6_0_2; // @[Top.scala 169:13]
  assign n125_I1_7_0_0 = n124_O_7_0_0; // @[Top.scala 169:13]
  assign n125_I1_7_0_1 = n124_O_7_0_1; // @[Top.scala 169:13]
  assign n125_I1_7_0_2 = n124_O_7_0_2; // @[Top.scala 169:13]
  assign n125_I1_8_0_0 = n124_O_8_0_0; // @[Top.scala 169:13]
  assign n125_I1_8_0_1 = n124_O_8_0_1; // @[Top.scala 169:13]
  assign n125_I1_8_0_2 = n124_O_8_0_2; // @[Top.scala 169:13]
  assign n125_I1_9_0_0 = n124_O_9_0_0; // @[Top.scala 169:13]
  assign n125_I1_9_0_1 = n124_O_9_0_1; // @[Top.scala 169:13]
  assign n125_I1_9_0_2 = n124_O_9_0_2; // @[Top.scala 169:13]
  assign n125_I1_10_0_0 = n124_O_10_0_0; // @[Top.scala 169:13]
  assign n125_I1_10_0_1 = n124_O_10_0_1; // @[Top.scala 169:13]
  assign n125_I1_10_0_2 = n124_O_10_0_2; // @[Top.scala 169:13]
  assign n125_I1_11_0_0 = n124_O_11_0_0; // @[Top.scala 169:13]
  assign n125_I1_11_0_1 = n124_O_11_0_1; // @[Top.scala 169:13]
  assign n125_I1_11_0_2 = n124_O_11_0_2; // @[Top.scala 169:13]
  assign n125_I1_12_0_0 = n124_O_12_0_0; // @[Top.scala 169:13]
  assign n125_I1_12_0_1 = n124_O_12_0_1; // @[Top.scala 169:13]
  assign n125_I1_12_0_2 = n124_O_12_0_2; // @[Top.scala 169:13]
  assign n125_I1_13_0_0 = n124_O_13_0_0; // @[Top.scala 169:13]
  assign n125_I1_13_0_1 = n124_O_13_0_1; // @[Top.scala 169:13]
  assign n125_I1_13_0_2 = n124_O_13_0_2; // @[Top.scala 169:13]
  assign n125_I1_14_0_0 = n124_O_14_0_0; // @[Top.scala 169:13]
  assign n125_I1_14_0_1 = n124_O_14_0_1; // @[Top.scala 169:13]
  assign n125_I1_14_0_2 = n124_O_14_0_2; // @[Top.scala 169:13]
  assign n125_I1_15_0_0 = n124_O_15_0_0; // @[Top.scala 169:13]
  assign n125_I1_15_0_1 = n124_O_15_0_1; // @[Top.scala 169:13]
  assign n125_I1_15_0_2 = n124_O_15_0_2; // @[Top.scala 169:13]
  assign n141_valid_up = n125_valid_down; // @[Top.scala 173:19]
  assign n141_I_0_0_0_0 = n125_O_0_0_0_0; // @[Top.scala 172:12]
  assign n141_I_0_0_0_1 = n125_O_0_0_0_1; // @[Top.scala 172:12]
  assign n141_I_0_0_0_2 = n125_O_0_0_0_2; // @[Top.scala 172:12]
  assign n141_I_0_0_1_0 = n125_O_0_0_1_0; // @[Top.scala 172:12]
  assign n141_I_0_0_1_1 = n125_O_0_0_1_1; // @[Top.scala 172:12]
  assign n141_I_0_0_1_2 = n125_O_0_0_1_2; // @[Top.scala 172:12]
  assign n141_I_0_0_2_0 = n125_O_0_0_2_0; // @[Top.scala 172:12]
  assign n141_I_0_0_2_1 = n125_O_0_0_2_1; // @[Top.scala 172:12]
  assign n141_I_0_0_2_2 = n125_O_0_0_2_2; // @[Top.scala 172:12]
  assign n141_I_1_0_0_0 = n125_O_1_0_0_0; // @[Top.scala 172:12]
  assign n141_I_1_0_0_1 = n125_O_1_0_0_1; // @[Top.scala 172:12]
  assign n141_I_1_0_0_2 = n125_O_1_0_0_2; // @[Top.scala 172:12]
  assign n141_I_1_0_1_0 = n125_O_1_0_1_0; // @[Top.scala 172:12]
  assign n141_I_1_0_1_1 = n125_O_1_0_1_1; // @[Top.scala 172:12]
  assign n141_I_1_0_1_2 = n125_O_1_0_1_2; // @[Top.scala 172:12]
  assign n141_I_1_0_2_0 = n125_O_1_0_2_0; // @[Top.scala 172:12]
  assign n141_I_1_0_2_1 = n125_O_1_0_2_1; // @[Top.scala 172:12]
  assign n141_I_1_0_2_2 = n125_O_1_0_2_2; // @[Top.scala 172:12]
  assign n141_I_2_0_0_0 = n125_O_2_0_0_0; // @[Top.scala 172:12]
  assign n141_I_2_0_0_1 = n125_O_2_0_0_1; // @[Top.scala 172:12]
  assign n141_I_2_0_0_2 = n125_O_2_0_0_2; // @[Top.scala 172:12]
  assign n141_I_2_0_1_0 = n125_O_2_0_1_0; // @[Top.scala 172:12]
  assign n141_I_2_0_1_1 = n125_O_2_0_1_1; // @[Top.scala 172:12]
  assign n141_I_2_0_1_2 = n125_O_2_0_1_2; // @[Top.scala 172:12]
  assign n141_I_2_0_2_0 = n125_O_2_0_2_0; // @[Top.scala 172:12]
  assign n141_I_2_0_2_1 = n125_O_2_0_2_1; // @[Top.scala 172:12]
  assign n141_I_2_0_2_2 = n125_O_2_0_2_2; // @[Top.scala 172:12]
  assign n141_I_3_0_0_0 = n125_O_3_0_0_0; // @[Top.scala 172:12]
  assign n141_I_3_0_0_1 = n125_O_3_0_0_1; // @[Top.scala 172:12]
  assign n141_I_3_0_0_2 = n125_O_3_0_0_2; // @[Top.scala 172:12]
  assign n141_I_3_0_1_0 = n125_O_3_0_1_0; // @[Top.scala 172:12]
  assign n141_I_3_0_1_1 = n125_O_3_0_1_1; // @[Top.scala 172:12]
  assign n141_I_3_0_1_2 = n125_O_3_0_1_2; // @[Top.scala 172:12]
  assign n141_I_3_0_2_0 = n125_O_3_0_2_0; // @[Top.scala 172:12]
  assign n141_I_3_0_2_1 = n125_O_3_0_2_1; // @[Top.scala 172:12]
  assign n141_I_3_0_2_2 = n125_O_3_0_2_2; // @[Top.scala 172:12]
  assign n141_I_4_0_0_0 = n125_O_4_0_0_0; // @[Top.scala 172:12]
  assign n141_I_4_0_0_1 = n125_O_4_0_0_1; // @[Top.scala 172:12]
  assign n141_I_4_0_0_2 = n125_O_4_0_0_2; // @[Top.scala 172:12]
  assign n141_I_4_0_1_0 = n125_O_4_0_1_0; // @[Top.scala 172:12]
  assign n141_I_4_0_1_1 = n125_O_4_0_1_1; // @[Top.scala 172:12]
  assign n141_I_4_0_1_2 = n125_O_4_0_1_2; // @[Top.scala 172:12]
  assign n141_I_4_0_2_0 = n125_O_4_0_2_0; // @[Top.scala 172:12]
  assign n141_I_4_0_2_1 = n125_O_4_0_2_1; // @[Top.scala 172:12]
  assign n141_I_4_0_2_2 = n125_O_4_0_2_2; // @[Top.scala 172:12]
  assign n141_I_5_0_0_0 = n125_O_5_0_0_0; // @[Top.scala 172:12]
  assign n141_I_5_0_0_1 = n125_O_5_0_0_1; // @[Top.scala 172:12]
  assign n141_I_5_0_0_2 = n125_O_5_0_0_2; // @[Top.scala 172:12]
  assign n141_I_5_0_1_0 = n125_O_5_0_1_0; // @[Top.scala 172:12]
  assign n141_I_5_0_1_1 = n125_O_5_0_1_1; // @[Top.scala 172:12]
  assign n141_I_5_0_1_2 = n125_O_5_0_1_2; // @[Top.scala 172:12]
  assign n141_I_5_0_2_0 = n125_O_5_0_2_0; // @[Top.scala 172:12]
  assign n141_I_5_0_2_1 = n125_O_5_0_2_1; // @[Top.scala 172:12]
  assign n141_I_5_0_2_2 = n125_O_5_0_2_2; // @[Top.scala 172:12]
  assign n141_I_6_0_0_0 = n125_O_6_0_0_0; // @[Top.scala 172:12]
  assign n141_I_6_0_0_1 = n125_O_6_0_0_1; // @[Top.scala 172:12]
  assign n141_I_6_0_0_2 = n125_O_6_0_0_2; // @[Top.scala 172:12]
  assign n141_I_6_0_1_0 = n125_O_6_0_1_0; // @[Top.scala 172:12]
  assign n141_I_6_0_1_1 = n125_O_6_0_1_1; // @[Top.scala 172:12]
  assign n141_I_6_0_1_2 = n125_O_6_0_1_2; // @[Top.scala 172:12]
  assign n141_I_6_0_2_0 = n125_O_6_0_2_0; // @[Top.scala 172:12]
  assign n141_I_6_0_2_1 = n125_O_6_0_2_1; // @[Top.scala 172:12]
  assign n141_I_6_0_2_2 = n125_O_6_0_2_2; // @[Top.scala 172:12]
  assign n141_I_7_0_0_0 = n125_O_7_0_0_0; // @[Top.scala 172:12]
  assign n141_I_7_0_0_1 = n125_O_7_0_0_1; // @[Top.scala 172:12]
  assign n141_I_7_0_0_2 = n125_O_7_0_0_2; // @[Top.scala 172:12]
  assign n141_I_7_0_1_0 = n125_O_7_0_1_0; // @[Top.scala 172:12]
  assign n141_I_7_0_1_1 = n125_O_7_0_1_1; // @[Top.scala 172:12]
  assign n141_I_7_0_1_2 = n125_O_7_0_1_2; // @[Top.scala 172:12]
  assign n141_I_7_0_2_0 = n125_O_7_0_2_0; // @[Top.scala 172:12]
  assign n141_I_7_0_2_1 = n125_O_7_0_2_1; // @[Top.scala 172:12]
  assign n141_I_7_0_2_2 = n125_O_7_0_2_2; // @[Top.scala 172:12]
  assign n141_I_8_0_0_0 = n125_O_8_0_0_0; // @[Top.scala 172:12]
  assign n141_I_8_0_0_1 = n125_O_8_0_0_1; // @[Top.scala 172:12]
  assign n141_I_8_0_0_2 = n125_O_8_0_0_2; // @[Top.scala 172:12]
  assign n141_I_8_0_1_0 = n125_O_8_0_1_0; // @[Top.scala 172:12]
  assign n141_I_8_0_1_1 = n125_O_8_0_1_1; // @[Top.scala 172:12]
  assign n141_I_8_0_1_2 = n125_O_8_0_1_2; // @[Top.scala 172:12]
  assign n141_I_8_0_2_0 = n125_O_8_0_2_0; // @[Top.scala 172:12]
  assign n141_I_8_0_2_1 = n125_O_8_0_2_1; // @[Top.scala 172:12]
  assign n141_I_8_0_2_2 = n125_O_8_0_2_2; // @[Top.scala 172:12]
  assign n141_I_9_0_0_0 = n125_O_9_0_0_0; // @[Top.scala 172:12]
  assign n141_I_9_0_0_1 = n125_O_9_0_0_1; // @[Top.scala 172:12]
  assign n141_I_9_0_0_2 = n125_O_9_0_0_2; // @[Top.scala 172:12]
  assign n141_I_9_0_1_0 = n125_O_9_0_1_0; // @[Top.scala 172:12]
  assign n141_I_9_0_1_1 = n125_O_9_0_1_1; // @[Top.scala 172:12]
  assign n141_I_9_0_1_2 = n125_O_9_0_1_2; // @[Top.scala 172:12]
  assign n141_I_9_0_2_0 = n125_O_9_0_2_0; // @[Top.scala 172:12]
  assign n141_I_9_0_2_1 = n125_O_9_0_2_1; // @[Top.scala 172:12]
  assign n141_I_9_0_2_2 = n125_O_9_0_2_2; // @[Top.scala 172:12]
  assign n141_I_10_0_0_0 = n125_O_10_0_0_0; // @[Top.scala 172:12]
  assign n141_I_10_0_0_1 = n125_O_10_0_0_1; // @[Top.scala 172:12]
  assign n141_I_10_0_0_2 = n125_O_10_0_0_2; // @[Top.scala 172:12]
  assign n141_I_10_0_1_0 = n125_O_10_0_1_0; // @[Top.scala 172:12]
  assign n141_I_10_0_1_1 = n125_O_10_0_1_1; // @[Top.scala 172:12]
  assign n141_I_10_0_1_2 = n125_O_10_0_1_2; // @[Top.scala 172:12]
  assign n141_I_10_0_2_0 = n125_O_10_0_2_0; // @[Top.scala 172:12]
  assign n141_I_10_0_2_1 = n125_O_10_0_2_1; // @[Top.scala 172:12]
  assign n141_I_10_0_2_2 = n125_O_10_0_2_2; // @[Top.scala 172:12]
  assign n141_I_11_0_0_0 = n125_O_11_0_0_0; // @[Top.scala 172:12]
  assign n141_I_11_0_0_1 = n125_O_11_0_0_1; // @[Top.scala 172:12]
  assign n141_I_11_0_0_2 = n125_O_11_0_0_2; // @[Top.scala 172:12]
  assign n141_I_11_0_1_0 = n125_O_11_0_1_0; // @[Top.scala 172:12]
  assign n141_I_11_0_1_1 = n125_O_11_0_1_1; // @[Top.scala 172:12]
  assign n141_I_11_0_1_2 = n125_O_11_0_1_2; // @[Top.scala 172:12]
  assign n141_I_11_0_2_0 = n125_O_11_0_2_0; // @[Top.scala 172:12]
  assign n141_I_11_0_2_1 = n125_O_11_0_2_1; // @[Top.scala 172:12]
  assign n141_I_11_0_2_2 = n125_O_11_0_2_2; // @[Top.scala 172:12]
  assign n141_I_12_0_0_0 = n125_O_12_0_0_0; // @[Top.scala 172:12]
  assign n141_I_12_0_0_1 = n125_O_12_0_0_1; // @[Top.scala 172:12]
  assign n141_I_12_0_0_2 = n125_O_12_0_0_2; // @[Top.scala 172:12]
  assign n141_I_12_0_1_0 = n125_O_12_0_1_0; // @[Top.scala 172:12]
  assign n141_I_12_0_1_1 = n125_O_12_0_1_1; // @[Top.scala 172:12]
  assign n141_I_12_0_1_2 = n125_O_12_0_1_2; // @[Top.scala 172:12]
  assign n141_I_12_0_2_0 = n125_O_12_0_2_0; // @[Top.scala 172:12]
  assign n141_I_12_0_2_1 = n125_O_12_0_2_1; // @[Top.scala 172:12]
  assign n141_I_12_0_2_2 = n125_O_12_0_2_2; // @[Top.scala 172:12]
  assign n141_I_13_0_0_0 = n125_O_13_0_0_0; // @[Top.scala 172:12]
  assign n141_I_13_0_0_1 = n125_O_13_0_0_1; // @[Top.scala 172:12]
  assign n141_I_13_0_0_2 = n125_O_13_0_0_2; // @[Top.scala 172:12]
  assign n141_I_13_0_1_0 = n125_O_13_0_1_0; // @[Top.scala 172:12]
  assign n141_I_13_0_1_1 = n125_O_13_0_1_1; // @[Top.scala 172:12]
  assign n141_I_13_0_1_2 = n125_O_13_0_1_2; // @[Top.scala 172:12]
  assign n141_I_13_0_2_0 = n125_O_13_0_2_0; // @[Top.scala 172:12]
  assign n141_I_13_0_2_1 = n125_O_13_0_2_1; // @[Top.scala 172:12]
  assign n141_I_13_0_2_2 = n125_O_13_0_2_2; // @[Top.scala 172:12]
  assign n141_I_14_0_0_0 = n125_O_14_0_0_0; // @[Top.scala 172:12]
  assign n141_I_14_0_0_1 = n125_O_14_0_0_1; // @[Top.scala 172:12]
  assign n141_I_14_0_0_2 = n125_O_14_0_0_2; // @[Top.scala 172:12]
  assign n141_I_14_0_1_0 = n125_O_14_0_1_0; // @[Top.scala 172:12]
  assign n141_I_14_0_1_1 = n125_O_14_0_1_1; // @[Top.scala 172:12]
  assign n141_I_14_0_1_2 = n125_O_14_0_1_2; // @[Top.scala 172:12]
  assign n141_I_14_0_2_0 = n125_O_14_0_2_0; // @[Top.scala 172:12]
  assign n141_I_14_0_2_1 = n125_O_14_0_2_1; // @[Top.scala 172:12]
  assign n141_I_14_0_2_2 = n125_O_14_0_2_2; // @[Top.scala 172:12]
  assign n141_I_15_0_0_0 = n125_O_15_0_0_0; // @[Top.scala 172:12]
  assign n141_I_15_0_0_1 = n125_O_15_0_0_1; // @[Top.scala 172:12]
  assign n141_I_15_0_0_2 = n125_O_15_0_0_2; // @[Top.scala 172:12]
  assign n141_I_15_0_1_0 = n125_O_15_0_1_0; // @[Top.scala 172:12]
  assign n141_I_15_0_1_1 = n125_O_15_0_1_1; // @[Top.scala 172:12]
  assign n141_I_15_0_1_2 = n125_O_15_0_1_2; // @[Top.scala 172:12]
  assign n141_I_15_0_2_0 = n125_O_15_0_2_0; // @[Top.scala 172:12]
  assign n141_I_15_0_2_1 = n125_O_15_0_2_1; // @[Top.scala 172:12]
  assign n141_I_15_0_2_2 = n125_O_15_0_2_2; // @[Top.scala 172:12]
  assign n183_clock = clock;
  assign n183_reset = reset;
  assign n183_valid_up = n141_valid_down; // @[Top.scala 176:19]
  assign n183_I_0_0_0 = n141_O_0_0_0; // @[Top.scala 175:12]
  assign n183_I_0_0_1 = n141_O_0_0_1; // @[Top.scala 175:12]
  assign n183_I_0_0_2 = n141_O_0_0_2; // @[Top.scala 175:12]
  assign n183_I_0_1_0 = n141_O_0_1_0; // @[Top.scala 175:12]
  assign n183_I_0_1_1 = n141_O_0_1_1; // @[Top.scala 175:12]
  assign n183_I_0_1_2 = n141_O_0_1_2; // @[Top.scala 175:12]
  assign n183_I_0_2_0 = n141_O_0_2_0; // @[Top.scala 175:12]
  assign n183_I_0_2_1 = n141_O_0_2_1; // @[Top.scala 175:12]
  assign n183_I_0_2_2 = n141_O_0_2_2; // @[Top.scala 175:12]
  assign n183_I_1_0_0 = n141_O_1_0_0; // @[Top.scala 175:12]
  assign n183_I_1_0_1 = n141_O_1_0_1; // @[Top.scala 175:12]
  assign n183_I_1_0_2 = n141_O_1_0_2; // @[Top.scala 175:12]
  assign n183_I_1_1_0 = n141_O_1_1_0; // @[Top.scala 175:12]
  assign n183_I_1_1_1 = n141_O_1_1_1; // @[Top.scala 175:12]
  assign n183_I_1_1_2 = n141_O_1_1_2; // @[Top.scala 175:12]
  assign n183_I_1_2_0 = n141_O_1_2_0; // @[Top.scala 175:12]
  assign n183_I_1_2_1 = n141_O_1_2_1; // @[Top.scala 175:12]
  assign n183_I_1_2_2 = n141_O_1_2_2; // @[Top.scala 175:12]
  assign n183_I_2_0_0 = n141_O_2_0_0; // @[Top.scala 175:12]
  assign n183_I_2_0_1 = n141_O_2_0_1; // @[Top.scala 175:12]
  assign n183_I_2_0_2 = n141_O_2_0_2; // @[Top.scala 175:12]
  assign n183_I_2_1_0 = n141_O_2_1_0; // @[Top.scala 175:12]
  assign n183_I_2_1_1 = n141_O_2_1_1; // @[Top.scala 175:12]
  assign n183_I_2_1_2 = n141_O_2_1_2; // @[Top.scala 175:12]
  assign n183_I_2_2_0 = n141_O_2_2_0; // @[Top.scala 175:12]
  assign n183_I_2_2_1 = n141_O_2_2_1; // @[Top.scala 175:12]
  assign n183_I_2_2_2 = n141_O_2_2_2; // @[Top.scala 175:12]
  assign n183_I_3_0_0 = n141_O_3_0_0; // @[Top.scala 175:12]
  assign n183_I_3_0_1 = n141_O_3_0_1; // @[Top.scala 175:12]
  assign n183_I_3_0_2 = n141_O_3_0_2; // @[Top.scala 175:12]
  assign n183_I_3_1_0 = n141_O_3_1_0; // @[Top.scala 175:12]
  assign n183_I_3_1_1 = n141_O_3_1_1; // @[Top.scala 175:12]
  assign n183_I_3_1_2 = n141_O_3_1_2; // @[Top.scala 175:12]
  assign n183_I_3_2_0 = n141_O_3_2_0; // @[Top.scala 175:12]
  assign n183_I_3_2_1 = n141_O_3_2_1; // @[Top.scala 175:12]
  assign n183_I_3_2_2 = n141_O_3_2_2; // @[Top.scala 175:12]
  assign n183_I_4_0_0 = n141_O_4_0_0; // @[Top.scala 175:12]
  assign n183_I_4_0_1 = n141_O_4_0_1; // @[Top.scala 175:12]
  assign n183_I_4_0_2 = n141_O_4_0_2; // @[Top.scala 175:12]
  assign n183_I_4_1_0 = n141_O_4_1_0; // @[Top.scala 175:12]
  assign n183_I_4_1_1 = n141_O_4_1_1; // @[Top.scala 175:12]
  assign n183_I_4_1_2 = n141_O_4_1_2; // @[Top.scala 175:12]
  assign n183_I_4_2_0 = n141_O_4_2_0; // @[Top.scala 175:12]
  assign n183_I_4_2_1 = n141_O_4_2_1; // @[Top.scala 175:12]
  assign n183_I_4_2_2 = n141_O_4_2_2; // @[Top.scala 175:12]
  assign n183_I_5_0_0 = n141_O_5_0_0; // @[Top.scala 175:12]
  assign n183_I_5_0_1 = n141_O_5_0_1; // @[Top.scala 175:12]
  assign n183_I_5_0_2 = n141_O_5_0_2; // @[Top.scala 175:12]
  assign n183_I_5_1_0 = n141_O_5_1_0; // @[Top.scala 175:12]
  assign n183_I_5_1_1 = n141_O_5_1_1; // @[Top.scala 175:12]
  assign n183_I_5_1_2 = n141_O_5_1_2; // @[Top.scala 175:12]
  assign n183_I_5_2_0 = n141_O_5_2_0; // @[Top.scala 175:12]
  assign n183_I_5_2_1 = n141_O_5_2_1; // @[Top.scala 175:12]
  assign n183_I_5_2_2 = n141_O_5_2_2; // @[Top.scala 175:12]
  assign n183_I_6_0_0 = n141_O_6_0_0; // @[Top.scala 175:12]
  assign n183_I_6_0_1 = n141_O_6_0_1; // @[Top.scala 175:12]
  assign n183_I_6_0_2 = n141_O_6_0_2; // @[Top.scala 175:12]
  assign n183_I_6_1_0 = n141_O_6_1_0; // @[Top.scala 175:12]
  assign n183_I_6_1_1 = n141_O_6_1_1; // @[Top.scala 175:12]
  assign n183_I_6_1_2 = n141_O_6_1_2; // @[Top.scala 175:12]
  assign n183_I_6_2_0 = n141_O_6_2_0; // @[Top.scala 175:12]
  assign n183_I_6_2_1 = n141_O_6_2_1; // @[Top.scala 175:12]
  assign n183_I_6_2_2 = n141_O_6_2_2; // @[Top.scala 175:12]
  assign n183_I_7_0_0 = n141_O_7_0_0; // @[Top.scala 175:12]
  assign n183_I_7_0_1 = n141_O_7_0_1; // @[Top.scala 175:12]
  assign n183_I_7_0_2 = n141_O_7_0_2; // @[Top.scala 175:12]
  assign n183_I_7_1_0 = n141_O_7_1_0; // @[Top.scala 175:12]
  assign n183_I_7_1_1 = n141_O_7_1_1; // @[Top.scala 175:12]
  assign n183_I_7_1_2 = n141_O_7_1_2; // @[Top.scala 175:12]
  assign n183_I_7_2_0 = n141_O_7_2_0; // @[Top.scala 175:12]
  assign n183_I_7_2_1 = n141_O_7_2_1; // @[Top.scala 175:12]
  assign n183_I_7_2_2 = n141_O_7_2_2; // @[Top.scala 175:12]
  assign n183_I_8_0_0 = n141_O_8_0_0; // @[Top.scala 175:12]
  assign n183_I_8_0_1 = n141_O_8_0_1; // @[Top.scala 175:12]
  assign n183_I_8_0_2 = n141_O_8_0_2; // @[Top.scala 175:12]
  assign n183_I_8_1_0 = n141_O_8_1_0; // @[Top.scala 175:12]
  assign n183_I_8_1_1 = n141_O_8_1_1; // @[Top.scala 175:12]
  assign n183_I_8_1_2 = n141_O_8_1_2; // @[Top.scala 175:12]
  assign n183_I_8_2_0 = n141_O_8_2_0; // @[Top.scala 175:12]
  assign n183_I_8_2_1 = n141_O_8_2_1; // @[Top.scala 175:12]
  assign n183_I_8_2_2 = n141_O_8_2_2; // @[Top.scala 175:12]
  assign n183_I_9_0_0 = n141_O_9_0_0; // @[Top.scala 175:12]
  assign n183_I_9_0_1 = n141_O_9_0_1; // @[Top.scala 175:12]
  assign n183_I_9_0_2 = n141_O_9_0_2; // @[Top.scala 175:12]
  assign n183_I_9_1_0 = n141_O_9_1_0; // @[Top.scala 175:12]
  assign n183_I_9_1_1 = n141_O_9_1_1; // @[Top.scala 175:12]
  assign n183_I_9_1_2 = n141_O_9_1_2; // @[Top.scala 175:12]
  assign n183_I_9_2_0 = n141_O_9_2_0; // @[Top.scala 175:12]
  assign n183_I_9_2_1 = n141_O_9_2_1; // @[Top.scala 175:12]
  assign n183_I_9_2_2 = n141_O_9_2_2; // @[Top.scala 175:12]
  assign n183_I_10_0_0 = n141_O_10_0_0; // @[Top.scala 175:12]
  assign n183_I_10_0_1 = n141_O_10_0_1; // @[Top.scala 175:12]
  assign n183_I_10_0_2 = n141_O_10_0_2; // @[Top.scala 175:12]
  assign n183_I_10_1_0 = n141_O_10_1_0; // @[Top.scala 175:12]
  assign n183_I_10_1_1 = n141_O_10_1_1; // @[Top.scala 175:12]
  assign n183_I_10_1_2 = n141_O_10_1_2; // @[Top.scala 175:12]
  assign n183_I_10_2_0 = n141_O_10_2_0; // @[Top.scala 175:12]
  assign n183_I_10_2_1 = n141_O_10_2_1; // @[Top.scala 175:12]
  assign n183_I_10_2_2 = n141_O_10_2_2; // @[Top.scala 175:12]
  assign n183_I_11_0_0 = n141_O_11_0_0; // @[Top.scala 175:12]
  assign n183_I_11_0_1 = n141_O_11_0_1; // @[Top.scala 175:12]
  assign n183_I_11_0_2 = n141_O_11_0_2; // @[Top.scala 175:12]
  assign n183_I_11_1_0 = n141_O_11_1_0; // @[Top.scala 175:12]
  assign n183_I_11_1_1 = n141_O_11_1_1; // @[Top.scala 175:12]
  assign n183_I_11_1_2 = n141_O_11_1_2; // @[Top.scala 175:12]
  assign n183_I_11_2_0 = n141_O_11_2_0; // @[Top.scala 175:12]
  assign n183_I_11_2_1 = n141_O_11_2_1; // @[Top.scala 175:12]
  assign n183_I_11_2_2 = n141_O_11_2_2; // @[Top.scala 175:12]
  assign n183_I_12_0_0 = n141_O_12_0_0; // @[Top.scala 175:12]
  assign n183_I_12_0_1 = n141_O_12_0_1; // @[Top.scala 175:12]
  assign n183_I_12_0_2 = n141_O_12_0_2; // @[Top.scala 175:12]
  assign n183_I_12_1_0 = n141_O_12_1_0; // @[Top.scala 175:12]
  assign n183_I_12_1_1 = n141_O_12_1_1; // @[Top.scala 175:12]
  assign n183_I_12_1_2 = n141_O_12_1_2; // @[Top.scala 175:12]
  assign n183_I_12_2_0 = n141_O_12_2_0; // @[Top.scala 175:12]
  assign n183_I_12_2_1 = n141_O_12_2_1; // @[Top.scala 175:12]
  assign n183_I_12_2_2 = n141_O_12_2_2; // @[Top.scala 175:12]
  assign n183_I_13_0_0 = n141_O_13_0_0; // @[Top.scala 175:12]
  assign n183_I_13_0_1 = n141_O_13_0_1; // @[Top.scala 175:12]
  assign n183_I_13_0_2 = n141_O_13_0_2; // @[Top.scala 175:12]
  assign n183_I_13_1_0 = n141_O_13_1_0; // @[Top.scala 175:12]
  assign n183_I_13_1_1 = n141_O_13_1_1; // @[Top.scala 175:12]
  assign n183_I_13_1_2 = n141_O_13_1_2; // @[Top.scala 175:12]
  assign n183_I_13_2_0 = n141_O_13_2_0; // @[Top.scala 175:12]
  assign n183_I_13_2_1 = n141_O_13_2_1; // @[Top.scala 175:12]
  assign n183_I_13_2_2 = n141_O_13_2_2; // @[Top.scala 175:12]
  assign n183_I_14_0_0 = n141_O_14_0_0; // @[Top.scala 175:12]
  assign n183_I_14_0_1 = n141_O_14_0_1; // @[Top.scala 175:12]
  assign n183_I_14_0_2 = n141_O_14_0_2; // @[Top.scala 175:12]
  assign n183_I_14_1_0 = n141_O_14_1_0; // @[Top.scala 175:12]
  assign n183_I_14_1_1 = n141_O_14_1_1; // @[Top.scala 175:12]
  assign n183_I_14_1_2 = n141_O_14_1_2; // @[Top.scala 175:12]
  assign n183_I_14_2_0 = n141_O_14_2_0; // @[Top.scala 175:12]
  assign n183_I_14_2_1 = n141_O_14_2_1; // @[Top.scala 175:12]
  assign n183_I_14_2_2 = n141_O_14_2_2; // @[Top.scala 175:12]
  assign n183_I_15_0_0 = n141_O_15_0_0; // @[Top.scala 175:12]
  assign n183_I_15_0_1 = n141_O_15_0_1; // @[Top.scala 175:12]
  assign n183_I_15_0_2 = n141_O_15_0_2; // @[Top.scala 175:12]
  assign n183_I_15_1_0 = n141_O_15_1_0; // @[Top.scala 175:12]
  assign n183_I_15_1_1 = n141_O_15_1_1; // @[Top.scala 175:12]
  assign n183_I_15_1_2 = n141_O_15_1_2; // @[Top.scala 175:12]
  assign n183_I_15_2_0 = n141_O_15_2_0; // @[Top.scala 175:12]
  assign n183_I_15_2_1 = n141_O_15_2_1; // @[Top.scala 175:12]
  assign n183_I_15_2_2 = n141_O_15_2_2; // @[Top.scala 175:12]
  assign n184_clock = clock;
  assign n184_reset = reset;
  assign n184_valid_up = n1_valid_down; // @[Top.scala 179:19]
  assign n184_I_0_0_0 = n1_O_0_0_0; // @[Top.scala 178:12]
  assign n184_I_1_0_0 = n1_O_1_0_0; // @[Top.scala 178:12]
  assign n184_I_2_0_0 = n1_O_2_0_0; // @[Top.scala 178:12]
  assign n184_I_3_0_0 = n1_O_3_0_0; // @[Top.scala 178:12]
  assign n184_I_4_0_0 = n1_O_4_0_0; // @[Top.scala 178:12]
  assign n184_I_5_0_0 = n1_O_5_0_0; // @[Top.scala 178:12]
  assign n184_I_6_0_0 = n1_O_6_0_0; // @[Top.scala 178:12]
  assign n184_I_7_0_0 = n1_O_7_0_0; // @[Top.scala 178:12]
  assign n184_I_8_0_0 = n1_O_8_0_0; // @[Top.scala 178:12]
  assign n184_I_9_0_0 = n1_O_9_0_0; // @[Top.scala 178:12]
  assign n184_I_10_0_0 = n1_O_10_0_0; // @[Top.scala 178:12]
  assign n184_I_11_0_0 = n1_O_11_0_0; // @[Top.scala 178:12]
  assign n184_I_12_0_0 = n1_O_12_0_0; // @[Top.scala 178:12]
  assign n184_I_13_0_0 = n1_O_13_0_0; // @[Top.scala 178:12]
  assign n184_I_14_0_0 = n1_O_14_0_0; // @[Top.scala 178:12]
  assign n184_I_15_0_0 = n1_O_15_0_0; // @[Top.scala 178:12]
  assign n185_clock = clock;
  assign n185_reset = reset;
  assign n185_valid_up = n183_valid_down & n184_valid_down; // @[Top.scala 183:19]
  assign n185_I0_0_0_0 = n183_O_0_0_0; // @[Top.scala 181:13]
  assign n185_I0_1_0_0 = n183_O_1_0_0; // @[Top.scala 181:13]
  assign n185_I0_2_0_0 = n183_O_2_0_0; // @[Top.scala 181:13]
  assign n185_I0_3_0_0 = n183_O_3_0_0; // @[Top.scala 181:13]
  assign n185_I0_4_0_0 = n183_O_4_0_0; // @[Top.scala 181:13]
  assign n185_I0_5_0_0 = n183_O_5_0_0; // @[Top.scala 181:13]
  assign n185_I0_6_0_0 = n183_O_6_0_0; // @[Top.scala 181:13]
  assign n185_I0_7_0_0 = n183_O_7_0_0; // @[Top.scala 181:13]
  assign n185_I0_8_0_0 = n183_O_8_0_0; // @[Top.scala 181:13]
  assign n185_I0_9_0_0 = n183_O_9_0_0; // @[Top.scala 181:13]
  assign n185_I0_10_0_0 = n183_O_10_0_0; // @[Top.scala 181:13]
  assign n185_I0_11_0_0 = n183_O_11_0_0; // @[Top.scala 181:13]
  assign n185_I0_12_0_0 = n183_O_12_0_0; // @[Top.scala 181:13]
  assign n185_I0_13_0_0 = n183_O_13_0_0; // @[Top.scala 181:13]
  assign n185_I0_14_0_0 = n183_O_14_0_0; // @[Top.scala 181:13]
  assign n185_I0_15_0_0 = n183_O_15_0_0; // @[Top.scala 181:13]
  assign n185_I1_0_0_0 = n184_O_0_0_0; // @[Top.scala 182:13]
  assign n185_I1_1_0_0 = n184_O_1_0_0; // @[Top.scala 182:13]
  assign n185_I1_2_0_0 = n184_O_2_0_0; // @[Top.scala 182:13]
  assign n185_I1_3_0_0 = n184_O_3_0_0; // @[Top.scala 182:13]
  assign n185_I1_4_0_0 = n184_O_4_0_0; // @[Top.scala 182:13]
  assign n185_I1_5_0_0 = n184_O_5_0_0; // @[Top.scala 182:13]
  assign n185_I1_6_0_0 = n184_O_6_0_0; // @[Top.scala 182:13]
  assign n185_I1_7_0_0 = n184_O_7_0_0; // @[Top.scala 182:13]
  assign n185_I1_8_0_0 = n184_O_8_0_0; // @[Top.scala 182:13]
  assign n185_I1_9_0_0 = n184_O_9_0_0; // @[Top.scala 182:13]
  assign n185_I1_10_0_0 = n184_O_10_0_0; // @[Top.scala 182:13]
  assign n185_I1_11_0_0 = n184_O_11_0_0; // @[Top.scala 182:13]
  assign n185_I1_12_0_0 = n184_O_12_0_0; // @[Top.scala 182:13]
  assign n185_I1_13_0_0 = n184_O_13_0_0; // @[Top.scala 182:13]
  assign n185_I1_14_0_0 = n184_O_14_0_0; // @[Top.scala 182:13]
  assign n185_I1_15_0_0 = n184_O_15_0_0; // @[Top.scala 182:13]
  assign n217_clock = clock;
  assign n217_valid_up = n185_valid_down; // @[Top.scala 186:19]
  assign n217_I_0_0_0 = n185_O_0_0_0; // @[Top.scala 185:12]
  assign n217_I_1_0_0 = n185_O_1_0_0; // @[Top.scala 185:12]
  assign n217_I_2_0_0 = n185_O_2_0_0; // @[Top.scala 185:12]
  assign n217_I_3_0_0 = n185_O_3_0_0; // @[Top.scala 185:12]
  assign n217_I_4_0_0 = n185_O_4_0_0; // @[Top.scala 185:12]
  assign n217_I_5_0_0 = n185_O_5_0_0; // @[Top.scala 185:12]
  assign n217_I_6_0_0 = n185_O_6_0_0; // @[Top.scala 185:12]
  assign n217_I_7_0_0 = n185_O_7_0_0; // @[Top.scala 185:12]
  assign n217_I_8_0_0 = n185_O_8_0_0; // @[Top.scala 185:12]
  assign n217_I_9_0_0 = n185_O_9_0_0; // @[Top.scala 185:12]
  assign n217_I_10_0_0 = n185_O_10_0_0; // @[Top.scala 185:12]
  assign n217_I_11_0_0 = n185_O_11_0_0; // @[Top.scala 185:12]
  assign n217_I_12_0_0 = n185_O_12_0_0; // @[Top.scala 185:12]
  assign n217_I_13_0_0 = n185_O_13_0_0; // @[Top.scala 185:12]
  assign n217_I_14_0_0 = n185_O_14_0_0; // @[Top.scala 185:12]
  assign n217_I_15_0_0 = n185_O_15_0_0; // @[Top.scala 185:12]
  assign n218_clock = clock;
  assign n218_valid_up = n217_valid_down; // @[Top.scala 189:19]
  assign n218_I_0_0_0 = n217_O_0_0_0; // @[Top.scala 188:12]
  assign n218_I_1_0_0 = n217_O_1_0_0; // @[Top.scala 188:12]
  assign n218_I_2_0_0 = n217_O_2_0_0; // @[Top.scala 188:12]
  assign n218_I_3_0_0 = n217_O_3_0_0; // @[Top.scala 188:12]
  assign n218_I_4_0_0 = n217_O_4_0_0; // @[Top.scala 188:12]
  assign n218_I_5_0_0 = n217_O_5_0_0; // @[Top.scala 188:12]
  assign n218_I_6_0_0 = n217_O_6_0_0; // @[Top.scala 188:12]
  assign n218_I_7_0_0 = n217_O_7_0_0; // @[Top.scala 188:12]
  assign n218_I_8_0_0 = n217_O_8_0_0; // @[Top.scala 188:12]
  assign n218_I_9_0_0 = n217_O_9_0_0; // @[Top.scala 188:12]
  assign n218_I_10_0_0 = n217_O_10_0_0; // @[Top.scala 188:12]
  assign n218_I_11_0_0 = n217_O_11_0_0; // @[Top.scala 188:12]
  assign n218_I_12_0_0 = n217_O_12_0_0; // @[Top.scala 188:12]
  assign n218_I_13_0_0 = n217_O_13_0_0; // @[Top.scala 188:12]
  assign n218_I_14_0_0 = n217_O_14_0_0; // @[Top.scala 188:12]
  assign n218_I_15_0_0 = n217_O_15_0_0; // @[Top.scala 188:12]
  assign n219_clock = clock;
  assign n219_valid_up = n218_valid_down; // @[Top.scala 192:19]
  assign n219_I_0_0_0 = n218_O_0_0_0; // @[Top.scala 191:12]
  assign n219_I_1_0_0 = n218_O_1_0_0; // @[Top.scala 191:12]
  assign n219_I_2_0_0 = n218_O_2_0_0; // @[Top.scala 191:12]
  assign n219_I_3_0_0 = n218_O_3_0_0; // @[Top.scala 191:12]
  assign n219_I_4_0_0 = n218_O_4_0_0; // @[Top.scala 191:12]
  assign n219_I_5_0_0 = n218_O_5_0_0; // @[Top.scala 191:12]
  assign n219_I_6_0_0 = n218_O_6_0_0; // @[Top.scala 191:12]
  assign n219_I_7_0_0 = n218_O_7_0_0; // @[Top.scala 191:12]
  assign n219_I_8_0_0 = n218_O_8_0_0; // @[Top.scala 191:12]
  assign n219_I_9_0_0 = n218_O_9_0_0; // @[Top.scala 191:12]
  assign n219_I_10_0_0 = n218_O_10_0_0; // @[Top.scala 191:12]
  assign n219_I_11_0_0 = n218_O_11_0_0; // @[Top.scala 191:12]
  assign n219_I_12_0_0 = n218_O_12_0_0; // @[Top.scala 191:12]
  assign n219_I_13_0_0 = n218_O_13_0_0; // @[Top.scala 191:12]
  assign n219_I_14_0_0 = n218_O_14_0_0; // @[Top.scala 191:12]
  assign n219_I_15_0_0 = n218_O_15_0_0; // @[Top.scala 191:12]
endmodule
